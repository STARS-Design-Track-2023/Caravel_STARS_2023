VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO outel8227
  CLASS BLOCK ;
  FOREIGN outel8227 ;
  ORIGIN 0.000 0.000 ;
  SIZE 212.745 BY 223.465 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 208.745 47.640 212.745 48.240 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.745 6.840 212.745 7.440 ;
    END
  END cs
  PIN dataBusIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END dataBusIn[0]
  PIN dataBusIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END dataBusIn[1]
  PIN dataBusIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 219.465 193.570 223.465 ;
    END
  END dataBusIn[2]
  PIN dataBusIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END dataBusIn[3]
  PIN dataBusIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 219.465 154.930 223.465 ;
    END
  END dataBusIn[4]
  PIN dataBusIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 219.465 45.450 223.465 ;
    END
  END dataBusIn[5]
  PIN dataBusIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END dataBusIn[6]
  PIN dataBusIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 208.745 27.240 212.745 27.840 ;
    END
  END dataBusIn[7]
  PIN dataBusOut[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 208.745 183.640 212.745 184.240 ;
    END
  END dataBusOut[0]
  PIN dataBusOut[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END dataBusOut[1]
  PIN dataBusOut[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dataBusOut[2]
  PIN dataBusOut[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 208.745 163.240 212.745 163.840 ;
    END
  END dataBusOut[3]
  PIN dataBusOut[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END dataBusOut[4]
  PIN dataBusOut[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END dataBusOut[5]
  PIN dataBusOut[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 208.745 204.040 212.745 204.640 ;
    END
  END dataBusOut[6]
  PIN dataBusOut[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 219.465 6.810 223.465 ;
    END
  END dataBusOut[7]
  PIN dataBusSelect
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.970 219.465 174.250 223.465 ;
    END
  END dataBusSelect
  PIN gpio[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 219.465 119.510 223.465 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 219.465 100.190 223.465 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 219.465 26.130 223.465 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END gpio[16]
  PIN gpio[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 208.745 146.240 212.745 146.840 ;
    END
  END gpio[17]
  PIN gpio[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gpio[18]
  PIN gpio[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    PORT
      LAYER met3 ;
        RECT 208.745 125.840 212.745 126.440 ;
    END
  END gpio[19]
  PIN gpio[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END gpio[1]
  PIN gpio[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 219.465 138.830 223.465 ;
    END
  END gpio[20]
  PIN gpio[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met3 ;
        RECT 208.745 68.040 212.745 68.640 ;
    END
  END gpio[21]
  PIN gpio[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END gpio[22]
  PIN gpio[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gpio[23]
  PIN gpio[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END gpio[24]
  PIN gpio[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.745 85.040 212.745 85.640 ;
    END
  END gpio[25]
  PIN gpio[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 219.465 209.670 223.465 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 219.465 64.770 223.465 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 219.465 80.870 223.465 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 208.745 105.440 212.745 106.040 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 212.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 212.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 207.000 212.245 ;
      LAYER met1 ;
        RECT 0.070 10.640 209.690 212.400 ;
      LAYER met2 ;
        RECT 0.100 219.185 6.250 220.050 ;
        RECT 7.090 219.185 25.570 220.050 ;
        RECT 26.410 219.185 44.890 220.050 ;
        RECT 45.730 219.185 64.210 220.050 ;
        RECT 65.050 219.185 80.310 220.050 ;
        RECT 81.150 219.185 99.630 220.050 ;
        RECT 100.470 219.185 118.950 220.050 ;
        RECT 119.790 219.185 138.270 220.050 ;
        RECT 139.110 219.185 154.370 220.050 ;
        RECT 155.210 219.185 173.690 220.050 ;
        RECT 174.530 219.185 193.010 220.050 ;
        RECT 193.850 219.185 209.110 220.050 ;
        RECT 0.100 4.280 209.670 219.185 ;
        RECT 0.650 4.000 15.910 4.280 ;
        RECT 16.750 4.000 35.230 4.280 ;
        RECT 36.070 4.000 54.550 4.280 ;
        RECT 55.390 4.000 70.650 4.280 ;
        RECT 71.490 4.000 89.970 4.280 ;
        RECT 90.810 4.000 109.290 4.280 ;
        RECT 110.130 4.000 128.610 4.280 ;
        RECT 129.450 4.000 144.710 4.280 ;
        RECT 145.550 4.000 164.030 4.280 ;
        RECT 164.870 4.000 183.350 4.280 ;
        RECT 184.190 4.000 202.670 4.280 ;
        RECT 203.510 4.000 209.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 213.840 209.695 214.705 ;
        RECT 3.990 205.040 209.695 213.840 ;
        RECT 3.990 203.640 208.345 205.040 ;
        RECT 3.990 194.840 209.695 203.640 ;
        RECT 4.400 193.440 209.695 194.840 ;
        RECT 3.990 184.640 209.695 193.440 ;
        RECT 3.990 183.240 208.345 184.640 ;
        RECT 3.990 174.440 209.695 183.240 ;
        RECT 4.400 173.040 209.695 174.440 ;
        RECT 3.990 164.240 209.695 173.040 ;
        RECT 3.990 162.840 208.345 164.240 ;
        RECT 3.990 154.040 209.695 162.840 ;
        RECT 4.400 152.640 209.695 154.040 ;
        RECT 3.990 147.240 209.695 152.640 ;
        RECT 3.990 145.840 208.345 147.240 ;
        RECT 3.990 137.040 209.695 145.840 ;
        RECT 4.400 135.640 209.695 137.040 ;
        RECT 3.990 126.840 209.695 135.640 ;
        RECT 3.990 125.440 208.345 126.840 ;
        RECT 3.990 116.640 209.695 125.440 ;
        RECT 4.400 115.240 209.695 116.640 ;
        RECT 3.990 106.440 209.695 115.240 ;
        RECT 3.990 105.040 208.345 106.440 ;
        RECT 3.990 96.240 209.695 105.040 ;
        RECT 4.400 94.840 209.695 96.240 ;
        RECT 3.990 86.040 209.695 94.840 ;
        RECT 3.990 84.640 208.345 86.040 ;
        RECT 3.990 75.840 209.695 84.640 ;
        RECT 4.400 74.440 209.695 75.840 ;
        RECT 3.990 69.040 209.695 74.440 ;
        RECT 3.990 67.640 208.345 69.040 ;
        RECT 3.990 58.840 209.695 67.640 ;
        RECT 4.400 57.440 209.695 58.840 ;
        RECT 3.990 48.640 209.695 57.440 ;
        RECT 3.990 47.240 208.345 48.640 ;
        RECT 3.990 38.440 209.695 47.240 ;
        RECT 4.400 37.040 209.695 38.440 ;
        RECT 3.990 28.240 209.695 37.040 ;
        RECT 3.990 26.840 208.345 28.240 ;
        RECT 3.990 18.040 209.695 26.840 ;
        RECT 4.400 16.640 209.695 18.040 ;
        RECT 3.990 10.715 209.695 16.640 ;
      LAYER met4 ;
        RECT 26.975 17.855 97.440 211.305 ;
        RECT 99.840 17.855 174.240 211.305 ;
        RECT 176.640 17.855 196.585 211.305 ;
  END
END outel8227
END LIBRARY

