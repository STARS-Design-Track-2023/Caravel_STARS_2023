* NGSPICE file created from silly_synthesizer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt silly_synthesizer VGND VPWR clk cs gpio[0] gpio[10] gpio[11] gpio[12] gpio[13]
+ gpio[14] gpio[15] gpio[16] gpio[1] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7]
+ gpio[8] gpio[9] nrst pwm
X_2037_ _0487_ _1084_ _0488_ _0405_ net263 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a32o_1
X_2106_ net247 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2939_ clknet_leaf_12_clk _0145_ net39 VGND VGND VPWR VPWR outputs.divider_buffer\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2655_ _0979_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_1606_ outputs.divider_buffer\[3\] _1214_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__nor2_1
X_2724_ clknet_leaf_32_clk inputs.random_update_clock.next_count\[1\] net27 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2586_ net225 net294 _0936_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__mux2_1
X_1537_ outputs.sig_gen.count\[12\] _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__or2_1
X_1468_ outputs.divider_buffer\[3\] VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__inv_2
X_1399_ inputs.random_update_clock.count\[16\] _1060_ net284 VGND VGND VPWR VPWR _1062_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold170 outputs.div.oscillator_out\[2\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold192 _0526_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 outputs.output_gen.count\[4\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2440_ _0658_ _0811_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1322_ _1005_ net16 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__and2b_1
X_2371_ _0561_ _0540_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2569_ net223 net127 _0925_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__mux2_1
X_2638_ outputs.shaper.count\[9\] net209 _0966_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2707_ clknet_leaf_37_clk net84 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1940_ _0417_ _0418_ _0423_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1871_ _0362_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2423_ net253 _0827_ _0645_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1305_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__clkbuf_4
X_2285_ _0696_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_2354_ _0231_ _0680_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _0506_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nand2_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2972_ clknet_leaf_6_clk _0178_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_1923_ _0410_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1854_ outputs.div.a\[10\] _0347_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor2_1
X_1785_ _0277_ _0285_ _0286_ _0252_ net154 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2406_ _0538_ _0536_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2268_ _0622_ _0679_ _0624_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
X_2199_ inputs.key_encoder.sync_keys\[12\] _0596_ _0586_ VGND VGND VPWR VPWR _0613_
+ sky130_fd_sc_hd__o21a_1
X_2337_ _0648_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold63 outputs.div.q\[19\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 outputs.div.oscillator_out\[6\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 outputs.div.q_out\[0\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold30 inputs.random_note_generator.out\[12\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 inputs.random_update_clock.count\[22\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _0060_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 outputs.div.a\[0\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ net296 inputs.down.in VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__and2b_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ outputs.scaled_buffer\[2\] net201 _0497_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__buf_2
X_2955_ clknet_leaf_5_clk _0161_ VGND VGND VPWR VPWR outputs.signal_buffer2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2886_ clknet_leaf_8_clk outputs.sig_gen.next_count\[15\] net44 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[15\] sky130_fd_sc_hd__dfrtp_2
X_1906_ outputs.div.m\[15\] _0386_ _0320_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o21a_1
X_1837_ _0324_ _0327_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o21ai_1
X_1768_ outputs.div.m\[3\] _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1699_ _0217_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR pwm sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1622_ _1193_ _1194_ _1096_ outputs.shaper.count\[16\] VGND VGND VPWR VPWR _1236_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ _0768_ _0983_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nand2_1
X_2740_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[17\] net29 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[17\] sky130_fd_sc_hd__dfrtp_1
X_1553_ _1175_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
X_1484_ outputs.divider_buffer\[0\] VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__inv_2
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2036_ outputs.div.count\[1\] outputs.div.count\[0\] VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or2_1
X_2105_ net246 outputs.div.divisor\[11\] _0522_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2938_ clknet_leaf_12_clk _0144_ net39 VGND VGND VPWR VPWR outputs.divider_buffer\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2869_ clknet_leaf_26_clk outputs.output_gen.next_count\[6\] net49 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2723_ clknet_leaf_32_clk inputs.random_update_clock.next_count\[0\] net27 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[0\] sky130_fd_sc_hd__dfstp_1
X_2654_ outputs.shaper.count\[17\] net230 _1089_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__mux2_1
X_2585_ _0943_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
X_1605_ outputs.divider_buffer\[1\] _1217_ _1216_ _1218_ VGND VGND VPWR VPWR _1219_
+ sky130_fd_sc_hd__o211ai_1
X_1536_ _1116_ _1159_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1467_ _1094_ _1098_ _1102_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__or4_1
X_1398_ net168 _1060_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[16\]
+ sky130_fd_sc_hd__xor2_1
X_2019_ outputs.div.oscillator_out\[11\] _0475_ _0468_ net118 _0479_ VGND VGND VPWR
+ VPWR _0066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold160 outputs.signal_buffer2\[5\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 outputs.signal_buffer2\[0\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 outputs.divider_buffer2\[17\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 outputs.divider_buffer2\[12\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1321_ _1012_ VGND VGND VPWR VPWR inputs.keypad\[6\] sky130_fd_sc_hd__clkbuf_1
X_2370_ _0561_ _0776_ _0722_ _0650_ _0648_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2706_ clknet_leaf_37_clk net76 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2568_ net229 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
X_2637_ _0970_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
X_1519_ outputs.sig_gen.count\[6\] outputs.sig_gen.count\[7\] _1144_ VGND VGND VPWR
+ VPWR _1150_ sky130_fd_sc_hd__and3_1
X_2499_ net298 _0896_ _0855_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ _0339_ _0342_ _0348_ _0350_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2353_ _0626_ _0759_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__o21a_1
X_2422_ _0816_ _0822_ _0826_ _0642_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1304_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__clkbuf_4
X_2284_ net279 _0695_ _0645_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1999_ outputs.div.q\[9\] _0248_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1922_ _0400_ _0402_ _0398_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o21ai_1
X_2971_ clknet_leaf_4_clk _0177_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1853_ outputs.div.a\[10\] _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__nand2_2
X_1784_ _0280_ _0284_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2405_ _0568_ _0549_ _0662_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__or3_1
X_2336_ inputs.frequency_lut.rng\[3\] _0656_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2267_ _0668_ _0678_ _0237_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
X_2198_ _0602_ _0610_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold86 outputs.sample_rate.count\[4\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 outputs.div.q\[21\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _0066_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0061_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _0087_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 inputs.keypad_synchronizer.half_sync\[10\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 inputs.random_note_generator.out\[9\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 inputs.random_update_clock.next_count\[22\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ _0498_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
X_2121_ inputs.frequency_lut.rng\[2\] VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2954_ clknet_leaf_6_clk _0160_ VGND VGND VPWR VPWR outputs.signal_buffer2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2885_ clknet_leaf_5_clk outputs.sig_gen.next_count\[14\] net42 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[14\] sky130_fd_sc_hd__dfrtp_2
X_1905_ outputs.div.a\[15\] VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1836_ _0331_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1698_ outputs.div.m\[8\] net308 _1294_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
X_1767_ outputs.div.m\[2\] _0253_ _0262_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2319_ _0591_ _0597_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1552_ _1130_ _1173_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and3_1
X_1621_ _1206_ _1207_ _1233_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__o31a_1
X_2670_ _0990_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1483_ outputs.divider_buffer\[13\] _1093_ _1111_ outputs.sig_gen.count\[14\] _1120_
+ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__o221ai_1
X_2104_ _0525_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ outputs.div.count\[1\] outputs.div.count\[0\] VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2937_ clknet_leaf_3_clk _0143_ net37 VGND VGND VPWR VPWR outputs.divider_buffer\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2868_ clknet_leaf_26_clk outputs.output_gen.next_count\[5\] net36 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2799_ clknet_leaf_22_clk _0033_ net45 VGND VGND VPWR VPWR outputs.div.a\[12\] sky130_fd_sc_hd__dfrtp_1
X_1819_ _0309_ _0311_ _0299_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2722_ clknet_leaf_32_clk _0020_ net27 VGND VGND VPWR VPWR inputs.octave_fsm.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_2653_ _0978_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
X_2584_ net300 outputs.sig_gen.count\[1\] _0936_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
X_1604_ outputs.divider_buffer\[2\] outputs.shaper.count\[1\] VGND VGND VPWR VPWR
+ _1218_ sky130_fd_sc_hd__or2b_1
X_1535_ _1116_ _1159_ _1161_ _1131_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[11\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1466_ _1103_ outputs.sig_gen.count\[10\] _1092_ outputs.sig_gen.count\[1\] VGND
+ VGND VPWR VPWR _1104_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1397_ _1060_ _1061_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[15\]
+ sky130_fd_sc_hd__nor2_1
X_2018_ outputs.div.q\[18\] _1083_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold183 outputs.signal_buffer2\[15\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 outputs.signal_buffer2\[4\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 outputs.signal_buffer2\[7\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 outputs.output_gen.count\[5\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 inputs.random_update_clock.count\[6\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1320_ _1005_ net15 VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2636_ outputs.shaper.count\[8\] net271 _0966_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2705_ clknet_leaf_37_clk net82 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1449_ _0997_ _1088_ VGND VGND VPWR VPWR outputs.sample_rate.next_count\[6\] sky130_fd_sc_hd__nor2_1
X_2567_ net228 outputs.div.oscillator_out\[11\] _0925_ VGND VGND VPWR VPWR _0934_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1518_ _1149_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_2498_ _0231_ _0534_ _0626_ _0829_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__a41o_1
XFILLER_0_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1303_ _0998_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2283_ _0534_ _0682_ _0688_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2352_ _0626_ _0732_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2421_ _0752_ _0825_ _0247_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1998_ _1002_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_4
X_2619_ outputs.shaper.count\[0\] net237 _0916_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ _0406_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__xnor2_1
X_2970_ clknet_leaf_4_clk _0176_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1852_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1783_ _0280_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2404_ _0809_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_2266_ _0601_ _0598_ _0609_ _0617_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and4_1
X_2335_ _0565_ _0743_ _0555_ _0662_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__o2bb2a_1
X_2197_ _0237_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold87 outputs.sample_rate.next_count\[4\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 outputs.sample_rate.count\[5\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _0068_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 outputs.div.oscillator_out\[16\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 outputs.div.q\[10\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 outputs.div.oscillator_out\[4\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 inputs.random_note_generator.out\[1\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 inputs.random_note_generator.out\[13\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 inputs.keypad_synchronizer.half_sync\[3\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__buf_2
X_2051_ outputs.scaled_buffer\[1\] net105 _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2884_ clknet_leaf_5_clk outputs.sig_gen.next_count\[13\] net42 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[13\] sky130_fd_sc_hd__dfrtp_1
X_1904_ net192 _1004_ outputs.div.next_div _0394_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_1
X_2953_ clknet_leaf_4_clk _0159_ VGND VGND VPWR VPWR outputs.signal_buffer2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_1835_ outputs.div.a\[8\] _0330_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1766_ _0264_ _0267_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__nand2_1
X_1697_ _0216_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2318_ _0576_ _0723_ _0724_ _0726_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__o311a_1
X_2249_ _0556_ _0535_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1551_ outputs.sig_gen.count\[15\] _1172_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_1
X_1482_ _1119_ outputs.sig_gen.count\[6\] outputs.divider_buffer\[16\] _1112_ VGND
+ VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o22a_1
X_1620_ _1200_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2103_ net275 outputs.div.divisor\[10\] _0522_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _0486_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2798_ clknet_leaf_22_clk _0032_ net47 VGND VGND VPWR VPWR outputs.div.a\[11\] sky130_fd_sc_hd__dfrtp_1
X_2936_ clknet_leaf_3_clk _0142_ net37 VGND VGND VPWR VPWR outputs.divider_buffer\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1818_ net185 _1004_ outputs.div.next_div _0316_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__a22o_1
X_2867_ clknet_leaf_26_clk outputs.output_gen.next_count\[4\] net35 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ outputs.div.m\[0\] _0253_ outputs.div.m\[1\] VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a21o_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2652_ outputs.shaper.count\[16\] net207 _1089_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2721_ clknet_leaf_35_clk _0019_ net24 VGND VGND VPWR VPWR inputs.octave_fsm.state\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_14_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2583_ _0942_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_1603_ outputs.shaper.count\[0\] VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__inv_2
X_1465_ outputs.divider_buffer\[10\] VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__inv_2
X_1534_ _1116_ _1159_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ outputs.div.oscillator_out\[10\] _0475_ _0468_ net146 _0478_ VGND VGND VPWR
+ VPWR _0065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ net187 _1058_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2919_ clknet_leaf_1_clk _0125_ VGND VGND VPWR VPWR outputs.div.divisor\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold151 outputs.signal_buffer2\[6\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 outputs.divider_buffer2\[15\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 outputs.div.divisor\[9\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold195 outputs.div.q\[2\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 outputs.signal_buffer2\[11\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 outputs.divider_buffer2\[4\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2635_ _0969_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2704_ clknet_leaf_37_clk inputs.random_note_generator.feedback net22 VGND VGND VPWR
+ VPWR inputs.random_note_generator.out\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1448_ net180 _0996_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor2_1
X_2566_ net244 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1517_ _1130_ _1146_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2497_ _0674_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1379_ inputs.random_update_clock.count\[10\] _1047_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2420_ _0786_ _0824_ _0624_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1302_ outputs.div.count\[3\] outputs.div.count\[4\] _0999_ _1000_ VGND VGND VPWR
+ VPWR _1001_ sky130_fd_sc_hd__a31o_1
X_2282_ _0578_ _0693_ _0603_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o21ai_1
X_2351_ _0617_ _0758_ _0611_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1997_ outputs.div.oscillator_out\[1\] _1090_ _0405_ net136 _0467_ VGND VGND VPWR
+ VPWR _0056_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2618_ _0960_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_2549_ _0924_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1920_ outputs.div.m\[17\] _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ outputs.div.m\[11\] _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2403_ outputs.div.divisor\[8\] _0808_ _0645_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux2_1
X_1782_ outputs.div.a\[3\] _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2265_ _0677_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
X_2334_ _0551_ _0547_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_1
X_2196_ _0607_ _0608_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold22 inputs.keypad_synchronizer.half_sync\[14\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 inputs.keypad_synchronizer.half_sync\[1\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold77 _1087_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 _0071_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0059_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _0057_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 outputs.div.q_out\[5\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 outputs.div.a\[4\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 inputs.key_encoder.octave_key_up VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2050_ _1089_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__buf_4
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2952_ clknet_leaf_4_clk _0158_ VGND VGND VPWR VPWR outputs.signal_buffer2\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2883_ clknet_leaf_5_clk outputs.sig_gen.next_count\[12\] net42 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[12\] sky130_fd_sc_hd__dfrtp_1
X_1903_ _0392_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__xnor2_1
X_1834_ outputs.div.a\[8\] _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
X_1765_ _0249_ _0267_ _0268_ _0252_ net203 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1696_ outputs.div.m\[7\] outputs.div.divisor\[7\] _1294_ VGND VGND VPWR VPWR _0216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2317_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__clkbuf_4
X_2179_ _0591_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
X_2248_ _0650_ _0656_ _0658_ _0660_ _0538_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__o32a_1
XFILLER_0_79_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ outputs.sig_gen.count\[15\] _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__or2_1
X_1481_ outputs.divider_buffer\[6\] VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2033_ _1084_ _1003_ outputs.div.count\[0\] VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_2102_ _0524_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_2935_ clknet_leaf_39_clk _0141_ net26 VGND VGND VPWR VPWR outputs.divider_buffer\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2797_ clknet_leaf_21_clk _0031_ net49 VGND VGND VPWR VPWR outputs.div.a\[10\] sky130_fd_sc_hd__dfrtp_1
X_2866_ clknet_leaf_26_clk outputs.output_gen.next_count\[3\] net35 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1748_ outputs.div.a\[25\] VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
X_1817_ _0314_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _1285_ _1286_ _1287_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__and4b_1
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2651_ _0977_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
X_2582_ net155 outputs.sig_gen.count\[0\] _0936_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__mux2_1
X_1602_ outputs.shaper.count\[1\] outputs.divider_buffer\[2\] VGND VGND VPWR VPWR
+ _1216_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2720_ clknet_leaf_32_clk _0018_ net27 VGND VGND VPWR VPWR inputs.octave_fsm.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1533_ _1160_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
X_1464_ outputs.divider_buffer\[3\] _1099_ outputs.divider_buffer\[9\] _1100_ _1101_
+ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1395_ inputs.random_update_clock.count\[15\] _1058_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and2_1
X_2016_ net134 _1083_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2918_ clknet_leaf_1_clk _0124_ VGND VGND VPWR VPWR outputs.div.divisor\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold152 outputs.signal_buffer2\[16\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold174 _0934_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
X_2849_ clknet_leaf_20_clk _0083_ net48 VGND VGND VPWR VPWR outputs.scaled_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold163 outputs.output_gen.count\[2\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 outputs.div.a\[7\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _0518_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 inputs.random_update_clock.count\[9\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 outputs.divider_buffer2\[3\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2703_ clknet_leaf_14_clk _0017_ net46 VGND VGND VPWR VPWR outputs.div.m\[17\] sky130_fd_sc_hd__dfrtp_2
X_2634_ outputs.shaper.count\[7\] net205 _0966_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__mux2_1
X_2565_ net243 outputs.div.oscillator_out\[10\] _0925_ VGND VGND VPWR VPWR _0933_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1516_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1447_ _0996_ net132 VGND VGND VPWR VPWR outputs.sample_rate.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_49_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1378_ _1047_ _1048_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[9\]
+ sky130_fd_sc_hd__nor2_1
X_2496_ inputs.frequency_lut.rng\[5\] _0892_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1301_ outputs.div.start VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
X_2350_ _0606_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and2_1
X_2281_ _0657_ _0656_ _0689_ _0692_ _0686_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1996_ outputs.div.q\[8\] _0248_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2617_ net159 net301 _0512_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2548_ net188 net225 _0855_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2479_ _0552_ _0657_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ outputs.div.m\[10\] _0321_ _0336_ _0320_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o31a_1
X_1781_ outputs.div.m\[4\] _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__xor2_2
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2402_ _0642_ _0802_ _0803_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2333_ _0569_ _0566_ _0741_ _0686_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2264_ net310 _0676_ _0645_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux2_1
X_2195_ _0594_ _0585_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1979_ outputs.div.a\[24\] _0427_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold45 outputs.sample_rate.count\[0\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_1
Xhold56 outputs.divider_buffer2\[9\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 inputs.keypad_synchronizer.half_sync\[13\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 inputs.random_note_generator.out\[10\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 inputs.random_note_generator.out\[11\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold67 outputs.div.q\[4\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold78 outputs.div.a\[24\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _0092_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2951_ clknet_leaf_5_clk _0157_ VGND VGND VPWR VPWR outputs.signal_buffer2\[8\] sky130_fd_sc_hd__dfxtp_1
X_1902_ _0380_ _0383_ _0378_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2882_ clknet_leaf_3_clk outputs.sig_gen.next_count\[11\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[11\] sky130_fd_sc_hd__dfrtp_1
X_1833_ outputs.div.m\[9\] _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__xor2_1
X_1764_ _0260_ _0266_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1695_ _0215_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
X_2316_ _0567_ _0658_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2178_ inputs.key_encoder.sync_keys\[12\] _0586_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__nor2b_2
X_2247_ _0554_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1480_ outputs.divider_buffer\[7\] _1115_ outputs.divider_buffer\[11\] _1116_ _1117_
+ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2032_ outputs.div.q\[26\] _0252_ _0249_ net264 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__a22o_1
X_2101_ net111 net253 _0522_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2934_ clknet_leaf_2_clk _0140_ net38 VGND VGND VPWR VPWR outputs.divider_buffer\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2865_ clknet_leaf_27_clk outputs.output_gen.next_count\[2\] net49 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2796_ clknet_leaf_22_clk _0030_ net49 VGND VGND VPWR VPWR outputs.div.a\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1747_ _0249_ _0250_ _0251_ _0252_ net140 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__a32o_1
X_1816_ _0301_ _0306_ _0299_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o21a_1
X_1678_ inputs.key_encoder.sync_keys\[12\] _1288_ _1290_ _1291_ VGND VGND VPWR VPWR
+ _1292_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2650_ outputs.shaper.count\[15\] net238 _1089_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__mux2_1
X_2581_ _0941_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
X_1601_ outputs.divider_buffer\[4\] _1213_ _1214_ outputs.divider_buffer\[3\] VGND
+ VGND VPWR VPWR _1215_ sky130_fd_sc_hd__a22o_1
X_1532_ _1130_ _1158_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1463_ outputs.divider_buffer\[4\] outputs.sig_gen.count\[4\] VGND VGND VPWR VPWR
+ _1101_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1394_ _1058_ net167 VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2015_ outputs.div.oscillator_out\[9\] _0475_ _0468_ net134 _0477_ VGND VGND VPWR
+ VPWR _0064_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2848_ clknet_leaf_20_clk _0082_ net48 VGND VGND VPWR VPWR outputs.scaled_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2917_ clknet_leaf_1_clk _0123_ VGND VGND VPWR VPWR outputs.div.divisor\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold175 outputs.signal_buffer2\[17\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ clknet_leaf_16_clk inputs.keypad\[10\] net51 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold142 outputs.div.q\[5\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 outputs.sig_gen.count\[17\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold120 outputs.div.a\[10\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _1073_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 outputs.divider_buffer2\[1\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _0517_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 outputs.div.divisor\[6\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2702_ clknet_leaf_14_clk _0016_ net46 VGND VGND VPWR VPWR outputs.div.m\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2633_ _0968_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
X_2564_ _0932_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1515_ outputs.sig_gen.count\[6\] _1144_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2495_ _0555_ _0657_ _0878_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1446_ outputs.sample_rate.count\[4\] _0995_ net131 VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__a21oi_1
X_1377_ net196 _1046_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ outputs.div.count\[1\] outputs.div.count\[0\] outputs.div.count\[2\] VGND
+ VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2280_ _0552_ _0564_ _0690_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2616_ _0959_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ net155 _1090_ _0405_ outputs.div.q\[8\] _0466_ VGND VGND VPWR VPWR _0055_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2547_ net235 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ outputs.output_gen.count\[6\] _1076_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2478_ _0551_ _0556_ _0543_ _0536_ inputs.frequency_lut.rng\[4\] VGND VGND VPWR VPWR
+ _0878_ sky130_fd_sc_hd__a41o_1
XFILLER_0_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1780_ _0253_ _0281_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2401_ _0230_ _0806_ _0674_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2332_ _0561_ _0706_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2194_ _0595_ _0585_ _0592_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or3b_1
X_2263_ _0534_ _0666_ _0672_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1978_ outputs.div.a\[24\] _0427_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 outputs.sample_rate.count\[2\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 outputs.div.oscillator_out\[14\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 outputs.div.q\[17\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0091_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 outputs.output_gen.count\[0\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
Xhold24 inputs.keypad_synchronizer.half_sync\[6\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 inputs.random_note_generator.out\[8\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1901_ _0390_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nand2_1
X_2950_ clknet_leaf_4_clk _0156_ VGND VGND VPWR VPWR outputs.signal_buffer2\[7\] sky130_fd_sc_hd__dfxtp_1
X_2881_ clknet_leaf_4_clk outputs.sig_gen.next_count\[10\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[10\] sky130_fd_sc_hd__dfrtp_2
X_1832_ outputs.div.m\[8\] _0321_ _0253_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1763_ _0260_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_1
X_1694_ outputs.div.m\[6\] net316 _1294_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2246_ _0535_ _0543_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and2b_1
X_2315_ _0561_ _0659_ _0685_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a21oi_1
X_2177_ _0588_ _0590_ inputs.key_encoder.sync_keys\[11\] inputs.key_encoder.sync_keys\[10\]
+ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a211o_2
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2100_ _0523_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2031_ net159 _0475_ _1003_ outputs.div.q\[25\] _0485_ VGND VGND VPWR VPWR _0072_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2864_ clknet_leaf_21_clk net91 net49 VGND VGND VPWR VPWR outputs.output_gen.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_2795_ clknet_leaf_23_clk _0029_ net45 VGND VGND VPWR VPWR outputs.div.a\[8\] sky130_fd_sc_hd__dfrtp_1
X_2933_ clknet_leaf_39_clk _0139_ net25 VGND VGND VPWR VPWR outputs.divider_buffer\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1815_ _0312_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or2_1
X_1746_ _1003_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1677_ inputs.key_encoder.sync_keys\[4\] inputs.key_encoder.sync_keys\[5\] inputs.key_encoder.sync_keys\[6\]
+ inputs.key_encoder.sync_keys\[7\] VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _0247_ _0625_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2580_ net230 net159 _0936_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__mux2_1
X_1600_ outputs.shaper.count\[2\] VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__inv_2
X_1531_ outputs.sig_gen.count\[10\] _1157_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nand2_1
X_1462_ outputs.sig_gen.count\[9\] VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1393_ inputs.random_update_clock.count\[13\] _1052_ net166 VGND VGND VPWR VPWR _1059_
+ sky130_fd_sc_hd__a21oi_1
X_2014_ net124 _1083_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2847_ clknet_leaf_21_clk _0081_ net48 VGND VGND VPWR VPWR outputs.scaled_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold110 outputs.div.a\[12\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2916_ clknet_leaf_1_clk _0122_ VGND VGND VPWR VPWR outputs.div.divisor\[9\] sky130_fd_sc_hd__dfxtp_1
X_2778_ clknet_leaf_0_clk inputs.keypad\[9\] net25 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold154 outputs.signal_buffer2\[9\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 outputs.div.divisor\[15\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 outputs.div.divisor\[9\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _0515_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 outputs.divider_buffer2\[7\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 inputs.random_update_clock.count\[3\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 inputs.random_update_clock.count\[4\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
Xhold132 inputs.random_update_clock.count\[15\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2632_ outputs.shaper.count\[6\] net206 _0966_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__mux2_1
X_2701_ clknet_leaf_14_clk _0015_ net45 VGND VGND VPWR VPWR outputs.div.m\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1445_ net141 _0995_ VGND VGND VPWR VPWR outputs.sample_rate.next_count\[4\] sky130_fd_sc_hd__xor2_1
XFILLER_0_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2563_ net209 outputs.div.oscillator_out\[9\] _0925_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1514_ outputs.sig_gen.count\[6\] _1144_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2494_ inputs.frequency_lut.rng\[5\] _0709_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ inputs.random_update_clock.count\[9\] inputs.random_update_clock.count\[8\]
+ _1042_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ outputs.div.q\[7\] _0248_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2615_ net109 outputs.sig_gen.count\[16\] _0512_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2546_ net234 outputs.div.oscillator_out\[1\] _0855_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2477_ _0877_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
X_1428_ _1076_ _1077_ VGND VGND VPWR VPWR outputs.output_gen.next_count\[5\] sky130_fd_sc_hd__nor2_1
X_1359_ inputs.random_update_clock.count\[9\] inputs.random_update_clock.count\[11\]
+ inputs.random_update_clock.count\[10\] inputs.random_update_clock.count\[8\] VGND
+ VGND VPWR VPWR _1034_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2400_ _0759_ _0805_ _0624_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2331_ _0738_ _0653_ _0739_ _0575_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a211o_1
X_2262_ _0247_ _0673_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__o21ai_1
X_2193_ _0600_ _0598_ _0606_ _0601_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__o211a_1
X_1977_ _1084_ _0457_ _0458_ _0405_ net133 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2529_ outputs.divider_buffer\[11\] net246 _0905_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold58 _1085_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0069_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 outputs.div.q\[16\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 outputs.output_gen.next_count\[1\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 inputs.keypad_synchronizer.half_sync\[15\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 inputs.keypad_synchronizer.half_sync\[2\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1900_ outputs.div.a\[14\] _0389_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or2_1
X_2880_ clknet_leaf_3_clk outputs.sig_gen.next_count\[9\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[9\] sky130_fd_sc_hd__dfrtp_2
X_1831_ _0327_ _0328_ net161 _1004_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1762_ _0264_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nand2_1
X_1693_ _0214_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2176_ _1289_ _0589_ inputs.key_encoder.sync_keys\[6\] inputs.key_encoder.sync_keys\[7\]
+ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a211o_1
X_2314_ _0572_ _0717_ _0554_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__o21a_1
X_2245_ _0551_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2030_ outputs.div.q\[24\] _1083_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2932_ clknet_leaf_0_clk _0138_ net25 VGND VGND VPWR VPWR outputs.divider_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2863_ clknet_leaf_27_clk outputs.output_gen.next_count\[0\] net35 VGND VGND VPWR
+ VPWR outputs.output_gen.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_1745_ outputs.div.m\[0\] outputs.div.q\[26\] VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or2_1
X_2794_ clknet_leaf_25_clk _0028_ net33 VGND VGND VPWR VPWR outputs.div.a\[7\] sky130_fd_sc_hd__dfrtp_1
X_1814_ _0309_ _0311_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1676_ inputs.key_encoder.sync_keys\[13\] inputs.key_encoder.sync_keys\[1\] inputs.key_encoder.sync_keys\[0\]
+ _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _0556_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__nor2_1
X_2228_ _0603_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1530_ outputs.sig_gen.count\[10\] _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__or2_1
X_1461_ outputs.sig_gen.count\[3\] VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ inputs.random_update_clock.count\[13\] inputs.random_update_clock.count\[14\]
+ _1052_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2013_ outputs.div.oscillator_out\[8\] _0475_ _0468_ net124 _0476_ VGND VGND VPWR
+ VPWR _0063_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ clknet_leaf_1_clk _0121_ VGND VGND VPWR VPWR outputs.div.divisor\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold100 outputs.div.oscillator_out\[0\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 outputs.div.q\[6\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 outputs.signal_buffer2\[2\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
X_2846_ clknet_leaf_20_clk _0080_ net47 VGND VGND VPWR VPWR outputs.scaled_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2777_ clknet_leaf_32_clk inputs.keypad\[8\] net27 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1728_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[0\] VGND VGND VPWR VPWR
+ _0237_ sky130_fd_sc_hd__nor2b_2
Xhold111 inputs.random_update_clock.count\[14\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold122 inputs.random_update_clock.count\[20\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 outputs.signal_buffer2\[13\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 outputs.signal_buffer2\[14\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 outputs.div.q\[3\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 outputs.signal_buffer2\[10\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 outputs.div.oscillator_out\[7\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ outputs.output_gen.count\[4\] _1272_ _1259_ outputs.output_gen.count\[3\]
+ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a22o_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2631_ _0967_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
X_2562_ _0931_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_2700_ clknet_leaf_13_clk _0014_ net45 VGND VGND VPWR VPWR outputs.div.m\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1444_ _0995_ _1086_ VGND VGND VPWR VPWR outputs.sample_rate.next_count\[3\] sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1513_ _1144_ _1145_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[5\] sky130_fd_sc_hd__nor2_1
X_2493_ _0891_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_1375_ _1039_ _1045_ _1046_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2829_ clknet_leaf_6_clk net125 net41 VGND VGND VPWR VPWR outputs.div.q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout50 net54 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1993_ outputs.div.q\[7\] _0252_ _0249_ net199 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2614_ _0958_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2545_ _0922_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2476_ net306 _0876_ _0855_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__mux2_1
X_1427_ net314 _1074_ net227 VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a21oi_1
X_1358_ inputs.random_update_clock.count\[12\] inputs.random_update_clock.count\[15\]
+ inputs.random_update_clock.count\[14\] inputs.random_update_clock.count\[13\] VGND
+ VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2330_ _0568_ _0538_ _0659_ _0663_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a31o_1
X_2192_ _0604_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
X_2261_ _0533_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__buf_2
XFILLER_0_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1976_ _0453_ _0456_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2528_ _0913_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold59 outputs.sample_rate.count\[1\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 outputs.div.oscillator_out\[15\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 outputs.div.oscillator_out\[3\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 inputs.random_note_generator.out\[5\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 inputs.random_note_generator.out\[6\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _0768_ _0858_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1830_ _0318_ _0326_ _1084_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ _0261_ _0263_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__nand2_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1692_ outputs.div.m\[5\] outputs.div.divisor\[5\] _1294_ VGND VGND VPWR VPWR _0214_
+ sky130_fd_sc_hd__mux2_1
X_2313_ _0549_ _0722_ _0569_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2175_ inputs.key_encoder.sync_keys\[4\] inputs.key_encoder.sync_keys\[5\] VGND VGND
+ VPWR VPWR _0589_ sky130_fd_sc_hd__nor2_1
X_2244_ _0556_ inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\] VGND VGND
+ VPWR VPWR _0657_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_75_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1959_ outputs.div.a\[21\] _0427_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2931_ clknet_leaf_0_clk _0137_ net26 VGND VGND VPWR VPWR outputs.divider_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2862_ clknet_leaf_15_clk outputs.div.next_start net50 VGND VGND VPWR VPWR outputs.div.start
+ sky130_fd_sc_hd__dfrtp_1
X_1744_ outputs.div.m\[0\] outputs.div.q\[26\] VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nand2_1
X_1813_ _0309_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nor2_1
X_2793_ clknet_leaf_24_clk _0027_ net32 VGND VGND VPWR VPWR outputs.div.a\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ inputs.key_encoder.sync_keys\[2\] inputs.key_encoder.sync_keys\[3\] VGND VGND
+ VPWR VPWR _1289_ sky130_fd_sc_hd__or2_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2089_ net252 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2158_ _0543_ _0536_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__nor2_1
X_2227_ _0626_ _0634_ _0640_ _0230_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1460_ _1095_ outputs.sig_gen.count\[9\] _1096_ outputs.sig_gen.count\[17\] _1097_
+ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a221o_1
X_1391_ _1057_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2012_ net116 _0248_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2845_ clknet_leaf_22_clk _0079_ net47 VGND VGND VPWR VPWR outputs.scaled_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2914_ clknet_leaf_34_clk _0120_ VGND VGND VPWR VPWR outputs.div.divisor\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold167 outputs.div.a\[21\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold156 outputs.div.count\[4\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 _0055_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _0054_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _0963_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1658_ outputs.scaled_buffer\[4\] _1250_ _1271_ _1246_ _1254_ VGND VGND VPWR VPWR
+ _1272_ sky130_fd_sc_hd__a221oi_2
X_2776_ clknet_leaf_24_clk inputs.keypad\[7\] net32 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1727_ _0231_ _0232_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a21oi_1
Xhold112 _1059_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold123 _1067_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _0937_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _0933_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ outputs.divider_buffer\[12\] _1201_ _1202_ outputs.divider_buffer\[11\] VGND
+ VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a22o_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2630_ outputs.shaper.count\[5\] net215 _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__mux2_1
X_2561_ net271 net277 _0925_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__mux2_1
X_2492_ net220 _0890_ _0855_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__mux2_1
X_1512_ outputs.sig_gen.count\[5\] _1142_ _1131_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1443_ net145 _0994_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1374_ inputs.random_update_clock.count\[8\] _1042_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__and2_1
X_2828_ clknet_leaf_6_clk net117 net41 VGND VGND VPWR VPWR outputs.div.q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2759_ clknet_leaf_25_clk net56 net34 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout51 net54 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout40 net55 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1992_ net199 _0413_ _0249_ net197 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2613_ net103 outputs.sig_gen.count\[15\] _0512_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__mux2_1
X_2544_ net237 net155 _0855_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2475_ _0642_ _0869_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1426_ outputs.output_gen.count\[5\] outputs.output_gen.count\[4\] _1074_ VGND VGND
+ VPWR VPWR _1076_ sky130_fd_sc_hd__and3_1
X_1357_ _1030_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2260_ _0602_ _0629_ _0633_ _0638_ _0238_ _0626_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux4_1
X_2191_ _0600_ _0593_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1975_ _0453_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold38 _0058_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2527_ outputs.divider_buffer\[10\] net275 _0905_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
Xhold27 inputs.random_note_generator.out\[0\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 inputs.random_note_generator.out\[7\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ inputs.random_update_clock.count\[21\] _1066_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or2_1
X_2458_ _0576_ _0569_ _0799_ _0859_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR
+ _0860_ sky130_fd_sc_hd__a311o_1
Xhold49 _0070_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _0552_ _0559_ _0564_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1760_ _0261_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__or2_1
X_1691_ _0213_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _0539_ _0541_ _0535_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2174_ inputs.key_encoder.sync_keys\[8\] inputs.key_encoder.sync_keys\[9\] VGND VGND
+ VPWR VPWR _0588_ sky130_fd_sc_hd__nor2_1
X_2243_ inputs.frequency_lut.rng\[0\] inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\]
+ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1958_ _0440_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__nand2_1
X_1889_ _0370_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2861_ clknet_leaf_17_clk outputs.div.next_div net54 VGND VGND VPWR VPWR outputs.div.div
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2930_ clknet_leaf_0_clk _0136_ net26 VGND VGND VPWR VPWR outputs.divider_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1743_ _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_4
X_1812_ outputs.div.m\[7\] _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__xnor2_1
X_2792_ clknet_leaf_25_clk _0026_ net32 VGND VGND VPWR VPWR outputs.div.a\[5\] sky130_fd_sc_hd__dfrtp_1
X_1674_ inputs.key_encoder.sync_keys\[11\] inputs.key_encoder.sync_keys\[8\] inputs.key_encoder.sync_keys\[9\]
+ inputs.key_encoder.sync_keys\[10\] VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__or4_4
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _0611_ _0638_ _0639_ _0624_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a211o_1
X_2088_ net251 outputs.div.divisor\[3\] _0513_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_1
X_2157_ _0562_ _0566_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _1043_ _1055_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2011_ _1089_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2844_ clknet_leaf_16_clk _0078_ net50 VGND VGND VPWR VPWR outputs.div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2913_ clknet_leaf_34_clk _0119_ VGND VGND VPWR VPWR outputs.div.divisor\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold146 outputs.div.q_out\[2\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 outputs.signal_buffer2\[12\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 outputs.signal_buffer2\[1\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ outputs.shaper.count\[10\] VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__inv_2
X_1657_ outputs.scaled_buffer\[3\] _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__xor2_1
Xhold124 outputs.div.a\[11\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ clknet_leaf_0_clk inputs.keypad\[6\] net25 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold157 inputs.random_update_clock.count\[7\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 inputs.random_update_clock.count\[0\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
X_1726_ _0233_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or2b_1
Xhold113 inputs.random_update_clock.count\[16\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold135 inputs.random_update_clock.count\[19\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\]
+ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1442_ _0994_ net113 VGND VGND VPWR VPWR outputs.sample_rate.next_count\[2\] sky130_fd_sc_hd__nor2_1
X_2560_ _0930_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
X_1511_ outputs.sig_gen.count\[4\] outputs.sig_gen.count\[5\] _1138_ VGND VGND VPWR
+ VPWR _1144_ sky130_fd_sc_hd__and3_1
X_2491_ _0231_ _0534_ _0851_ _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1373_ inputs.random_update_clock.count\[8\] _1042_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_1
X_2827_ clknet_leaf_6_clk net108 net41 VGND VGND VPWR VPWR outputs.div.q\[14\] sky130_fd_sc_hd__dfrtp_1
X_2758_ clknet_leaf_33_clk net79 net32 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1709_ outputs.div.m\[13\] outputs.div.divisor\[13\] _0218_ VGND VGND VPWR VPWR _0223_
+ sky130_fd_sc_hd__mux2_1
X_2689_ clknet_leaf_23_clk _0003_ net33 VGND VGND VPWR VPWR outputs.div.m\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2612_ _0957_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ net197 _0413_ _0249_ net122 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2543_ _0921_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_1425_ net236 _1074_ VGND VGND VPWR VPWR outputs.output_gen.next_count\[4\] sky130_fd_sc_hd__xor2_1
X_2474_ _0727_ _0870_ _0874_ _0674_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__a211o_1
X_1356_ inputs.random_update_clock.count\[1\] inputs.random_update_clock.count\[0\]
+ inputs.random_update_clock.count\[3\] inputs.random_update_clock.count\[2\] VGND
+ VGND VPWR VPWR _1031_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2190_ _0603_ _0587_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or2_1
X_1974_ _0454_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2526_ _0912_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_2388_ _0568_ _0549_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nor2_1
Xhold39 inputs.key_encoder.sync_keys\[15\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 inputs.random_note_generator.out\[14\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 inputs.random_note_generator.out\[4\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2457_ _0685_ _0745_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nor2_1
X_1408_ _1066_ net178 VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1339_ _1021_ VGND VGND VPWR VPWR inputs.keypad\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ outputs.div.m\[4\] outputs.div.divisor\[4\] _1294_ VGND VGND VPWR VPWR _0213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _0716_ _0719_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o21a_1
X_2242_ _0561_ _0549_ _0650_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2173_ inputs.key_encoder.sync_keys\[12\] _1288_ _1291_ _0586_ VGND VGND VPWR VPWR
+ _0587_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ _0433_ _0436_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1888_ _0378_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2509_ _0903_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2860_ clknet_leaf_20_clk net172 net47 VGND VGND VPWR VPWR outputs.div.q_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1811_ outputs.div.m\[6\] _0281_ _0296_ _0253_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__o31a_1
X_2791_ clknet_leaf_25_clk _0025_ net34 VGND VGND VPWR VPWR outputs.div.a\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1742_ _1082_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__buf_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1673_ inputs.key_encoder.sync_keys\[14\] inputs.key_encoder.sync_keys\[15\] inputs.key_encoder.octave_key_up
+ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__nor3_2
XFILLER_0_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2225_ _0607_ _0609_ _0614_ _0611_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a31oi_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
X_2087_ net280 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_2156_ _0564_ _0567_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2989_ clknet_leaf_4_clk _0195_ net40 VGND VGND VPWR VPWR outputs.shaper.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2010_ outputs.div.oscillator_out\[7\] _1090_ _0468_ net116 _0474_ VGND VGND VPWR
+ VPWR _0062_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2912_ clknet_leaf_34_clk _0118_ VGND VGND VPWR VPWR outputs.div.divisor\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2843_ clknet_leaf_16_clk _0077_ net50 VGND VGND VPWR VPWR outputs.div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2774_ clknet_leaf_25_clk inputs.keypad\[5\] net34 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ inputs.octave_fsm.octave_key_up inputs.down.det_edge VGND VGND VPWR VPWR _0234_
+ sky130_fd_sc_hd__or2b_1
Xhold125 outputs.sample_rate.count\[6\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
Xhold158 outputs.div.q\[1\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _0089_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 outputs.div.a\[16\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ outputs.shaper.count\[11\] VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__inv_2
X_1656_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] outputs.scaled_buffer\[2\]
+ net21 VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__o31a_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold169 outputs.divider_buffer2\[6\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 outputs.div.a\[6\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 inputs.random_update_clock.count\[11\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0545_ _0550_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_1
X_2208_ _0615_ _0621_ _0238_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1441_ outputs.sample_rate.count\[1\] outputs.sample_rate.count\[0\] net112 VGND
+ VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1510_ _1142_ _1143_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[4\] sky130_fd_sc_hd__nor2_1
X_2490_ _0886_ _0888_ _0603_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1372_ _1042_ _1044_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2826_ clknet_leaf_7_clk net151 net41 VGND VGND VPWR VPWR outputs.div.q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1708_ _0222_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_2688_ clknet_leaf_34_clk _0002_ net33 VGND VGND VPWR VPWR outputs.div.m\[2\] sky130_fd_sc_hd__dfrtp_1
X_2757_ clknet_leaf_28_clk net57 net34 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1639_ outputs.scaled_buffer\[6\] _1247_ _1252_ outputs.scaled_buffer\[7\] VGND VGND
+ VPWR VPWR _1253_ sky130_fd_sc_hd__or4b_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout42 net55 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xfanout53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xfanout31 net36 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1990_ net122 _0413_ _0249_ net210 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a22o_1
X_2611_ net101 outputs.sig_gen.count\[14\] _0947_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2542_ outputs.divider_buffer\[17\] net248 _0916_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1424_ _1074_ _1075_ VGND VGND VPWR VPWR outputs.output_gen.next_count\[3\] sky130_fd_sc_hd__nor2_1
X_1355_ inputs.random_update_clock.count\[4\] inputs.random_update_clock.count\[6\]
+ inputs.random_update_clock.count\[7\] inputs.random_update_clock.count\[5\] VGND
+ VGND VPWR VPWR _1030_ sky130_fd_sc_hd__or4bb_1
X_2473_ _0871_ _0873_ _0727_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2809_ clknet_leaf_17_clk _0043_ net51 VGND VGND VPWR VPWR outputs.div.a\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1973_ outputs.div.a\[23\] _0427_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2525_ outputs.divider_buffer\[9\] net111 _0905_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1338_ net1 net7 VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__and2b_1
X_2387_ _0724_ _0792_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or2_1
Xhold18 inputs.random_note_generator.out\[3\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 inputs.random_note_generator.out\[2\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ inputs.random_update_clock.count\[19\] _1065_ net177 VGND VGND VPWR VPWR _1067_
+ sky130_fd_sc_hd__a21oi_1
X_2456_ _0542_ _0648_ _0857_ _0562_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2310_ _0716_ _0719_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__a21oi_1
X_2172_ inputs.key_encoder.sync_keys\[13\] _1287_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__and2b_1
X_2241_ _0561_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__nand2_1
X_1956_ _0402_ _0426_ _0428_ _0429_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o211ai_1
X_1887_ _0375_ _0377_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2508_ outputs.divider_buffer\[1\] net241 _0497_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__mux2_1
X_2439_ _0842_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2790_ clknet_leaf_26_clk _0024_ net35 VGND VGND VPWR VPWR outputs.div.a\[3\] sky130_fd_sc_hd__dfrtp_1
X_1810_ outputs.div.a\[6\] VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1741_ _0234_ _0247_ _0243_ _0233_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1672_ outputs.output_gen.count\[7\] _1283_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__clkbuf_4
X_2224_ _0635_ _0637_ _0616_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2086_ outputs.divider_buffer2\[2\] net279 _0513_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1939_ net295 _0413_ outputs.div.next_div _0425_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a22o_1
X_2988_ clknet_leaf_4_clk _0194_ net40 VGND VGND VPWR VPWR outputs.shaper.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2911_ clknet_leaf_34_clk _0117_ VGND VGND VPWR VPWR outputs.div.divisor\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold115 outputs.div.a\[23\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 outputs.div.oscillator_out\[17\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
X_2842_ clknet_leaf_16_clk _0076_ net51 VGND VGND VPWR VPWR outputs.div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold126 outputs.div.a\[1\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
X_2773_ clknet_leaf_33_clk inputs.keypad\[4\] net32 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1724_ inputs.down.det_edge inputs.octave_fsm.octave_key_up VGND VGND VPWR VPWR _0233_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold159 _0049_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 outputs.div.a\[15\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ _1111_ outputs.shaper.count\[13\] _1199_ outputs.divider_buffer\[13\] VGND
+ VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a2bb2o_1
X_1655_ outputs.output_gen.count\[3\] _1259_ _1263_ outputs.output_gen.count\[2\]
+ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__o221a_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold148 outputs.div.a\[2\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2069_ outputs.div.q\[1\] outputs.div.q\[0\] _0507_ _0508_ VGND VGND VPWR VPWR _0509_
+ sky130_fd_sc_hd__or4_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2138_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__clkbuf_4
X_2207_ _0618_ _0619_ _0620_ _0604_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or4b_1
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440_ net114 net100 VGND VGND VPWR VPWR outputs.sample_rate.next_count\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1371_ net212 _1040_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__o21ai_1
X_2825_ clknet_leaf_9_clk net99 net43 VGND VGND VPWR VPWR outputs.div.q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1638_ outputs.scaled_buffer\[5\] outputs.scaled_buffer\[4\] _1188_ VGND VGND VPWR
+ VPWR _1252_ sky130_fd_sc_hd__or3_1
X_1707_ outputs.div.m\[12\] net276 _0218_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
X_2687_ clknet_leaf_34_clk _0001_ net33 VGND VGND VPWR VPWR outputs.div.m\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2756_ clknet_leaf_33_clk net61 net32 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1569_ _1185_ VGND VGND VPWR VPWR inputs.mode_edge.ff_in sky130_fd_sc_hd__inv_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout54 net55 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout32 net36 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2610_ _0956_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_2541_ _0920_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2472_ _0650_ _0745_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__o21ai_1
X_1423_ net268 _1072_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__nor2_1
X_1354_ inputs.random_update_clock.count\[4\] inputs.random_update_clock.count\[5\]
+ _1026_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__and3_1
X_2808_ clknet_leaf_17_clk _0042_ net51 VGND VGND VPWR VPWR outputs.div.a\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2739_ clknet_leaf_31_clk inputs.random_update_clock.next_count\[16\] net29 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1972_ outputs.div.a\[23\] _0427_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2524_ _0911_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2455_ _0652_ _0817_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and2_1
X_1337_ _1020_ VGND VGND VPWR VPWR inputs.keypad\[14\] sky130_fd_sc_hd__clkbuf_1
Xhold19 inputs.keypad_synchronizer.half_sync\[16\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ inputs.random_update_clock.count\[19\] inputs.random_update_clock.count\[20\]
+ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and3_1
X_2386_ _0722_ _0764_ _0551_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2171_ inputs.key_encoder.sync_keys\[10\] _0584_ inputs.key_encoder.sync_keys\[11\]
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__o21bai_4
X_2240_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1955_ outputs.div.a\[20\] outputs.div.a\[19\] _0427_ VGND VGND VPWR VPWR _0439_
+ sky130_fd_sc_hd__o21ai_1
X_1886_ _0375_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2507_ _0902_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_2438_ outputs.div.divisor\[10\] _0841_ _0645_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2369_ _0536_ _0540_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__and2_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1671_ _1275_ _1279_ _1283_ outputs.output_gen.count\[7\] _1284_ VGND VGND VPWR VPWR
+ _1285_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1740_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ net242 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
X_2154_ inputs.frequency_lut.rng\[3\] VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_4
X_2223_ _0596_ _0591_ _0592_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2987_ clknet_leaf_4_clk _0193_ net37 VGND VGND VPWR VPWR outputs.shaper.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1938_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__xnor2_1
X_1869_ _0353_ _0348_ _0349_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2841_ clknet_leaf_16_clk _0075_ net51 VGND VGND VPWR VPWR outputs.div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ clknet_leaf_34_clk _0116_ VGND VGND VPWR VPWR outputs.div.divisor\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold105 _0072_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 outputs.sample_rate.count\[7\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 outputs.div.q_out\[7\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 outputs.div.a\[13\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold138 outputs.sig_gen.count\[0\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ outputs.output_gen.count\[2\] _1263_ _1265_ _1267_ VGND VGND VPWR VPWR _1268_
+ sky130_fd_sc_hd__a22o_1
X_1723_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\] VGND VGND VPWR VPWR
+ _0232_ sky130_fd_sc_hd__or2b_1
X_2772_ clknet_leaf_32_clk inputs.keypad\[3\] net27 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1585_ outputs.shaper.count\[12\] VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__inv_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2206_ _0585_ _0598_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2068_ outputs.div.q\[3\] outputs.div.q\[2\] outputs.div.q\[5\] outputs.div.q\[4\]
+ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2137_ inputs.frequency_lut.rng\[3\] VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1032_ _1035_ _1036_ _1037_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__nand4_2
X_2824_ clknet_leaf_9_clk net93 net44 VGND VGND VPWR VPWR outputs.div.q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1637_ inputs.wavetype_fsm.state\[0\] inputs.wavetype_fsm.state\[1\] VGND VGND VPWR
+ VPWR _1251_ sky130_fd_sc_hd__nand2_1
X_1706_ _0221_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2686_ clknet_leaf_23_clk _0000_ net32 VGND VGND VPWR VPWR outputs.div.m\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2755_ clknet_leaf_32_clk net65 net28 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1499_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] outputs.sig_gen.count\[2\]
+ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1568_ net115 inputs.key_encoder.mode_key VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or2b_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout44 net55 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_4
Xfanout55 net19 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xfanout33 net36 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xfanout22 net24 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2540_ outputs.divider_buffer\[16\] net266 _0916_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1422_ outputs.output_gen.count\[3\] _1072_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ _0568_ _0557_ _0575_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__a21oi_1
X_1353_ inputs.random_update_clock.count\[4\] _1026_ net293 VGND VGND VPWR VPWR _1028_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2807_ clknet_leaf_17_clk _0041_ net53 VGND VGND VPWR VPWR outputs.div.a\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2738_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[15\] net30 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2669_ _0989_ _0562_ _0983_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1971_ _0440_ _0441_ _0451_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2454_ _0856_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
X_2523_ outputs.divider_buffer\[8\] net245 _0905_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__mux2_1
X_2385_ _0791_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1405_ net190 _1065_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[19\]
+ sky130_fd_sc_hd__xor2_1
Xinput1 cs VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_1336_ net1 net6 VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2170_ inputs.key_encoder.sync_keys\[8\] _0583_ inputs.key_encoder.sync_keys\[9\]
+ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__o21ba_1
X_1954_ _0277_ _0437_ _0438_ _0405_ net222 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ outputs.div.m\[14\] _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2506_ outputs.divider_buffer\[0\] net255 _0497_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux2_1
X_2368_ net208 _0513_ _0763_ _0775_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__o22a_1
X_2437_ _0534_ _0831_ _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__a21o_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1011_ VGND VGND VPWR VPWR inputs.keypad\[5\] sky130_fd_sc_hd__clkbuf_1
X_2299_ _0650_ _0656_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__nor3_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1670_ outputs.output_gen.count\[6\] _1278_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2222_ _0609_ _0631_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand2_1
X_2084_ net241 outputs.div.divisor\[1\] _0513_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_1
X_2153_ _0537_ _0540_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1937_ _0417_ _0421_ _0415_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o21ai_1
X_2986_ clknet_leaf_5_clk _0192_ net37 VGND VGND VPWR VPWR outputs.shaper.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1868_ _0360_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nand2_1
X_1799_ _0295_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2840_ clknet_leaf_16_clk _0074_ net51 VGND VGND VPWR VPWR outputs.div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2771_ clknet_leaf_32_clk inputs.keypad\[2\] net28 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold117 _0094_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _1095_ outputs.shaper.count\[8\] _1197_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a21o_1
Xhold106 outputs.div.a\[8\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ outputs.output_gen.count\[1\] _1264_ _1266_ outputs.output_gen.count\[0\]
+ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__a211o_1
Xhold128 inputs.wavetype_fsm.state\[1\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_4
Xhold139 inputs.random_update_clock.count\[2\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2205_ _0591_ _0608_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2067_ outputs.div.q\[7\] outputs.div.q\[6\] outputs.div.q\[8\] VGND VGND VPWR VPWR
+ _0507_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2136_ _0547_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2969_ clknet_leaf_5_clk _0175_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2823_ clknet_leaf_10_clk net121 net44 VGND VGND VPWR VPWR outputs.div.q\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1705_ outputs.div.m\[11\] net278 _0218_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2754_ clknet_leaf_32_clk net69 net28 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1636_ _1249_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2685_ clknet_leaf_26_clk net184 net35 VGND VGND VPWR VPWR inputs.wavetype_fsm.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1567_ _1183_ _1184_ VGND VGND VPWR VPWR inputs.random_note_generator.feedback sky130_fd_sc_hd__xnor2_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1134_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_2119_ inputs.key_encoder.sync_keys\[13\] _1287_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__nand2_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout45 net55 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xfanout23 net24 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XFILLER_0_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ _1072_ net219 VGND VGND VPWR VPWR outputs.output_gen.next_count\[2\] sky130_fd_sc_hd__nor2_1
X_2470_ _0555_ _0550_ _0810_ _0576_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__o211ai_1
X_1352_ net176 _1026_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2806_ clknet_leaf_18_clk _0040_ net53 VGND VGND VPWR VPWR outputs.div.a\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2668_ _0537_ _1182_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__xor2_1
X_2737_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[14\] net30 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_2599_ net277 outputs.sig_gen.count\[8\] _0947_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__mux2_1
X_1619_ _1197_ _1232_ _1203_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1970_ outputs.div.a\[22\] outputs.div.a\[21\] outputs.div.a\[20\] outputs.div.a\[19\]
+ _0427_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o41a_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2522_ _0910_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2453_ outputs.div.divisor\[11\] _0854_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__mux2_1
X_2384_ outputs.div.divisor\[7\] _0790_ _0645_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1404_ _1039_ _1064_ _1065_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[18\]
+ sky130_fd_sc_hd__nor3_1
X_1335_ _1019_ VGND VGND VPWR VPWR inputs.keypad\[13\] sky130_fd_sc_hd__clkbuf_1
Xinput2 gpio[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1953_ _0431_ _0435_ _0436_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21o_1
X_1884_ outputs.div.m\[13\] outputs.div.m\[12\] _0357_ _0320_ VGND VGND VPWR VPWR
+ _0376_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2505_ _0901_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2367_ _0770_ _0774_ _0513_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a21bo_1
X_1318_ _1005_ net14 VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and2b_1
X_2436_ _0674_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__nor2_1
X_2298_ _0538_ _0707_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__and2_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _0564_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nand2_1
X_2221_ _0601_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2083_ _0514_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1936_ outputs.div.a\[18\] _0414_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__xnor2_2
X_2985_ clknet_leaf_7_clk _0191_ net42 VGND VGND VPWR VPWR outputs.shaper.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1867_ _0356_ _0359_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1798_ outputs.div.m\[6\] _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__xnor2_1
X_2419_ _0611_ _0804_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2770_ clknet_leaf_32_clk inputs.keypad\[1\] net27 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1721_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold107 outputs.div.count\[2\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ _1095_ outputs.shaper.count\[8\] outputs.divider_buffer\[10\] _1196_ VGND
+ VGND VPWR VPWR _1197_ sky130_fd_sc_hd__a2bb2o_1
X_1652_ outputs.scaled_buffer\[0\] _1250_ _1254_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__a21oi_1
Xhold129 inputs.wavetype_fsm.next_state\[1\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 outputs.div.a\[5\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__buf_2
X_2204_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2066_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1919_ _0320_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and2_1
X_2968_ clknet_leaf_4_clk _0174_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2899_ clknet_leaf_0_clk _0105_ VGND VGND VPWR VPWR outputs.divider_buffer2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2822_ clknet_leaf_10_clk net137 net50 VGND VGND VPWR VPWR outputs.div.q\[9\] sky130_fd_sc_hd__dfrtp_1
X_1704_ _0220_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2684_ clknet_leaf_26_clk inputs.wavetype_fsm.next_state\[0\] net35 VGND VGND VPWR
+ VPWR inputs.wavetype_fsm.state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2753_ clknet_leaf_32_clk net66 net27 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1497_ _1131_ _1132_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__and3_1
X_1635_ inputs.wavetype_fsm.state\[0\] inputs.wavetype_fsm.state\[1\] VGND VGND VPWR
+ VPWR _1249_ sky130_fd_sc_hd__and2b_1
X_1566_ net319 inputs.random_note_generator.out\[10\] VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__xor2_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2049_ _0496_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
X_2118_ _0532_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout46 net55 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout24 net19 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1420_ outputs.output_gen.count\[1\] net90 net218 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__a21oi_1
X_1351_ _1026_ _1027_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_2805_ clknet_leaf_18_clk _0039_ net53 VGND VGND VPWR VPWR outputs.div.a\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1618_ _1204_ _1205_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__nor2_1
X_2667_ _0988_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2736_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[13\] net31 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[13\] sky130_fd_sc_hd__dfrtp_1
X_1549_ _1170_ _1168_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nor2_1
X_2598_ _0950_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2521_ outputs.divider_buffer\[7\] net231 _0905_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2452_ _0512_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__buf_4
X_1403_ inputs.random_update_clock.count\[18\] _1063_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2_1
X_2383_ _0783_ _0789_ _0674_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux2_1
X_1334_ net1 net9 VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__and2b_1
Xinput3 gpio[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_2719_ clknet_leaf_37_clk net72 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ _0431_ _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nand3_1
X_1883_ outputs.div.a\[13\] VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2504_ outputs.div.divisor\[17\] _0900_ _0855_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux2_1
X_2435_ _0836_ _0838_ _0578_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ _1010_ VGND VGND VPWR VPWR inputs.keypad\[4\] sky130_fd_sc_hd__buf_1
X_2366_ _0578_ _0773_ _0534_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a21oi_1
X_2297_ _0651_ _0663_ _0706_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_66_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2082_ net255 net317 _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
X_2151_ _0536_ _0542_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
X_2220_ _0629_ _0633_ _0238_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux2_1
X_2984_ clknet_leaf_8_clk _0190_ net43 VGND VGND VPWR VPWR outputs.shaper.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1935_ net256 _0413_ outputs.div.next_div _0422_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1866_ _0356_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or2_1
X_1797_ _0281_ _0296_ _0253_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2418_ _0585_ _0594_ _0606_ _0601_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__o211a_2
X_2349_ _0613_ _0605_ _0627_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 outputs.div.q_out\[3\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ outputs.output_gen.count\[1\] _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__or2_1
X_1720_ inputs.octave_fsm.state\[2\] _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__nand2_1
X_1582_ outputs.shaper.count\[9\] VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__inv_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold119 inputs.random_update_clock.count\[1\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
X_2065_ outputs.div.div _0998_ _1001_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and3_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2134_ inputs.frequency_lut.rng\[2\] _0539_ _0541_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and3_1
X_2203_ _0599_ _0614_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2967_ clknet_leaf_5_clk _0173_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1918_ outputs.div.m\[16\] outputs.div.m\[15\] _0386_ VGND VGND VPWR VPWR _0407_
+ sky130_fd_sc_hd__or3_1
X_1849_ _0277_ _0343_ _0344_ _0252_ net175 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a32o_1
X_2898_ clknet_leaf_1_clk _0104_ VGND VGND VPWR VPWR outputs.divider_buffer2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2821_ clknet_leaf_15_clk net156 net50 VGND VGND VPWR VPWR outputs.div.q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2683_ clknet_leaf_9_clk outputs.sample_rate.next_count\[7\] net55 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[7\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
X_1634_ outputs.scaled_buffer\[4\] _1188_ net21 _1247_ VGND VGND VPWR VPWR _1248_
+ sky130_fd_sc_hd__a31o_1
X_1703_ outputs.div.m\[10\] outputs.div.divisor\[10\] _0218_ VGND VGND VPWR VPWR _0220_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2752_ clknet_leaf_28_clk net58 net34 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1496_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] VGND VGND VPWR VPWR
+ _1133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1182_ inputs.random_note_generator.out\[13\] VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__xor2_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2048_ outputs.scaled_buffer\[0\] net129 _0218_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
X_2117_ net248 outputs.div.divisor\[17\] _0522_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout47 net49 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xfanout25 net26 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xfanout36 net19 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ net198 _1024_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
X_2804_ clknet_leaf_18_clk _0038_ net52 VGND VGND VPWR VPWR outputs.div.a\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1617_ _1210_ _1212_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__and3b_1
X_2597_ net221 outputs.sig_gen.count\[7\] _0947_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2666_ _0987_ _0537_ _0983_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__mux2_1
X_2735_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[12\] net30 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[12\] sky130_fd_sc_hd__dfrtp_1
X_1548_ _1170_ _1168_ _1171_ _1131_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[14\]
+ sky130_fd_sc_hd__o211a_1
X_1479_ outputs.divider_buffer\[8\] outputs.sig_gen.count\[8\] VGND VGND VPWR VPWR
+ _1117_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2520_ _0909_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
X_2451_ _0534_ _0849_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ net307 _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1333_ _1018_ VGND VGND VPWR VPWR inputs.keypad\[12\] sky130_fd_sc_hd__clkbuf_1
X_3003_ clknet_leaf_28_clk net62 net35 VGND VGND VPWR VPWR outputs.pwm_output sky130_fd_sc_hd__dfrtp_1
Xinput4 gpio[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_2382_ _0247_ _0787_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2718_ clknet_leaf_37_clk net87 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2649_ _0976_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ outputs.div.a\[20\] _0427_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__xnor2_1
X_1882_ net182 _1004_ outputs.div.next_div _0374_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2365_ _0768_ _0660_ _0771_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a31o_1
X_2434_ _0685_ _0648_ _0837_ _0725_ _0718_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2503_ _0898_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nand2_1
X_1316_ _1005_ net13 VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__and2b_1
X_2296_ _0554_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2081_ _0512_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__clkbuf_4
X_2150_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_4
X_1934_ _0417_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__xor2_1
X_2983_ clknet_leaf_10_clk _0189_ net44 VGND VGND VPWR VPWR outputs.shaper.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1865_ outputs.div.m\[12\] _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__xor2_1
X_1796_ outputs.div.m\[5\] outputs.div.m\[4\] VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2417_ _0576_ _0819_ _0821_ _0674_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a31o_1
X_2348_ _0585_ _0593_ _0597_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o21a_1
X_2279_ _0568_ _0541_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold109 _0090_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ _1191_ _1193_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__or3b_1
XFILLER_0_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1650_ outputs.scaled_buffer\[0\] _1246_ _1250_ outputs.scaled_buffer\[1\] _1254_
+ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__a221oi_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2202_ _0595_ _0591_ _0600_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_2
X_2064_ _0504_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2133_ _0535_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2966_ clknet_leaf_7_clk _0172_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_1917_ outputs.div.a\[16\] VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__inv_2
X_2897_ clknet_leaf_0_clk _0103_ VGND VGND VPWR VPWR outputs.divider_buffer2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1848_ _0339_ _0342_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1779_ outputs.div.m\[3\] outputs.div.m\[2\] outputs.div.m\[0\] outputs.div.m\[1\]
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or4_2
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2820_ clknet_leaf_20_clk net200 net52 VGND VGND VPWR VPWR outputs.div.q\[7\] sky130_fd_sc_hd__dfrtp_2
X_2751_ clknet_leaf_30_clk inputs.up.ff_in net27 VGND VGND VPWR VPWR inputs.octave_fsm.octave_key_up
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2682_ clknet_leaf_9_clk outputs.sample_rate.next_count\[6\] net43 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[6\] sky130_fd_sc_hd__dfrtp_1
X_1633_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__inv_2
X_1702_ _0219_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1564_ inputs.random_note_generator.out\[15\] VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__buf_2
X_1495_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] VGND VGND VPWR VPWR
+ _1132_ sky130_fd_sc_hd__or2_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2047_ _0495_ _0492_ _1090_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout37 net40 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
X_2116_ net267 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
Xfanout26 net19 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
X_2949_ clknet_leaf_5_clk _0155_ VGND VGND VPWR VPWR outputs.signal_buffer2\[6\] sky130_fd_sc_hd__dfxtp_1
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2803_ clknet_leaf_15_clk _0037_ net50 VGND VGND VPWR VPWR outputs.div.a\[16\] sky130_fd_sc_hd__dfrtp_1
X_2734_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[11\] net30 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2596_ _0949_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
X_1547_ _1170_ _1168_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__nand2_1
X_1616_ _1226_ _1227_ _1228_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__a31o_1
X_2665_ _0543_ _1182_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__xor2_1
X_1478_ outputs.sig_gen.count\[11\] VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2450_ _0230_ _0787_ _0852_ _0642_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__a211o_1
X_1401_ _1039_ net285 _1063_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[17\]
+ sky130_fd_sc_hd__nor3_1
X_2381_ _0229_ _0700_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 gpio[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1332_ net1 net5 VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__and2b_1
X_3002_ clknet_leaf_35_clk _0208_ net24 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[5\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2717_ clknet_leaf_37_clk net85 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2648_ net273 net254 _0966_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__mux2_1
X_2579_ _0940_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ _0277_ _0434_ _0435_ _0405_ net281 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a32o_1
X_1881_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2502_ _0727_ _0768_ _0533_ _0862_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__or4_1
X_2364_ _0562_ _0557_ _0567_ _0717_ _0768_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a311oi_1
X_1315_ _1009_ VGND VGND VPWR VPWR inputs.keypad\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2433_ _0547_ _0776_ _0555_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__o21ai_1
X_2295_ inputs.frequency_lut.rng\[1\] inputs.frequency_lut.rng\[2\] VGND VGND VPWR
+ VPWR _0706_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2080_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1933_ _0402_ _0418_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__o21ba_1
X_2982_ clknet_leaf_10_clk _0188_ net44 VGND VGND VPWR VPWR outputs.shaper.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1864_ _0320_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__nand2_1
X_1795_ outputs.div.a\[5\] VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2347_ _0755_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
X_2416_ _0562_ _0564_ _0820_ _0727_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__o211ai_1
X_2278_ _0538_ _0536_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1580_ _1192_ outputs.shaper.count\[15\] VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2132_ _0538_ inputs.frequency_lut.rng\[1\] VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and2_1
X_2201_ _0601_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and2_1
X_2063_ net303 net171 _0497_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2965_ clknet_leaf_8_clk _0171_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_1916_ _0277_ _0403_ _0404_ _0405_ net158 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1847_ _0339_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or2_1
X_2896_ clknet_leaf_0_clk _0102_ VGND VGND VPWR VPWR outputs.divider_buffer2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_1778_ _0273_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2681_ clknet_leaf_9_clk outputs.sample_rate.next_count\[5\] net43 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1701_ outputs.div.m\[9\] net217 _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2750_ clknet_leaf_31_clk net88 net31 VGND VGND VPWR VPWR inputs.up.ff_out sky130_fd_sc_hd__dfrtp_1
X_1494_ net193 _1131_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[0\] sky130_fd_sc_hd__nand2_1
X_1632_ inputs.wavetype_fsm.state\[1\] inputs.wavetype_fsm.state\[0\] VGND VGND VPWR
+ VPWR _1246_ sky130_fd_sc_hd__nor2b_4
X_1563_ net183 _1179_ VGND VGND VPWR VPWR inputs.wavetype_fsm.next_state\[1\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2115_ net266 outputs.div.divisor\[16\] _0522_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux2_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2046_ net211 VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__inv_2
Xfanout49 net55 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
Xfanout38 net40 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2948_ clknet_leaf_8_clk _0154_ VGND VGND VPWR VPWR outputs.signal_buffer2\[5\] sky130_fd_sc_hd__dfxtp_1
X_2879_ clknet_leaf_3_clk outputs.sig_gen.next_count\[8\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2802_ clknet_leaf_20_clk _0036_ net47 VGND VGND VPWR VPWR outputs.div.a\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2733_ clknet_leaf_29_clk inputs.random_update_clock.next_count\[10\] net30 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[10\] sky130_fd_sc_hd__dfrtp_1
X_2664_ _0986_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2595_ net107 outputs.sig_gen.count\[6\] _0947_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__mux2_1
X_1546_ outputs.sig_gen.count\[14\] VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__inv_2
X_1615_ _1126_ outputs.shaper.count\[6\] outputs.divider_buffer\[8\] _1211_ VGND VGND
+ VPWR VPWR _1229_ sky130_fd_sc_hd__a2bb2o_1
X_1477_ outputs.sig_gen.count\[7\] VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__inv_2
X_2029_ net109 _0475_ _1003_ outputs.div.q\[24\] _0484_ VGND VGND VPWR VPWR _0071_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold260 outputs.div.divisor\[2\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331_ _1017_ VGND VGND VPWR VPWR inputs.keypad\[11\] sky130_fd_sc_hd__clkbuf_1
X_1400_ inputs.random_update_clock.count\[16\] inputs.random_update_clock.count\[17\]
+ _1060_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__and3_1
X_2380_ _0751_ _0786_ _0624_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3001_ clknet_leaf_36_clk _0207_ net24 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput6 gpio[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2647_ _0975_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2716_ clknet_leaf_37_clk net67 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2578_ net207 net109 _0936_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux2_1
X_1529_ _1100_ _1154_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1880_ _0362_ _0364_ _0360_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__o21ai_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2501_ inputs.octave_fsm.state\[2\] _0823_ _0228_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__or3b_1
X_2363_ _0572_ _0717_ _0562_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o21ai_1
X_1314_ _1005_ net12 VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__and2b_1
X_2294_ _0561_ _0564_ _0704_ _0663_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2432_ _0685_ _0833_ _0834_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1932_ _0406_ _0409_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a21oi_1
X_2981_ clknet_leaf_12_clk _0187_ net39 VGND VGND VPWR VPWR outputs.shaper.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1863_ outputs.div.m\[11\] outputs.div.m\[10\] _0321_ _0336_ VGND VGND VPWR VPWR
+ _0357_ sky130_fd_sc_hd__or4_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1794_ _0277_ _0293_ _0294_ _0252_ net173 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a32o_1
X_2415_ _0555_ _0549_ _0572_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2346_ outputs.div.divisor\[5\] _0754_ _0645_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2277_ _0685_ _0647_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2062_ _0503_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2200_ _0613_ _0598_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nand2_1
X_2131_ _0537_ _0542_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o21a_1
X_2964_ clknet_leaf_10_clk _0170_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ _1002_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
X_1846_ _0318_ _0326_ _0340_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o31ai_4
X_1777_ _0260_ _0266_ _0278_ _0264_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o211a_1
X_2895_ clknet_leaf_0_clk _0101_ VGND VGND VPWR VPWR outputs.divider_buffer2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ _0556_ _0537_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2680_ clknet_leaf_9_clk net142 net43 VGND VGND VPWR VPWR outputs.sample_rate.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1631_ _1188_ net21 outputs.scaled_buffer\[4\] VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21oi_1
X_1700_ _1089_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_4
X_1493_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_1562_ _1181_ VGND VGND VPWR VPWR inputs.wavetype_fsm.next_state\[0\] sky130_fd_sc_hd__clkbuf_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ _0494_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2114_ _0530_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2947_ clknet_leaf_8_clk _0153_ VGND VGND VPWR VPWR outputs.signal_buffer2\[4\] sky130_fd_sc_hd__dfxtp_1
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout28 net36 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
X_2878_ clknet_leaf_3_clk outputs.sig_gen.next_count\[7\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[7\] sky130_fd_sc_hd__dfrtp_2
X_1829_ _0318_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2801_ clknet_leaf_14_clk _0035_ net46 VGND VGND VPWR VPWR outputs.div.a\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2594_ _0948_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
X_1614_ _1126_ outputs.shaper.count\[6\] VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2732_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[9\] net30 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_2663_ _0985_ _0543_ _0983_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1545_ _1169_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_1476_ _1111_ outputs.sig_gen.count\[14\] outputs.divider_buffer\[16\] _1112_ _1113_
+ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2028_ outputs.div.q\[23\] _1083_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold261 outputs.div.divisor\[6\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold250 inputs.up.ff_out VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1330_ net1 net4 VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__and2b_1
Xinput7 gpio[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3000_ clknet_leaf_37_clk _0206_ net23 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_2646_ outputs.shaper.count\[13\] net232 _0966_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
X_2577_ _0939_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2715_ clknet_leaf_37_clk net89 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1459_ outputs.divider_buffer\[12\] outputs.sig_gen.count\[12\] VGND VGND VPWR VPWR
+ _1097_ sky130_fd_sc_hd__xor2_1
X_1528_ _1100_ _1154_ _1156_ _1131_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[9\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2500_ _0897_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2431_ _0561_ _0799_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1313_ _1008_ VGND VGND VPWR VPWR inputs.keypad\[2\] sky130_fd_sc_hd__clkbuf_1
X_2293_ _0656_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__inv_2
X_2362_ _0576_ _0765_ _0767_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2629_ _1089_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2980_ clknet_leaf_12_clk _0186_ net39 VGND VGND VPWR VPWR outputs.shaper.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1931_ _0406_ _0409_ _0398_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__o21a_1
X_1862_ outputs.div.a\[11\] VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__inv_2
X_1793_ _0288_ _0286_ _0292_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a21o_1
Xinput10 gpio[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2414_ _0567_ _0817_ _0818_ _0691_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR
+ _0819_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2276_ _0683_ _0684_ _0687_ _0578_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__o211a_1
X_2345_ _0642_ _0749_ _0750_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2061_ outputs.scaled_buffer\[6\] net138 _0497_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2130_ _0543_ _0535_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_1
X_2963_ clknet_leaf_10_clk _0169_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1914_ _0400_ _0402_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1845_ _0324_ _0331_ _0332_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o21ai_1
X_1776_ outputs.div.a\[2\] _0271_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nand2_1
X_2894_ clknet_leaf_0_clk _0100_ VGND VGND VPWR VPWR outputs.divider_buffer2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2328_ _0737_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ _0230_ _0671_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ _1231_ _1237_ _1238_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_53_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1492_ _1105_ _1110_ _1114_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__or4_4
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _1179_ _1180_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__and2_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2044_ _0998_ _0492_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__and3_1
X_2113_ net195 net220 _0522_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2946_ clknet_leaf_10_clk _0152_ VGND VGND VPWR VPWR outputs.signal_buffer2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2877_ clknet_leaf_2_clk outputs.sig_gen.next_count\[6\] net37 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout29 net31 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
X_1828_ _0324_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2_2
XFILLER_0_40_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1759_ outputs.div.m\[2\] _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__xnor2_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2800_ clknet_leaf_22_clk _0034_ net47 VGND VGND VPWR VPWR outputs.div.a\[13\] sky130_fd_sc_hd__dfrtp_1
X_2731_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[8\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_2593_ net150 outputs.sig_gen.count\[5\] _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__mux2_1
X_1544_ _1130_ _1167_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__and3_1
X_1613_ _1119_ outputs.shaper.count\[5\] VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2662_ _0556_ _1182_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__xor2_1
X_1475_ outputs.divider_buffer\[2\] outputs.sig_gen.count\[2\] VGND VGND VPWR VPWR
+ _1113_ sky130_fd_sc_hd__xor2_1
X_2027_ net103 _0475_ _1003_ outputs.div.q\[23\] _0483_ VGND VGND VPWR VPWR _0070_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ clknet_leaf_0_clk _0135_ net26 VGND VGND VPWR VPWR outputs.divider_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold240 outputs.div.a\[19\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 outputs.div.divisor\[13\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 outputs.div.divisor\[0\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput8 gpio[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2714_ clknet_leaf_37_clk net75 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2576_ net238 net103 _0936_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__mux2_1
X_2645_ _0974_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
X_1527_ outputs.sig_gen.count\[9\] _1153_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1458_ outputs.divider_buffer\[17\] VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__inv_2
X_1389_ inputs.random_update_clock.count\[13\] _1052_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2361_ _0768_ _0559_ _0564_ _0654_ _0578_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a41o_1
X_2430_ _0551_ _0652_ _0817_ _0685_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1312_ _1005_ net11 VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__and2b_1
X_2292_ _0700_ _0702_ _0230_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2628_ _0965_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
X_2559_ net205 net221 _0925_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ _0400_ _0410_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1861_ net179 _1004_ outputs.div.next_div _0355_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a22o_1
X_1792_ _0288_ _0286_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 gpio[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_12_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2413_ _0568_ _0549_ _0572_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__or3_1
X_2344_ _0247_ _0752_ _0642_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2275_ _0569_ _0559_ _0566_ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _0502_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2962_ clknet_leaf_10_clk _0168_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1913_ _0400_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2893_ clknet_leaf_0_clk _0099_ VGND VGND VPWR VPWR outputs.divider_buffer2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1775_ _1084_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ _0333_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2327_ net311 _0736_ _0645_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__mux2_1
X_2258_ _0669_ _0670_ _0626_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2189_ inputs.key_encoder.sync_keys\[13\] _1287_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__and2_2
XFILLER_0_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1560_ inputs.wavetype_fsm.state\[0\] inputs.mode_edge.det_edge VGND VGND VPWR VPWR
+ _1180_ sky130_fd_sc_hd__or2_1
X_1491_ _1118_ _1121_ _1125_ _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__or4_1
X_2112_ net270 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2043_ outputs.div.start _0489_ outputs.div.count\[3\] VGND VGND VPWR VPWR _0493_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2945_ clknet_leaf_10_clk _0151_ VGND VGND VPWR VPWR outputs.signal_buffer2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2876_ clknet_leaf_2_clk outputs.sig_gen.next_count\[5\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1827_ _0319_ _0323_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1758_ outputs.div.m\[0\] outputs.div.m\[1\] outputs.div.a\[25\] VGND VGND VPWR VPWR
+ _0262_ sky130_fd_sc_hd__o21ba_1
X_1689_ _0212_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2730_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[7\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_2661_ _0984_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2592_ _0512_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__buf_4
X_1474_ outputs.sig_gen.count\[16\] VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__inv_2
X_1543_ outputs.sig_gen.count\[13\] _1164_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__nand2_1
X_1612_ _1222_ _1223_ _1224_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2026_ outputs.div.q\[22\] _1083_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ clknet_leaf_20_clk net139 net47 VGND VGND VPWR VPWR outputs.div.q_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2928_ clknet_leaf_1_clk _0134_ net26 VGND VGND VPWR VPWR outputs.divider_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold263 outputs.div.divisor\[3\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _1062_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 inputs.random_update_clock.count\[18\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 inputs.down.ff_out VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 gpio[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_0_52_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2644_ outputs.shaper.count\[12\] net223 _0966_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__mux2_1
X_2713_ clknet_leaf_37_clk net68 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2575_ _0938_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_1457_ outputs.divider_buffer\[9\] VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__inv_2
X_1526_ _1155_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1388_ inputs.random_update_clock.count\[13\] _1052_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__or2_1
X_2009_ outputs.div.q\[14\] _0248_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1311_ _1007_ VGND VGND VPWR VPWR inputs.keypad\[1\] sky130_fd_sc_hd__clkbuf_1
X_2360_ _0686_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__clkbuf_4
X_2291_ _0670_ _0701_ _0626_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2627_ outputs.shaper.count\[4\] net249 _0916_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2558_ _0929_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_1509_ net290 _1138_ _1131_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o21ai_1
X_2489_ _0872_ _0887_ _0577_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_35_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1860_ _0351_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1791_ _0289_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 gpio[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2274_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__clkbuf_4
X_2343_ _0699_ _0751_ _0624_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__mux2_1
X_2412_ _0722_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_1989_ net210 _0413_ _0249_ net250 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2961_ clknet_leaf_10_clk _0167_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1912_ _0380_ _0383_ _0392_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o31a_2
X_1843_ outputs.div.a\[9\] _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2892_ clknet_leaf_1_clk _0098_ VGND VGND VPWR VPWR outputs.divider_buffer2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
X_1774_ net299 _1004_ _0275_ _0276_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2326_ _0674_ _0721_ _0728_ _0734_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__o32a_1
X_2257_ _0610_ _0621_ _0611_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2188_ _0585_ _0594_ _0598_ _0599_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1490_ _1126_ outputs.sig_gen.count\[7\] _1103_ outputs.sig_gen.count\[10\] _1127_
+ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2042_ _0491_ _1001_ _0490_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2111_ outputs.divider_buffer2\[14\] net269 _0522_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
Xhold1 inputs.keypad_synchronizer.half_sync\[7\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2944_ clknet_leaf_12_clk _0150_ VGND VGND VPWR VPWR outputs.signal_buffer2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2875_ clknet_leaf_2_clk outputs.sig_gen.next_count\[4\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[4\] sky130_fd_sc_hd__dfrtp_2
X_1826_ _0319_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1757_ outputs.div.a\[1\] VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__inv_2
X_1688_ outputs.div.m\[3\] net292 _1294_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _0555_ _0717_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1611_ _1119_ outputs.shaper.count\[5\] outputs.shaper.count\[4\] _1108_ VGND VGND
+ VPWR VPWR _1225_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2660_ _0982_ _0556_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__mux2_1
X_2591_ _0946_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
X_1542_ outputs.sig_gen.count\[13\] _1164_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__or2_1
X_1473_ outputs.divider_buffer\[14\] VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2025_ net101 _0475_ _1003_ outputs.div.q\[22\] _0482_ VGND VGND VPWR VPWR _0069_
+ sky130_fd_sc_hd__a221o_1
X_2927_ clknet_leaf_1_clk _0133_ net38 VGND VGND VPWR VPWR outputs.divider_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2858_ clknet_leaf_20_clk net144 net48 VGND VGND VPWR VPWR outputs.div.q_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold231 outputs.divider_buffer2\[14\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 outputs.div.divisor\[8\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 outputs.divider_buffer2\[10\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 outputs.div.divisor\[0\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ clknet_leaf_26_clk _0023_ net35 VGND VGND VPWR VPWR outputs.div.a\[2\] sky130_fd_sc_hd__dfrtp_1
X_1809_ _0277_ _0307_ _0308_ _0252_ net169 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a32o_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold264 inputs.random_note_generator.out\[12\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2574_ net254 net101 _0936_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__mux2_1
X_2643_ _0973_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
X_2712_ clknet_leaf_37_clk net71 net23 VGND VGND VPWR VPWR inputs.random_note_generator.out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1456_ _1092_ outputs.sig_gen.count\[1\] outputs.divider_buffer\[13\] _1093_ VGND
+ VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a2bb2o_1
X_1525_ _1130_ _1152_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1387_ _1054_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2008_ net107 _1090_ _0468_ outputs.div.q\[14\] _0473_ VGND VGND VPWR VPWR _0061_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _1005_ net10 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__and2b_1
X_2290_ _0602_ _0629_ _0238_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2557_ net206 net107 _0925_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__mux2_1
X_2626_ _0964_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1439_ net100 VGND VGND VPWR VPWR outputs.sample_rate.next_count\[0\] sky130_fd_sc_hd__inv_2
X_1508_ outputs.sig_gen.count\[4\] _1138_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__and2_1
X_2488_ _0656_ _0800_ _0575_ _0557_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 gpio[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ outputs.div.m\[5\] _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2411_ _0768_ _0813_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2273_ inputs.frequency_lut.rng\[4\] VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__clkbuf_4
X_2342_ _0618_ _0731_ _0238_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1988_ outputs.div.q\[2\] _0413_ _0249_ net213 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2609_ net302 outputs.sig_gen.count\[13\] _0947_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2960_ clknet_leaf_9_clk _0166_ VGND VGND VPWR VPWR outputs.signal_buffer2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1911_ _0378_ _0390_ _0391_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1842_ outputs.div.m\[10\] _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__xnor2_2
X_1773_ _0269_ _0274_ _1084_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2891_ clknet_leaf_1_clk _0097_ VGND VGND VPWR VPWR outputs.divider_buffer2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2325_ _0247_ _0625_ _0674_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o21ai_1
X_2256_ _0615_ _0668_ _0237_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux2_1
X_2187_ _0587_ _0591_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or3_4
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2041_ outputs.div.count\[3\] VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__inv_2
X_2110_ _0528_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
Xhold2 inputs.keypad_synchronizer.half_sync\[5\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2943_ clknet_leaf_15_clk _0149_ VGND VGND VPWR VPWR outputs.signal_buffer2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2874_ clknet_leaf_2_clk outputs.sig_gen.next_count\[3\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1825_ outputs.div.m\[8\] _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__xor2_1
X_1756_ _0250_ _0257_ _0256_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1687_ _0211_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
X_2308_ _0554_ _0564_ _0690_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2239_ _0535_ _0541_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2590_ net98 outputs.sig_gen.count\[4\] _0936_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__mux2_1
X_1610_ _1108_ outputs.shaper.count\[4\] VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1541_ _1166_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
X_1472_ _1106_ outputs.sig_gen.count\[3\] _1107_ outputs.sig_gen.count\[15\] _1109_
+ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2024_ outputs.div.q\[21\] _1083_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2857_ clknet_leaf_19_clk net123 net53 VGND VGND VPWR VPWR outputs.div.q_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2926_ clknet_leaf_1_clk _0132_ net38 VGND VGND VPWR VPWR outputs.divider_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _0073_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 outputs.div.oscillator_out\[10\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _0918_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 outputs.div.divisor\[16\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 outputs.div.divisor\[12\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
XFILLER_0_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2788_ clknet_leaf_24_clk _0022_ net33 VGND VGND VPWR VPWR outputs.div.a\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1808_ _0301_ _0306_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1739_ inputs.octave_fsm.state\[2\] _0228_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__and2_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2711_ clknet_leaf_37_clk net81 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2573_ net233 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2642_ net259 net228 _0966_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__mux2_1
X_1524_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1455_ outputs.sig_gen.count\[13\] VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__inv_2
X_1386_ _1052_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2007_ outputs.div.q\[13\] _0248_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2909_ clknet_leaf_34_clk _0115_ VGND VGND VPWR VPWR outputs.div.divisor\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2556_ _0928_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_2625_ outputs.shaper.count\[3\] net262 _0916_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__mux2_1
X_1507_ _1141_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2487_ inputs.frequency_lut.rng\[5\] _0686_ _0569_ _0717_ VGND VGND VPWR VPWR _0886_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1438_ _1084_ VGND VGND VPWR VPWR outputs.div.next_div sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1369_ inputs.random_update_clock.count\[6\] inputs.random_update_clock.count\[7\]
+ _1029_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 gpio[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_2341_ _0231_ _0671_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nand2_1
X_2410_ _0569_ _0652_ _0800_ _0814_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR
+ _0815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2272_ _0559_ _0658_ _0576_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1987_ net213 _0413_ _0249_ net261 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a22o_1
X_2608_ _0955_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_2539_ _0919_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1910_ _0398_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nand2_1
X_2890_ clknet_leaf_1_clk _0096_ VGND VGND VPWR VPWR outputs.divider_buffer2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1841_ _0321_ _0336_ _0320_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o21a_1
X_1772_ _0269_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2324_ _0230_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
X_2255_ _0601_ _0606_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and3_1
X_2186_ _0585_ _0592_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _0999_ _1084_ _0490_ _0405_ net162 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a32o_1
Xhold3 inputs.keypad_synchronizer.half_sync\[0\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2942_ clknet_leaf_12_clk _0148_ net39 VGND VGND VPWR VPWR outputs.divider_buffer\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2873_ clknet_leaf_11_clk outputs.sig_gen.next_count\[2\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1755_ net181 _1004_ outputs.div.next_div _0259_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a22o_1
X_1824_ _0320_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__nand2_1
X_1686_ outputs.div.m\[2\] net315 _1294_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2238_ _0535_ _0543_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or2b_1
X_2307_ _0543_ _0535_ _0556_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__and3b_2
X_2169_ inputs.key_encoder.sync_keys\[6\] _0582_ inputs.key_encoder.sync_keys\[7\]
+ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1540_ _1130_ _1163_ _1165_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1471_ _1108_ outputs.sig_gen.count\[5\] _1096_ outputs.sig_gen.count\[17\] VGND
+ VGND VPWR VPWR _1109_ sky130_fd_sc_hd__o22ai_1
X_2023_ outputs.div.oscillator_out\[13\] _0475_ _1003_ net152 _0481_ VGND VGND VPWR
+ VPWR _0068_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2856_ clknet_leaf_19_clk net164 net53 VGND VGND VPWR VPWR outputs.div.q_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2925_ clknet_leaf_1_clk _0131_ net38 VGND VGND VPWR VPWR outputs.divider_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1807_ _0301_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold222 outputs.div.oscillator_out\[8\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 outputs.divider_buffer2\[16\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _1280_ _1281_ _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__o21a_1
Xhold233 outputs.div.a\[9\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 outputs.div.a\[3\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ clknet_leaf_23_clk _0021_ net33 VGND VGND VPWR VPWR outputs.div.a\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold200 outputs.divider_buffer2\[0\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 outputs.div.divisor\[1\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1738_ _0235_ _0231_ _0236_ _0245_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2710_ clknet_leaf_37_clk net70 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2572_ net232 outputs.div.oscillator_out\[13\] _0936_ VGND VGND VPWR VPWR _0937_
+ sky130_fd_sc_hd__mux2_1
X_2641_ _0972_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
X_1454_ outputs.divider_buffer\[1\] VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1523_ outputs.sig_gen.count\[8\] _1150_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and2_1
X_1385_ inputs.random_update_clock.count\[11\] inputs.random_update_clock.count\[10\]
+ _1047_ inputs.random_update_clock.count\[12\] VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2006_ net150 _1090_ _0468_ outputs.div.q\[13\] _0472_ VGND VGND VPWR VPWR _0060_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2839_ clknet_leaf_15_clk net265 net50 VGND VGND VPWR VPWR outputs.div.q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2908_ clknet_leaf_34_clk _0114_ VGND VGND VPWR VPWR outputs.div.divisor\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
X_2624_ net189 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1437_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__clkbuf_4
X_2555_ net215 net150 _0925_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__mux2_1
X_1506_ _1130_ _1139_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__and3_1
X_2486_ _0885_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1299_ outputs.sample_rate.count\[7\] _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__nand2_1
X_1368_ _1040_ _1041_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 gpio[6] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2271_ _0555_ _0545_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__nor2_1
X_2340_ _0727_ _0740_ _0742_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1986_ net261 _0413_ outputs.div.next_div _0465_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ net127 outputs.sig_gen.count\[12\] _0947_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ outputs.divider_buffer\[15\] net195 _0916_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
X_2469_ _0686_ _0767_ _0862_ _0859_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ outputs.div.m\[9\] outputs.div.m\[8\] VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1771_ _0272_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2323_ _0679_ _0732_ _0624_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__mux2_1
X_2254_ _0598_ _0599_ _0616_ _0632_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2185_ _0595_ _0585_ _0593_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1969_ _0445_ _0448_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 inputs.keypad_synchronizer.half_sync\[11\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2941_ clknet_leaf_14_clk _0147_ net46 VGND VGND VPWR VPWR outputs.divider_buffer\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_2872_ clknet_leaf_12_clk outputs.sig_gen.next_count\[1\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[1\] sky130_fd_sc_hd__dfrtp_4
X_1823_ outputs.div.m\[7\] outputs.div.m\[6\] _0281_ _0296_ VGND VGND VPWR VPWR _0321_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_29_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1754_ _0250_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__xor2_1
X_1685_ _0210_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2306_ _0685_ _0550_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__nor2_1
X_2237_ _0536_ _0558_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2099_ net245 outputs.div.divisor\[8\] _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2168_ inputs.key_encoder.sync_keys\[4\] _0581_ inputs.key_encoder.sync_keys\[5\]
+ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1470_ outputs.divider_buffer\[5\] VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2022_ outputs.div.q\[20\] _1083_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold201 outputs.div.a\[18\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
X_2855_ clknet_leaf_19_clk net202 net53 VGND VGND VPWR VPWR outputs.div.q_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2924_ clknet_leaf_12_clk _0130_ VGND VGND VPWR VPWR outputs.div.divisor\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1806_ _0273_ _0279_ _0303_ _0292_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o41a_1
X_2786_ clknet_leaf_28_clk outputs.output_gen.pwm_unff net35 VGND VGND VPWR VPWR outputs.output_gen.pwm_ff
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold245 outputs.div.oscillator_out\[1\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
X_1599_ outputs.shaper.count\[3\] VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__inv_2
Xhold234 outputs.div.q_out\[4\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _0531_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ outputs.scaled_buffer\[7\] _1250_ _1254_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a21oi_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 outputs.div.divisor\[11\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold256 outputs.div.divisor\[4\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1737_ _0242_ _0244_ _0233_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2640_ net282 net243 _0966_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1453_ _1090_ _1091_ VGND VGND VPWR VPWR outputs.sample_rate.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_2571_ _0512_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__buf_4
X_1522_ outputs.sig_gen.count\[8\] _1150_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2005_ outputs.div.q\[12\] _0248_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1384_ inputs.random_update_clock.count\[11\] inputs.random_update_clock.count\[10\]
+ inputs.random_update_clock.count\[12\] _1047_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2907_ clknet_leaf_1_clk _0113_ VGND VGND VPWR VPWR outputs.div.divisor\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2838_ clknet_leaf_9_clk net160 net44 VGND VGND VPWR VPWR outputs.div.q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2769_ clknet_leaf_25_clk inputs.keypad\[0\] net34 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2554_ _0927_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
X_2623_ outputs.shaper.count\[2\] net188 _0916_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1436_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__buf_2
X_1505_ _1099_ _1136_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nand2_1
X_2485_ net269 _0884_ _0855_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__mux2_1
X_1367_ net216 _1029_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1298_ outputs.sample_rate.count\[6\] _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 gpio[7] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_0_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2270_ _0680_ _0681_ _0230_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1985_ _0457_ _0461_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2606_ _0954_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_2537_ net287 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1419_ outputs.output_gen.count\[2\] outputs.output_gen.count\[1\] outputs.output_gen.count\[0\]
+ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and3_1
X_2399_ _0784_ _0804_ _0611_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
X_2468_ _0823_ _0825_ _0230_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ outputs.div.a\[2\] _0271_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2184_ _0591_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or2_2
X_2253_ _0649_ _0655_ _0661_ _0665_ _0576_ _0578_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux4_1
X_2322_ _0698_ _0731_ _0611_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ _0277_ _0449_ _0450_ _0405_ net170 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1899_ outputs.div.a\[14\] _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 inputs.keypad_synchronizer.half_sync\[12\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2940_ clknet_leaf_12_clk _0146_ net46 VGND VGND VPWR VPWR outputs.divider_buffer\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2871_ clknet_leaf_1_clk outputs.sig_gen.next_count\[0\] net38 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[0\] sky130_fd_sc_hd__dfstp_2
X_1822_ _0253_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__buf_2
X_1753_ _0256_ _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1684_ outputs.div.m\[1\] outputs.div.divisor\[1\] _1294_ VGND VGND VPWR VPWR _0210_
+ sky130_fd_sc_hd__mux2_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0715_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_2167_ inputs.key_encoder.sync_keys\[1\] _0580_ inputs.key_encoder.sync_keys\[3\]
+ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a21oi_1
X_2236_ _0547_ _0647_ _0648_ _0538_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2098_ _0512_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2021_ net127 _0475_ _1003_ outputs.div.q\[20\] _0480_ VGND VGND VPWR VPWR _0067_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2923_ clknet_leaf_13_clk _0129_ VGND VGND VPWR VPWR outputs.div.divisor\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2854_ clknet_leaf_19_clk net106 net52 VGND VGND VPWR VPWR outputs.div.q_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold235 outputs.sig_gen.count\[4\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 outputs.output_gen.count\[3\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 outputs.div.divisor\[2\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
X_1805_ _0289_ _0291_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21o_1
Xhold202 outputs.divider_buffer2\[5\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2785_ clknet_leaf_28_clk inputs.keypad\[16\] net34 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1736_ _0228_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold246 outputs.sig_gen.count\[17\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ outputs.divider_buffer\[8\] _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__or2_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ outputs.scaled_buffer\[6\] net21 _1252_ _1247_ VGND VGND VPWR VPWR _1281_
+ sky130_fd_sc_hd__a31o_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold257 outputs.div.divisor\[12\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _0628_ _0630_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2570_ _0935_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1452_ net204 _0997_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1521_ _1150_ _1151_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[7\] sky130_fd_sc_hd__nor2_1
X_1383_ net191 _1049_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[11\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2004_ net98 _1090_ _0468_ outputs.div.q\[12\] _0471_ VGND VGND VPWR VPWR _0059_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2906_ clknet_leaf_12_clk _0112_ VGND VGND VPWR VPWR outputs.divider_buffer2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2837_ clknet_leaf_9_clk net110 net43 VGND VGND VPWR VPWR outputs.div.q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2699_ clknet_leaf_13_clk _0013_ net45 VGND VGND VPWR VPWR outputs.div.m\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2768_ clknet_leaf_28_clk net74 net36 VGND VGND VPWR VPWR inputs.key_encoder.octave_key_up
+ sky130_fd_sc_hd__dfrtp_1
X_1719_ inputs.octave_fsm.state\[1\] inputs.octave_fsm.state\[0\] VGND VGND VPWR VPWR
+ _0228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ net249 net98 _0925_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__mux2_1
X_2622_ _0962_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1504_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1435_ _1081_ _1001_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nor2_1
X_2484_ _0231_ _0534_ _0830_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__a31o_1
X_1366_ inputs.random_update_clock.count\[6\] _1029_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1297_ outputs.sample_rate.count\[4\] outputs.sample_rate.count\[5\] _0995_ VGND
+ VGND VPWR VPWR _0996_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 gpio[8] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1984_ outputs.div.m\[17\] outputs.div.a\[25\] _0407_ _0454_ _0459_ VGND VGND VPWR
+ VPWR _0464_ sky130_fd_sc_hd__o311a_1
XFILLER_0_55_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2605_ net304 outputs.sig_gen.count\[11\] _0947_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__mux2_1
X_2536_ outputs.divider_buffer\[14\] net286 _0916_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
X_2467_ _0868_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1418_ outputs.output_gen.count\[1\] net90 VGND VGND VPWR VPWR outputs.output_gen.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
X_1349_ inputs.random_update_clock.count\[3\] _1024_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__and2_1
X_2398_ _0597_ _0609_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2321_ _0729_ _0730_ _0604_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2252_ _0565_ _0663_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a21oi_1
X_2183_ _0596_ _0592_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1967_ _0443_ _0446_ _0448_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1898_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2519_ outputs.divider_buffer\[6\] net224 _0905_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 inputs.keypad_synchronizer.half_sync\[4\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2870_ clknet_leaf_22_clk net149 net49 VGND VGND VPWR VPWR outputs.output_gen.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
X_1821_ outputs.div.a\[7\] VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1752_ _0254_ _0255_ outputs.div.a\[0\] VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a21oi_1
X_1683_ _0209_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ net318 _0714_ _0645_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ _0521_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_2166_ inputs.key_encoder.sync_keys\[2\] VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__inv_2
X_2235_ _0551_ _0544_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2999_ clknet_leaf_37_clk _0205_ net23 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ net118 _1083_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2853_ clknet_leaf_22_clk net130 net47 VGND VGND VPWR VPWR outputs.div.q_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2922_ clknet_leaf_13_clk _0128_ VGND VGND VPWR VPWR outputs.div.divisor\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold247 outputs.div.oscillator_out\[13\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ net21 _1252_ outputs.scaled_buffer\[6\] VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__a21oi_1
Xhold258 outputs.div.divisor\[15\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 outputs.div.divisor\[14\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 outputs.divider_buffer2\[2\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _0516_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
X_1804_ _0287_ _0283_ _0291_ _0289_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o22a_1
Xhold203 _0519_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
X_2784_ clknet_leaf_38_clk inputs.keypad\[15\] net25 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1735_ inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[1\]
+ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1597_ outputs.shaper.count\[7\] VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2149_ _0535_ _0540_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or2_1
X_2218_ _0594_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1520_ outputs.sig_gen.count\[7\] _1147_ _1131_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1451_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1382_ _1051_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2003_ outputs.div.q\[11\] _0248_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2836_ clknet_leaf_8_clk net104 net43 VGND VGND VPWR VPWR outputs.div.q\[23\] sky130_fd_sc_hd__dfrtp_1
X_2905_ clknet_leaf_13_clk _0111_ VGND VGND VPWR VPWR outputs.divider_buffer2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1718_ _0227_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
X_1649_ _1260_ _1261_ _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__o21a_1
X_2698_ clknet_leaf_23_clk _0012_ net45 VGND VGND VPWR VPWR outputs.div.m\[12\] sky130_fd_sc_hd__dfrtp_2
X_2767_ clknet_leaf_33_clk net80 net34 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2552_ _0926_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_2621_ outputs.shaper.count\[1\] net234 _0916_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__mux2_1
X_1503_ _1099_ _1136_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2483_ _0727_ _0881_ _0882_ _0859_ _0603_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__o221a_1
X_1296_ outputs.sample_rate.count\[3\] _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__and2_1
X_1434_ outputs.sample_rate.count\[6\] outputs.sample_rate.count\[7\] _0996_ VGND
+ VGND VPWR VPWR _1081_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1365_ _1028_ _1029_ _1039_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2819_ clknet_leaf_19_clk _0053_ net52 VGND VGND VPWR VPWR outputs.div.q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 gpio[9] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1983_ _1084_ _0462_ _0463_ _0405_ net274 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a32o_1
X_2604_ _0953_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2535_ _0917_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2466_ net312 _0867_ _0855_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux2_1
X_1417_ net90 VGND VGND VPWR VPWR outputs.output_gen.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2397_ _0231_ _0733_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nand2_1
X_1348_ _1024_ _1025_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2251_ _0564_ _0567_ _0555_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__a21oi_1
X_2320_ _0585_ _0597_ _0616_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2182_ _0595_ _1291_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1966_ _0443_ _0446_ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1897_ outputs.div.m\[15\] _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2518_ _0908_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_2449_ _0230_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 outputs.output_gen.pwm_ff VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ _0301_ _0306_ _0314_ _0317_ _0313_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o32a_2
XFILLER_0_80_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1751_ outputs.div.a\[0\] _0254_ _0255_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__and3_1
X_1682_ outputs.div.m\[0\] net297 _1294_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2303_ _0642_ _0703_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o21ai_1
X_2234_ _0554_ _0558_ _0540_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2096_ net231 outputs.div.divisor\[7\] _0513_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__mux2_1
X_2165_ _0553_ _0560_ _0571_ _0574_ _0576_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1949_ _0430_ _0433_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2998_ clknet_leaf_36_clk _0204_ net24 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2852_ clknet_leaf_22_clk _0086_ net47 VGND VGND VPWR VPWR outputs.scaled_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2921_ clknet_leaf_13_clk _0127_ VGND VGND VPWR VPWR outputs.div.divisor\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1803_ _0288_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__nand2_1
X_2783_ clknet_leaf_28_clk inputs.keypad\[14\] net36 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold226 outputs.div.a\[20\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 outputs.shaper.count\[11\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ _1189_ _1195_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__or3_1
Xhold248 outputs.scaled_buffer\[7\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _0529_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ outputs.output_gen.count\[5\] _1256_ _1278_ outputs.output_gen.count\[6\]
+ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a22o_1
Xhold259 outputs.output_gen.count\[4\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 outputs.div.divisor\[3\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1734_ inputs.octave_fsm.state\[1\] inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\]
+ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2217_ _0585_ _0598_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__or2_1
X_2079_ net43 _1081_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__and2_1
X_2148_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1450_ _1081_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1381_ _1043_ _1049_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__and3_1
X_2002_ net92 _1090_ _0468_ outputs.div.q\[11\] _0470_ VGND VGND VPWR VPWR _0058_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2835_ clknet_leaf_8_clk net102 net41 VGND VGND VPWR VPWR outputs.div.q\[22\] sky130_fd_sc_hd__dfrtp_1
X_2904_ clknet_leaf_13_clk _0110_ VGND VGND VPWR VPWR outputs.divider_buffer2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2766_ clknet_leaf_28_clk net77 net31 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1579_ _1192_ outputs.shaper.count\[15\] _1190_ outputs.divider_buffer\[15\] VGND
+ VGND VPWR VPWR _1193_ sky130_fd_sc_hd__a2bb2o_1
X_1717_ outputs.div.m\[17\] outputs.div.divisor\[17\] _0218_ VGND VGND VPWR VPWR _0227_
+ sky130_fd_sc_hd__mux2_1
X_1648_ outputs.scaled_buffer\[2\] _1250_ _1254_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__a21oi_1
X_2697_ clknet_leaf_13_clk _0011_ net45 VGND VGND VPWR VPWR outputs.div.m\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2620_ _0961_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2551_ net262 net92 _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
X_1502_ _1137_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1433_ net148 _1078_ VGND VGND VPWR VPWR outputs.output_gen.next_count\[7\] sky130_fd_sc_hd__xnor2_1
X_2482_ _0686_ _0569_ _0537_ _0546_ _0577_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a41o_1
X_1295_ outputs.sample_rate.count\[2\] outputs.sample_rate.count\[1\] outputs.sample_rate.count\[0\]
+ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__and3_1
X_1364_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__buf_2
X_2818_ clknet_leaf_19_clk _0052_ net52 VGND VGND VPWR VPWR outputs.div.q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2749_ clknet_leaf_30_clk inputs.down.ff_in net27 VGND VGND VPWR VPWR inputs.down.det_edge
+ sky130_fd_sc_hd__dfrtp_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 nrst VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ _0454_ _0457_ _0461_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2603_ net309 outputs.sig_gen.count\[10\] _0947_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ outputs.divider_buffer\[13\] net272 _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2396_ _0793_ _0795_ _0798_ _0801_ _0686_ _0727_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux4_1
X_1347_ net174 inputs.random_update_clock.count\[0\] net194 VGND VGND VPWR VPWR _1025_
+ sky130_fd_sc_hd__a21oi_1
X_1416_ _1071_ VGND VGND VPWR VPWR inputs.down.in sky130_fd_sc_hd__clkbuf_1
X_2465_ _0642_ _0861_ _0864_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire21 _1244_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2250_ _0551_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2181_ _1288_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1965_ outputs.div.a\[22\] _0427_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1896_ _0320_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__nand2_1
X_2517_ outputs.divider_buffer\[5\] net257 _0905_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2379_ _0238_ _0784_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__o21ai_1
X_2448_ _0624_ _0824_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold8 inputs.keypad_synchronizer.half_sync\[9\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ outputs.div.m\[0\] outputs.div.m\[1\] _0253_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1681_ _1081_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _0646_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
X_2302_ _0674_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__or2_1
X_2164_ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__clkbuf_4
X_2095_ _0520_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1948_ _0430_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1879_ _0370_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2997_ clknet_leaf_36_clk _0203_ net24 VGND VGND VPWR VPWR inputs.frequency_lut.rng\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2920_ clknet_leaf_12_clk _0126_ VGND VGND VPWR VPWR outputs.div.divisor\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2851_ clknet_leaf_20_clk _0085_ net47 VGND VGND VPWR VPWR outputs.scaled_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ _0287_ _0283_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__nand2_1
X_1733_ _0236_ _0241_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__xnor2_1
X_2782_ clknet_leaf_38_clk inputs.keypad\[13\] net24 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold249 outputs.div.oscillator_out\[11\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 outputs.div.a\[17\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 outputs.signal_buffer2\[8\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ _1198_ _1200_ _1203_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__or4_1
Xhold227 outputs.shaper.count\[10\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ outputs.scaled_buffer\[6\] _1250_ _1277_ _1246_ _1254_ VGND VGND VPWR VPWR
+ _1278_ sky130_fd_sc_hd__a221oi_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold238 inputs.random_update_clock.count\[5\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ _0551_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2216_ _0597_ _0627_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2078_ net171 _0506_ _0510_ outputs.div.q\[7\] VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1380_ inputs.random_update_clock.count\[10\] _1047_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2001_ outputs.div.q\[10\] _0248_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and2_1
X_2903_ clknet_leaf_12_clk _0109_ VGND VGND VPWR VPWR outputs.divider_buffer2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2834_ clknet_leaf_7_clk net153 net41 VGND VGND VPWR VPWR outputs.div.q\[21\] sky130_fd_sc_hd__dfrtp_1
X_1716_ _0226_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2696_ clknet_leaf_23_clk _0010_ net45 VGND VGND VPWR VPWR outputs.div.m\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2765_ clknet_leaf_35_clk net78 net28 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1578_ outputs.divider_buffer\[16\] VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__inv_2
X_1647_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] net21 _1247_ VGND VGND
+ VPWR VPWR _1261_ sky130_fd_sc_hd__a31o_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2550_ _0512_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1501_ _1130_ _1135_ _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1432_ _1080_ VGND VGND VPWR VPWR outputs.output_gen.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_1363_ _1032_ _1035_ _1036_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2481_ _0765_ _0879_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2679_ clknet_leaf_16_clk outputs.sample_rate.next_count\[3\] net51 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_2817_ clknet_leaf_18_clk _0051_ net52 VGND VGND VPWR VPWR outputs.div.q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2748_ clknet_leaf_31_clk inputs.down.in net31 VGND VGND VPWR VPWR inputs.down.ff_out
+ sky130_fd_sc_hd__dfrtp_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ _0454_ _0457_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ _1089_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__clkbuf_4
X_2602_ _0952_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2464_ _0247_ _0806_ _0865_ _0533_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__o211a_1
X_1346_ inputs.random_update_clock.count\[1\] inputs.random_update_clock.count\[0\]
+ inputs.random_update_clock.count\[2\] VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and3_1
X_1415_ inputs.key_encoder.octave_key_up inputs.key_encoder.sync_keys\[15\] VGND VGND
+ VPWR VPWR _1071_ sky130_fd_sc_hd__and2b_1
X_2395_ _0552_ _0799_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ _0587_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1964_ net283 _0413_ _0446_ _0447_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1895_ outputs.div.m\[14\] outputs.div.m\[13\] outputs.div.m\[12\] _0357_ VGND VGND
+ VPWR VPWR _0386_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_13_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2516_ _0907_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
X_2447_ _0611_ _0626_ _0823_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__or3_1
X_1329_ _1016_ VGND VGND VPWR VPWR inputs.keypad\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2378_ _0611_ _0758_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold9 inputs.keypad_synchronizer.half_sync\[8\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1680_ _1293_ VGND VGND VPWR VPWR outputs.output_gen.pwm_unff sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2301_ _0705_ _0708_ _0710_ _0711_ _0685_ _0577_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
X_2232_ net317 _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2163_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2094_ net224 net208 _0513_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux2_1
X_2996_ clknet_leaf_9_clk _0202_ net44 VGND VGND VPWR VPWR outputs.shaper.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1947_ _0431_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1878_ _0367_ _0369_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2850_ clknet_leaf_20_clk _0084_ net48 VGND VGND VPWR VPWR outputs.scaled_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold206 outputs.div.q\[0\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1663_ outputs.scaled_buffer\[5\] _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__xnor2_1
Xhold217 outputs.divider_buffer2\[13\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1801_ _0299_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2781_ clknet_leaf_38_clk inputs.keypad\[12\] net25 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ inputs.octave_fsm.state\[1\] _0235_ _0238_ _0240_ VGND VGND VPWR VPWR _0241_
+ sky130_fd_sc_hd__o31a_1
Xhold228 outputs.div.a\[22\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 outputs.sig_gen.count\[2\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ _1204_ _1205_ _1206_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__or4_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2077_ net138 _0506_ _0510_ outputs.div.q\[6\] VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__o22a_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2146_ _0555_ _0557_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o21ai_1
X_2215_ _0596_ _0592_ _0627_ _0619_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a311o_1
XFILLER_0_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2979_ clknet_leaf_15_clk _0185_ net50 VGND VGND VPWR VPWR outputs.shaper.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2000_ outputs.div.oscillator_out\[2\] _1090_ _0468_ net120 _0469_ VGND VGND VPWR
+ VPWR _0057_ sky130_fd_sc_hd__a221o_1
X_2833_ clknet_leaf_7_clk net128 net41 VGND VGND VPWR VPWR outputs.div.q\[20\] sky130_fd_sc_hd__dfrtp_1
X_2902_ clknet_leaf_12_clk _0108_ VGND VGND VPWR VPWR outputs.divider_buffer2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ outputs.div.m\[16\] net298 _0218_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
X_1646_ outputs.scaled_buffer\[0\] net21 outputs.scaled_buffer\[1\] VGND VGND VPWR
+ VPWR _1260_ sky130_fd_sc_hd__a21oi_1
X_2695_ clknet_leaf_13_clk _0009_ net45 VGND VGND VPWR VPWR outputs.div.m\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2764_ clknet_leaf_38_clk net60 net25 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1577_ outputs.divider_buffer\[15\] _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__nor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2129_ inputs.frequency_lut.rng\[1\] VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__buf_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1500_ outputs.sig_gen.count\[0\] outputs.sig_gen.count\[1\] outputs.sig_gen.count\[2\]
+ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nand3_1
X_2480_ _0552_ _0537_ _0872_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__o21a_1
X_1431_ _1078_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__and2_1
X_1362_ inputs.random_update_clock.count\[20\] inputs.random_update_clock.count\[22\]
+ inputs.random_update_clock.count\[21\] VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2816_ clknet_leaf_19_clk _0050_ net52 VGND VGND VPWR VPWR outputs.div.q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2678_ clknet_leaf_16_clk outputs.sample_rate.next_count\[2\] net51 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1629_ _1219_ _1210_ _1239_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__or4b_1
X_2747_ clknet_leaf_25_clk inputs.mode_edge.ff_in net34 VGND VGND VPWR VPWR inputs.mode_edge.det_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1980_ _0459_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
X_2601_ outputs.div.oscillator_out\[9\] outputs.sig_gen.count\[9\] _0947_ VGND VGND
+ VPWR VPWR _0952_ sky130_fd_sc_hd__mux2_1
X_2532_ _0915_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2463_ _0229_ _0823_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__or2_1
X_1414_ net94 net88 inputs.key_encoder.sync_keys\[14\] VGND VGND VPWR VPWR inputs.key_encoder.mode_key
+ sky130_fd_sc_hd__nor3b_1
X_1345_ net174 net157 VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
X_2394_ _0554_ _0544_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1963_ _0445_ _0439_ _0442_ _1001_ _1294_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a311oi_1
X_1894_ _0277_ _0384_ _0385_ _0252_ net126 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2515_ outputs.divider_buffer\[4\] net239 _0905_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__mux2_1
X_2446_ _0843_ _0845_ _0847_ _0848_ _0576_ _0578_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__mux4_1
X_1328_ net1 net3 VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2377_ _1288_ _0592_ _0627_ _0636_ _0628_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__a311o_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _0512_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2300_ _0573_ _0648_ _0653_ _0561_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2093_ net258 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_2162_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__clkbuf_4
X_2995_ clknet_leaf_9_clk _0201_ net43 VGND VGND VPWR VPWR outputs.shaper.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1946_ outputs.div.a\[19\] _0414_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or2_1
X_1877_ _0367_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2429_ _0540_ _0541_ _0800_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _0295_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold218 outputs.shaper.count\[14\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold207 outputs.signal_buffer2\[3\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ outputs.scaled_buffer\[4\] _1188_ net21 VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2780_ clknet_leaf_38_clk inputs.keypad\[11\] net25 VGND VGND VPWR VPWR inputs.keypad_synchronizer.half_sync\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1731_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] _0239_ _0231_ _0233_
+ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o32a_1
Xhold229 inputs.random_update_clock.count\[17\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ outputs.divider_buffer\[13\] _1199_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nor2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _0604_ _0605_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__nor2_1
X_2076_ net143 _0506_ _0510_ outputs.div.q\[5\] VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__o22a_1
X_2145_ _0537_ _0558_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nand2_2
X_2978_ clknet_leaf_9_clk _0184_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_1929_ _0415_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold90 outputs.sample_rate.count\[3\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
X_2832_ clknet_leaf_6_clk net119 net41 VGND VGND VPWR VPWR outputs.div.q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2901_ clknet_leaf_2_clk _0107_ VGND VGND VPWR VPWR outputs.divider_buffer2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2763_ clknet_leaf_38_clk net59 net25 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1576_ outputs.shaper.count\[14\] VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1714_ _0225_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
X_1645_ outputs.scaled_buffer\[3\] _1250_ _1258_ _1246_ _1254_ VGND VGND VPWR VPWR
+ _1259_ sky130_fd_sc_hd__a221oi_2
X_2694_ clknet_leaf_23_clk _0008_ net45 VGND VGND VPWR VPWR outputs.div.m\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2059_ outputs.scaled_buffer\[5\] net143 _0497_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2128_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__nand2_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ outputs.output_gen.count\[6\] _1076_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1361_ inputs.random_update_clock.count\[16\] inputs.random_update_clock.count\[19\]
+ inputs.random_update_clock.count\[18\] inputs.random_update_clock.count\[17\] VGND
+ VGND VPWR VPWR _1036_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2815_ clknet_leaf_19_clk net214 net52 VGND VGND VPWR VPWR outputs.div.q\[2\] sky130_fd_sc_hd__dfrtp_1
X_2746_ clknet_leaf_25_clk net95 net34 VGND VGND VPWR VPWR inputs.mode_edge.ff_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2677_ clknet_leaf_17_clk outputs.sample_rate.next_count\[1\] net51 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1628_ _1224_ _1227_ _1240_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__and4_1
X_1559_ inputs.wavetype_fsm.state\[0\] inputs.mode_edge.det_edge VGND VGND VPWR VPWR
+ _1179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2600_ _0951_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2531_ outputs.divider_buffer\[12\] net226 _0905_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1413_ net96 _1069_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[22\]
+ sky130_fd_sc_hd__xnor2_1
X_2462_ _0768_ _0796_ _0862_ _0863_ _0578_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__a311o_1
X_2393_ _0540_ _0547_ _0764_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ net157 VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2729_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[6\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1962_ _0439_ _0442_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1893_ _0380_ _0383_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2514_ _0906_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_2376_ _0777_ _0779_ _0781_ _0782_ _0686_ _0578_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__mux4_1
X_2445_ _0562_ _0540_ _0537_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1327_ _1015_ VGND VGND VPWR VPWR inputs.keypad\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0534_ _0579_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2092_ net257 outputs.div.divisor\[5\] _0513_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__mux2_1
X_2161_ inputs.frequency_lut.rng\[4\] VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__inv_2
X_2994_ clknet_leaf_8_clk _0200_ net43 VGND VGND VPWR VPWR outputs.shaper.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1945_ outputs.div.a\[19\] _0414_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1876_ outputs.div.m\[13\] _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _0657_ _0764_ inputs.frequency_lut.rng\[3\] VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__o21a_1
X_2359_ _0542_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold208 outputs.div.count\[1\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 outputs.div.a\[25\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
X_1592_ outputs.divider_buffer\[12\] _1201_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nor2_1
X_1661_ outputs.output_gen.count\[5\] _1256_ _1269_ _1273_ _1274_ VGND VGND VPWR VPWR
+ _1275_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ inputs.octave_fsm.state\[1\] _0233_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nor2_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0556_ _0543_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nor2_1
X_2213_ _0600_ _0591_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or2b_1
X_2075_ outputs.div.q_out\[4\] _0506_ _0510_ net122 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2977_ clknet_leaf_8_clk _0183_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1928_ outputs.div.a\[17\] _0414_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or2_1
X_1859_ _0353_ _0344_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold91 outputs.div.q\[18\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 _0064_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
X_2900_ clknet_leaf_3_clk _0106_ VGND VGND VPWR VPWR outputs.divider_buffer2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2831_ clknet_leaf_6_clk net147 net41 VGND VGND VPWR VPWR outputs.div.q\[18\] sky130_fd_sc_hd__dfrtp_1
X_1713_ outputs.div.m\[15\] net313 _0218_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2762_ clknet_leaf_33_clk net86 net32 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1575_ _1111_ outputs.shaper.count\[13\] VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__and2_1
X_1644_ outputs.scaled_buffer\[2\] _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__xnor2_1
X_2693_ clknet_leaf_34_clk _0007_ net33 VGND VGND VPWR VPWR outputs.div.m\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _0538_ inputs.frequency_lut.rng\[1\] VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2058_ _0501_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1360_ _1033_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2676_ clknet_leaf_16_clk outputs.sample_rate.next_count\[0\] net51 VGND VGND VPWR
+ VPWR outputs.sample_rate.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_2814_ clknet_leaf_18_clk _0048_ net52 VGND VGND VPWR VPWR outputs.div.q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2745_ clknet_leaf_29_clk net97 net31 VGND VGND VPWR VPWR inputs.random_update_clock.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1558_ net186 _1177_ _1178_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[17\]
+ sky130_fd_sc_hd__a21oi_1
X_1627_ _1220_ _1223_ _1228_ _1212_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__and4b_1
X_1489_ _1107_ outputs.sig_gen.count\[15\] _1119_ outputs.sig_gen.count\[6\] VGND
+ VGND VPWR VPWR _1127_ sky130_fd_sc_hd__a2bb2o_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2530_ _0914_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1343_ _1023_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_2392_ _0552_ _0547_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a21o_1
X_1412_ _1070_ VGND VGND VPWR VPWR inputs.random_update_clock.next_count\[21\] sky130_fd_sc_hd__clkbuf_1
X_2461_ _0552_ _0657_ _0656_ _0766_ _0576_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__o311a_1
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2728_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[5\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_2659_ _1039_ _0642_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nand2_4
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ _0443_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__nand2_1
X_1892_ _0380_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2513_ outputs.divider_buffer\[3\] net251 _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_1326_ _1005_ net18 VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__and2b_1
X_2444_ _0818_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2375_ _0552_ _0542_ _0662_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2160_ _0562_ _0547_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ net240 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_2993_ clknet_leaf_7_clk _0199_ net42 VGND VGND VPWR VPWR outputs.shaper.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1944_ _0402_ _0426_ _0428_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o211a_1
X_1875_ outputs.div.m\[12\] _0357_ _0320_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ _0761_ _0830_ _0247_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1309_ _1006_ VGND VGND VPWR VPWR inputs.keypad\[0\] sky130_fd_sc_hd__clkbuf_1
X_2289_ _0669_ _0699_ _0623_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux2_1
X_2358_ _0568_ _0537_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold209 outputs.div.q\[25\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
X_1591_ outputs.divider_buffer\[11\] _1202_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__nor2_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ outputs.output_gen.count\[4\] _1272_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__or2_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ inputs.octave_fsm.state\[0\] inputs.octave_fsm.state\[2\] inputs.octave_fsm.state\[1\]
+ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__a21oi_4
X_2143_ _0556_ _0543_ _0536_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2074_ net163 _0506_ _0510_ outputs.div.q\[3\] VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__o22a_1
X_2976_ clknet_leaf_7_clk _0182_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_1927_ outputs.div.a\[17\] _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__nand2_1
X_1858_ _0352_ _0338_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1789_ outputs.div.m\[4\] _0281_ _0253_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold92 _0065_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 _0063_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 outputs.div.q\[9\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ clknet_leaf_6_clk net135 net41 VGND VGND VPWR VPWR outputs.div.q\[17\] sky130_fd_sc_hd__dfrtp_1
X_1712_ _0224_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1643_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] net21 VGND VGND VPWR
+ VPWR _1257_ sky130_fd_sc_hd__o21ai_1
X_2692_ clknet_leaf_34_clk _0006_ net33 VGND VGND VPWR VPWR outputs.div.m\[6\] sky130_fd_sc_hd__dfrtp_1
X_2761_ clknet_leaf_0_clk net63 net25 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ outputs.scaled_buffer\[0\] outputs.scaled_buffer\[1\] outputs.scaled_buffer\[3\]
+ outputs.scaled_buffer\[2\] VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__or4_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ outputs.scaled_buffer\[4\] net289 _0497_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2126_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__clkbuf_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2959_ clknet_leaf_8_clk _0165_ VGND VGND VPWR VPWR outputs.signal_buffer2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2813_ clknet_leaf_18_clk _0047_ net52 VGND VGND VPWR VPWR outputs.div.q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1626_ _1096_ outputs.shaper.count\[16\] outputs.shaper.count\[0\] _1092_ VGND VGND
+ VPWR VPWR _1240_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2675_ _0993_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2744_ clknet_leaf_28_clk inputs.random_update_clock.next_count\[21\] net31 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[21\] sky130_fd_sc_hd__dfrtp_1
X_1557_ net186 _1177_ _1131_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__o21ai_1
X_1488_ outputs.divider_buffer\[7\] VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__inv_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2109_ net272 outputs.div.divisor\[13\] _0522_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2460_ _0555_ _0657_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nand2_1
X_1342_ net1 outputs.pwm_output VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__and2b_1
X_2391_ _0660_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__nand2_1
X_1411_ _1043_ _1068_ _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2589_ _0945_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_1609_ outputs.divider_buffer\[4\] _1213_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__or2_1
X_2658_ _0980_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__xnor2_1
X_2727_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[4\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ outputs.div.a\[21\] _0414_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1891_ _0362_ _0364_ _0372_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o31a_1
X_2512_ _1089_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__buf_4
X_2443_ _0549_ _0662_ _0562_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1325_ _1014_ VGND VGND VPWR VPWR inputs.keypad\[8\] sky130_fd_sc_hd__clkbuf_1
X_2374_ _0707_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ net239 outputs.div.divisor\[4\] _0513_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2992_ clknet_leaf_7_clk _0198_ net42 VGND VGND VPWR VPWR outputs.shaper.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1943_ _0406_ _0409_ _0417_ _0419_ _0423_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ outputs.div.a\[12\] VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2426_ _0805_ _0829_ _0624_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1308_ _1005_ net2 VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__and2b_1
X_2288_ _0678_ _0698_ _0237_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_1
X_2357_ _0568_ _0722_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1590_ outputs.divider_buffer\[10\] _1196_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor2_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2073_ net201 _0506_ _0510_ outputs.div.q\[2\] VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__o22a_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _0612_ _0622_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux2_1
X_2142_ inputs.frequency_lut.rng\[0\] VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__clkbuf_4
X_2975_ clknet_leaf_7_clk _0181_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1926_ outputs.div.m\[17\] _0407_ _0320_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o21a_2
X_1857_ outputs.div.a\[9\] VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__inv_2
X_1788_ outputs.div.a\[4\] VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2409_ _0650_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold82 _0056_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 outputs.div.a\[14\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 outputs.output_gen.count\[7\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 inputs.mode_edge.ff_out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1642_ _1245_ _1248_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o21a_1
X_1711_ outputs.div.m\[14\] net269 _0218_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
X_2691_ clknet_leaf_34_clk _0005_ net32 VGND VGND VPWR VPWR outputs.div.m\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2760_ clknet_leaf_32_clk net64 net28 VGND VGND VPWR VPWR inputs.key_encoder.sync_keys\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1573_ _1187_ VGND VGND VPWR VPWR inputs.up.ff_in sky130_fd_sc_hd__clkbuf_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ _0500_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_2125_ _0538_ inputs.frequency_lut.rng\[1\] VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2958_ clknet_leaf_8_clk _0164_ VGND VGND VPWR VPWR outputs.signal_buffer2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ _0395_ _0397_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2889_ clknet_leaf_1_clk _0095_ VGND VGND VPWR VPWR outputs.divider_buffer2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2812_ clknet_leaf_15_clk _0046_ net50 VGND VGND VPWR VPWR outputs.div.a\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2743_ clknet_leaf_31_clk inputs.random_update_clock.next_count\[20\] net31 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1556_ _1112_ _1174_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__nor2_1
X_1625_ _1229_ _1225_ _1215_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__or4b_1
XFILLER_0_26_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2674_ _0992_ _0727_ _0983_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1487_ _1122_ outputs.sig_gen.count\[0\] _1123_ outputs.sig_gen.count\[11\] _1124_
+ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__a221o_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2039_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2108_ _0527_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ inputs.random_update_clock.count\[21\] _1066_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1341_ _1022_ VGND VGND VPWR VPWR inputs.keypad\[16\] sky130_fd_sc_hd__buf_1
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2390_ _0551_ _0536_ _0540_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand3_1
X_2726_ clknet_leaf_32_clk inputs.random_update_clock.next_count\[3\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2588_ net92 outputs.sig_gen.count\[3\] _0936_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__mux2_1
X_1539_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__inv_2
X_1608_ _1215_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or2_1
X_2657_ _0562_ _1182_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold190 outputs.divider_buffer2\[8\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1890_ _0360_ _0381_ _0371_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a21o_1
X_2511_ _0904_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
X_2442_ _0569_ _0550_ _0844_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2373_ _0563_ _0704_ _0568_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1324_ _1005_ net17 VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2709_ clknet_leaf_37_clk net83 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1942_ outputs.div.a\[18\] outputs.div.a\[17\] _0427_ VGND VGND VPWR VPWR _0428_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ clknet_leaf_5_clk _0197_ net42 VGND VGND VPWR VPWR outputs.shaper.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1873_ _0277_ _0365_ _0366_ _0252_ net165 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2356_ inputs.frequency_lut.rng\[0\] inputs.frequency_lut.rng\[2\] VGND VGND VPWR
+ VPWR _0764_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2425_ _0238_ _0823_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1307_ net1 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_4
X_2287_ _0635_ _0620_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2210_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2072_ net105 _0506_ _0510_ outputs.div.q\[1\] VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__o22a_1
X_2141_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_4
X_2974_ clknet_leaf_7_clk _0180_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_1925_ _1003_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1856_ _0348_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nand2_1
X_1787_ _0287_ _0283_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2408_ _0810_ _0812_ _0577_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21o_1
X_2339_ _0686_ _0744_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold61 outputs.div.q\[15\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 outputs.div.oscillator_out\[12\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 outputs.div.q_out\[1\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 outputs.div.q_out\[6\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 outputs.output_gen.next_count\[7\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1710_ _0223_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_1641_ outputs.scaled_buffer\[5\] _1250_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2690_ clknet_leaf_34_clk _0004_ net32 VGND VGND VPWR VPWR outputs.div.m\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1572_ net305 inputs.key_encoder.octave_key_up VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__and2b_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ inputs.frequency_lut.rng\[0\] VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__inv_2
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2055_ outputs.scaled_buffer\[3\] net163 _0497_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2957_ clknet_leaf_7_clk _0163_ VGND VGND VPWR VPWR outputs.signal_buffer2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2888_ clknet_leaf_11_clk outputs.sig_gen.next_count\[17\] net44 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[17\] sky130_fd_sc_hd__dfrtp_1
X_1908_ _0395_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
X_1839_ net288 _1004_ _0334_ _0335_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
X_2811_ clknet_leaf_15_clk _0045_ net50 VGND VGND VPWR VPWR outputs.div.a\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2742_ clknet_leaf_31_clk inputs.random_update_clock.next_count\[19\] net31 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1555_ _1112_ _1174_ _1176_ _1131_ VGND VGND VPWR VPWR outputs.sig_gen.next_count\[16\]
+ sky130_fd_sc_hd__o211a_1
X_1624_ _1096_ outputs.shaper.count\[16\] outputs.shaper.count\[17\] VGND VGND VPWR
+ VPWR _1238_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2673_ _0768_ _1182_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
X_1486_ _1122_ outputs.sig_gen.count\[0\] _1108_ outputs.sig_gen.count\[5\] VGND VGND
+ VPWR VPWR _1124_ sky130_fd_sc_hd__a2bb2o_1
X_2107_ net226 net276 _0522_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ outputs.div.count\[2\] outputs.div.count\[1\] outputs.div.count\[0\] VGND
+ VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1340_ net1 net8 VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
X_2725_ clknet_leaf_32_clk inputs.random_update_clock.next_count\[2\] net29 VGND VGND
+ VPWR VPWR inputs.random_update_clock.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_2656_ _0727_ _0768_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2587_ _0944_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_1538_ outputs.sig_gen.count\[12\] _1162_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1607_ _1216_ _1219_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a21oi_1
X_1469_ outputs.divider_buffer\[15\] VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold180 _0923_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold191 outputs.divider_buffer2\[11\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ outputs.divider_buffer\[2\] net291 _0497_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1323_ _1013_ VGND VGND VPWR VPWR inputs.keypad\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2372_ _0552_ _0764_ _0778_ _0652_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__a22oi_1
X_2441_ _0554_ _0650_ _0656_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2639_ _0971_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2708_ clknet_leaf_37_clk net73 net22 VGND VGND VPWR VPWR inputs.random_note_generator.out\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1941_ _0414_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__buf_2
X_2990_ clknet_leaf_6_clk _0196_ net42 VGND VGND VPWR VPWR outputs.shaper.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1872_ _0362_ _0364_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1306_ _1004_ VGND VGND VPWR VPWR outputs.div.next_start sky130_fd_sc_hd__inv_2
X_2424_ _0828_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
X_2355_ _0231_ _0761_ _0762_ _0534_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__o211a_1
X_2286_ inputs.key_encoder.sync_keys\[12\] _1288_ _0596_ _0593_ _0586_ VGND VGND VPWR
+ VPWR _0697_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2140_ inputs.frequency_lut.rng\[3\] VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__inv_2
X_2071_ net129 _0506_ _0510_ outputs.div.q\[0\] VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__o22a_1
X_2973_ clknet_leaf_5_clk _0179_ VGND VGND VPWR VPWR outputs.div.oscillator_out\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_1924_ net260 _1004_ outputs.div.next_div _0412_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__a22o_1
X_1855_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1786_ outputs.div.a\[3\] VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2407_ _0547_ _0811_ _0569_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__o21ai_1
X_2338_ _0685_ _0564_ _0746_ inputs.frequency_lut.rng\[5\] VGND VGND VPWR VPWR _0747_
+ sky130_fd_sc_hd__a31o_1
X_2269_ _0612_ _0634_ _0626_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold40 inputs.key_encoder.mode_key VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _0067_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 outputs.div.oscillator_out\[5\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0062_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0088_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _0093_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1640_ net21 _1251_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_21_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ _1186_ VGND VGND VPWR VPWR inputs.down.ff_in sky130_fd_sc_hd__clkbuf_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__clkbuf_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ _0499_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2956_ clknet_leaf_7_clk _0162_ VGND VGND VPWR VPWR outputs.signal_buffer2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2887_ clknet_leaf_8_clk outputs.sig_gen.next_count\[16\] net44 VGND VGND VPWR VPWR
+ outputs.sig_gen.count\[16\] sky130_fd_sc_hd__dfrtp_1
X_1907_ outputs.div.m\[16\] _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__xnor2_1
X_1838_ _0324_ _0327_ _0333_ _1084_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1769_ outputs.div.a\[2\] _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2810_ clknet_leaf_16_clk _0044_ net54 VGND VGND VPWR VPWR outputs.div.a\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2672_ _0983_ _0981_ _0991_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__o21ai_1
X_2741_ clknet_leaf_30_clk inputs.random_update_clock.next_count\[18\] net29 VGND
+ VGND VPWR VPWR inputs.random_update_clock.count\[18\] sky130_fd_sc_hd__dfrtp_1
X_1554_ _1112_ _1174_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__nand2_1
X_1623_ _1189_ _1195_ _1235_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__o31ai_1
X_1485_ outputs.divider_buffer\[11\] VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__inv_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

