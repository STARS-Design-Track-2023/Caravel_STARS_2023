// This is the unpowered netlist.
module silly_synthesizer (clk,
    cs,
    nrst,
    pwm,
    gpio);
 input clk;
 input cs;
 input nrst;
 output pwm;
 input [16:0] gpio;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \inputs.down.det_edge ;
 wire \inputs.down.ff_in ;
 wire \inputs.down.ff_out ;
 wire \inputs.down.in ;
 wire \inputs.frequency_lut.rng[0] ;
 wire \inputs.frequency_lut.rng[1] ;
 wire \inputs.frequency_lut.rng[2] ;
 wire \inputs.frequency_lut.rng[3] ;
 wire \inputs.frequency_lut.rng[4] ;
 wire \inputs.frequency_lut.rng[5] ;
 wire \inputs.key_encoder.mode_key ;
 wire \inputs.key_encoder.octave_key_up ;
 wire \inputs.key_encoder.sync_keys[0] ;
 wire \inputs.key_encoder.sync_keys[10] ;
 wire \inputs.key_encoder.sync_keys[11] ;
 wire \inputs.key_encoder.sync_keys[12] ;
 wire \inputs.key_encoder.sync_keys[13] ;
 wire \inputs.key_encoder.sync_keys[14] ;
 wire \inputs.key_encoder.sync_keys[15] ;
 wire \inputs.key_encoder.sync_keys[1] ;
 wire \inputs.key_encoder.sync_keys[2] ;
 wire \inputs.key_encoder.sync_keys[3] ;
 wire \inputs.key_encoder.sync_keys[4] ;
 wire \inputs.key_encoder.sync_keys[5] ;
 wire \inputs.key_encoder.sync_keys[6] ;
 wire \inputs.key_encoder.sync_keys[7] ;
 wire \inputs.key_encoder.sync_keys[8] ;
 wire \inputs.key_encoder.sync_keys[9] ;
 wire \inputs.keypad[0] ;
 wire \inputs.keypad[10] ;
 wire \inputs.keypad[11] ;
 wire \inputs.keypad[12] ;
 wire \inputs.keypad[13] ;
 wire \inputs.keypad[14] ;
 wire \inputs.keypad[15] ;
 wire \inputs.keypad[16] ;
 wire \inputs.keypad[1] ;
 wire \inputs.keypad[2] ;
 wire \inputs.keypad[3] ;
 wire \inputs.keypad[4] ;
 wire \inputs.keypad[5] ;
 wire \inputs.keypad[6] ;
 wire \inputs.keypad[7] ;
 wire \inputs.keypad[8] ;
 wire \inputs.keypad[9] ;
 wire \inputs.keypad_synchronizer.half_sync[0] ;
 wire \inputs.keypad_synchronizer.half_sync[10] ;
 wire \inputs.keypad_synchronizer.half_sync[11] ;
 wire \inputs.keypad_synchronizer.half_sync[12] ;
 wire \inputs.keypad_synchronizer.half_sync[13] ;
 wire \inputs.keypad_synchronizer.half_sync[14] ;
 wire \inputs.keypad_synchronizer.half_sync[15] ;
 wire \inputs.keypad_synchronizer.half_sync[16] ;
 wire \inputs.keypad_synchronizer.half_sync[1] ;
 wire \inputs.keypad_synchronizer.half_sync[2] ;
 wire \inputs.keypad_synchronizer.half_sync[3] ;
 wire \inputs.keypad_synchronizer.half_sync[4] ;
 wire \inputs.keypad_synchronizer.half_sync[5] ;
 wire \inputs.keypad_synchronizer.half_sync[6] ;
 wire \inputs.keypad_synchronizer.half_sync[7] ;
 wire \inputs.keypad_synchronizer.half_sync[8] ;
 wire \inputs.keypad_synchronizer.half_sync[9] ;
 wire \inputs.mode_edge.det_edge ;
 wire \inputs.mode_edge.ff_in ;
 wire \inputs.mode_edge.ff_out ;
 wire \inputs.octave_fsm.octave_key_up ;
 wire \inputs.octave_fsm.state[0] ;
 wire \inputs.octave_fsm.state[1] ;
 wire \inputs.octave_fsm.state[2] ;
 wire \inputs.random_note_generator.feedback ;
 wire \inputs.random_note_generator.out[0] ;
 wire \inputs.random_note_generator.out[10] ;
 wire \inputs.random_note_generator.out[11] ;
 wire \inputs.random_note_generator.out[12] ;
 wire \inputs.random_note_generator.out[13] ;
 wire \inputs.random_note_generator.out[14] ;
 wire \inputs.random_note_generator.out[15] ;
 wire \inputs.random_note_generator.out[1] ;
 wire \inputs.random_note_generator.out[2] ;
 wire \inputs.random_note_generator.out[3] ;
 wire \inputs.random_note_generator.out[4] ;
 wire \inputs.random_note_generator.out[5] ;
 wire \inputs.random_note_generator.out[6] ;
 wire \inputs.random_note_generator.out[7] ;
 wire \inputs.random_note_generator.out[8] ;
 wire \inputs.random_note_generator.out[9] ;
 wire \inputs.random_update_clock.count[0] ;
 wire \inputs.random_update_clock.count[10] ;
 wire \inputs.random_update_clock.count[11] ;
 wire \inputs.random_update_clock.count[12] ;
 wire \inputs.random_update_clock.count[13] ;
 wire \inputs.random_update_clock.count[14] ;
 wire \inputs.random_update_clock.count[15] ;
 wire \inputs.random_update_clock.count[16] ;
 wire \inputs.random_update_clock.count[17] ;
 wire \inputs.random_update_clock.count[18] ;
 wire \inputs.random_update_clock.count[19] ;
 wire \inputs.random_update_clock.count[1] ;
 wire \inputs.random_update_clock.count[20] ;
 wire \inputs.random_update_clock.count[21] ;
 wire \inputs.random_update_clock.count[22] ;
 wire \inputs.random_update_clock.count[2] ;
 wire \inputs.random_update_clock.count[3] ;
 wire \inputs.random_update_clock.count[4] ;
 wire \inputs.random_update_clock.count[5] ;
 wire \inputs.random_update_clock.count[6] ;
 wire \inputs.random_update_clock.count[7] ;
 wire \inputs.random_update_clock.count[8] ;
 wire \inputs.random_update_clock.count[9] ;
 wire \inputs.random_update_clock.next_count[0] ;
 wire \inputs.random_update_clock.next_count[10] ;
 wire \inputs.random_update_clock.next_count[11] ;
 wire \inputs.random_update_clock.next_count[12] ;
 wire \inputs.random_update_clock.next_count[13] ;
 wire \inputs.random_update_clock.next_count[14] ;
 wire \inputs.random_update_clock.next_count[15] ;
 wire \inputs.random_update_clock.next_count[16] ;
 wire \inputs.random_update_clock.next_count[17] ;
 wire \inputs.random_update_clock.next_count[18] ;
 wire \inputs.random_update_clock.next_count[19] ;
 wire \inputs.random_update_clock.next_count[1] ;
 wire \inputs.random_update_clock.next_count[20] ;
 wire \inputs.random_update_clock.next_count[21] ;
 wire \inputs.random_update_clock.next_count[22] ;
 wire \inputs.random_update_clock.next_count[2] ;
 wire \inputs.random_update_clock.next_count[3] ;
 wire \inputs.random_update_clock.next_count[4] ;
 wire \inputs.random_update_clock.next_count[5] ;
 wire \inputs.random_update_clock.next_count[6] ;
 wire \inputs.random_update_clock.next_count[7] ;
 wire \inputs.random_update_clock.next_count[8] ;
 wire \inputs.random_update_clock.next_count[9] ;
 wire \inputs.up.ff_in ;
 wire \inputs.up.ff_out ;
 wire \inputs.wavetype_fsm.next_state[0] ;
 wire \inputs.wavetype_fsm.next_state[1] ;
 wire \inputs.wavetype_fsm.state[0] ;
 wire \inputs.wavetype_fsm.state[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \outputs.div.a[0] ;
 wire \outputs.div.a[10] ;
 wire \outputs.div.a[11] ;
 wire \outputs.div.a[12] ;
 wire \outputs.div.a[13] ;
 wire \outputs.div.a[14] ;
 wire \outputs.div.a[15] ;
 wire \outputs.div.a[16] ;
 wire \outputs.div.a[17] ;
 wire \outputs.div.a[18] ;
 wire \outputs.div.a[19] ;
 wire \outputs.div.a[1] ;
 wire \outputs.div.a[20] ;
 wire \outputs.div.a[21] ;
 wire \outputs.div.a[22] ;
 wire \outputs.div.a[23] ;
 wire \outputs.div.a[24] ;
 wire \outputs.div.a[25] ;
 wire \outputs.div.a[2] ;
 wire \outputs.div.a[3] ;
 wire \outputs.div.a[4] ;
 wire \outputs.div.a[5] ;
 wire \outputs.div.a[6] ;
 wire \outputs.div.a[7] ;
 wire \outputs.div.a[8] ;
 wire \outputs.div.a[9] ;
 wire \outputs.div.count[0] ;
 wire \outputs.div.count[1] ;
 wire \outputs.div.count[2] ;
 wire \outputs.div.count[3] ;
 wire \outputs.div.count[4] ;
 wire \outputs.div.div ;
 wire \outputs.div.divisor[0] ;
 wire \outputs.div.divisor[10] ;
 wire \outputs.div.divisor[11] ;
 wire \outputs.div.divisor[12] ;
 wire \outputs.div.divisor[13] ;
 wire \outputs.div.divisor[14] ;
 wire \outputs.div.divisor[15] ;
 wire \outputs.div.divisor[16] ;
 wire \outputs.div.divisor[17] ;
 wire \outputs.div.divisor[1] ;
 wire \outputs.div.divisor[2] ;
 wire \outputs.div.divisor[3] ;
 wire \outputs.div.divisor[4] ;
 wire \outputs.div.divisor[5] ;
 wire \outputs.div.divisor[6] ;
 wire \outputs.div.divisor[7] ;
 wire \outputs.div.divisor[8] ;
 wire \outputs.div.divisor[9] ;
 wire \outputs.div.m[0] ;
 wire \outputs.div.m[10] ;
 wire \outputs.div.m[11] ;
 wire \outputs.div.m[12] ;
 wire \outputs.div.m[13] ;
 wire \outputs.div.m[14] ;
 wire \outputs.div.m[15] ;
 wire \outputs.div.m[16] ;
 wire \outputs.div.m[17] ;
 wire \outputs.div.m[1] ;
 wire \outputs.div.m[2] ;
 wire \outputs.div.m[3] ;
 wire \outputs.div.m[4] ;
 wire \outputs.div.m[5] ;
 wire \outputs.div.m[6] ;
 wire \outputs.div.m[7] ;
 wire \outputs.div.m[8] ;
 wire \outputs.div.m[9] ;
 wire \outputs.div.next_div ;
 wire \outputs.div.next_start ;
 wire \outputs.div.oscillator_out[0] ;
 wire \outputs.div.oscillator_out[10] ;
 wire \outputs.div.oscillator_out[11] ;
 wire \outputs.div.oscillator_out[12] ;
 wire \outputs.div.oscillator_out[13] ;
 wire \outputs.div.oscillator_out[14] ;
 wire \outputs.div.oscillator_out[15] ;
 wire \outputs.div.oscillator_out[16] ;
 wire \outputs.div.oscillator_out[17] ;
 wire \outputs.div.oscillator_out[1] ;
 wire \outputs.div.oscillator_out[2] ;
 wire \outputs.div.oscillator_out[3] ;
 wire \outputs.div.oscillator_out[4] ;
 wire \outputs.div.oscillator_out[5] ;
 wire \outputs.div.oscillator_out[6] ;
 wire \outputs.div.oscillator_out[7] ;
 wire \outputs.div.oscillator_out[8] ;
 wire \outputs.div.oscillator_out[9] ;
 wire \outputs.div.q[0] ;
 wire \outputs.div.q[10] ;
 wire \outputs.div.q[11] ;
 wire \outputs.div.q[12] ;
 wire \outputs.div.q[13] ;
 wire \outputs.div.q[14] ;
 wire \outputs.div.q[15] ;
 wire \outputs.div.q[16] ;
 wire \outputs.div.q[17] ;
 wire \outputs.div.q[18] ;
 wire \outputs.div.q[19] ;
 wire \outputs.div.q[1] ;
 wire \outputs.div.q[20] ;
 wire \outputs.div.q[21] ;
 wire \outputs.div.q[22] ;
 wire \outputs.div.q[23] ;
 wire \outputs.div.q[24] ;
 wire \outputs.div.q[25] ;
 wire \outputs.div.q[26] ;
 wire \outputs.div.q[2] ;
 wire \outputs.div.q[3] ;
 wire \outputs.div.q[4] ;
 wire \outputs.div.q[5] ;
 wire \outputs.div.q[6] ;
 wire \outputs.div.q[7] ;
 wire \outputs.div.q[8] ;
 wire \outputs.div.q[9] ;
 wire \outputs.div.q_out[0] ;
 wire \outputs.div.q_out[1] ;
 wire \outputs.div.q_out[2] ;
 wire \outputs.div.q_out[3] ;
 wire \outputs.div.q_out[4] ;
 wire \outputs.div.q_out[5] ;
 wire \outputs.div.q_out[6] ;
 wire \outputs.div.q_out[7] ;
 wire \outputs.div.start ;
 wire \outputs.divider_buffer[0] ;
 wire \outputs.divider_buffer[10] ;
 wire \outputs.divider_buffer[11] ;
 wire \outputs.divider_buffer[12] ;
 wire \outputs.divider_buffer[13] ;
 wire \outputs.divider_buffer[14] ;
 wire \outputs.divider_buffer[15] ;
 wire \outputs.divider_buffer[16] ;
 wire \outputs.divider_buffer[17] ;
 wire \outputs.divider_buffer[1] ;
 wire \outputs.divider_buffer[2] ;
 wire \outputs.divider_buffer[3] ;
 wire \outputs.divider_buffer[4] ;
 wire \outputs.divider_buffer[5] ;
 wire \outputs.divider_buffer[6] ;
 wire \outputs.divider_buffer[7] ;
 wire \outputs.divider_buffer[8] ;
 wire \outputs.divider_buffer[9] ;
 wire \outputs.output_gen.count[0] ;
 wire \outputs.output_gen.count[1] ;
 wire \outputs.output_gen.count[2] ;
 wire \outputs.output_gen.count[3] ;
 wire \outputs.output_gen.count[4] ;
 wire \outputs.output_gen.count[5] ;
 wire \outputs.output_gen.count[6] ;
 wire \outputs.output_gen.count[7] ;
 wire \outputs.output_gen.next_count[0] ;
 wire \outputs.output_gen.next_count[1] ;
 wire \outputs.output_gen.next_count[2] ;
 wire \outputs.output_gen.next_count[3] ;
 wire \outputs.output_gen.next_count[4] ;
 wire \outputs.output_gen.next_count[5] ;
 wire \outputs.output_gen.next_count[6] ;
 wire \outputs.output_gen.next_count[7] ;
 wire \outputs.output_gen.pwm_ff ;
 wire \outputs.output_gen.pwm_unff ;
 wire \outputs.pwm_output ;
 wire \outputs.sample_rate.count[0] ;
 wire \outputs.sample_rate.count[1] ;
 wire \outputs.sample_rate.count[2] ;
 wire \outputs.sample_rate.count[3] ;
 wire \outputs.sample_rate.count[4] ;
 wire \outputs.sample_rate.count[5] ;
 wire \outputs.sample_rate.count[6] ;
 wire \outputs.sample_rate.count[7] ;
 wire \outputs.sample_rate.next_count[0] ;
 wire \outputs.sample_rate.next_count[1] ;
 wire \outputs.sample_rate.next_count[2] ;
 wire \outputs.sample_rate.next_count[3] ;
 wire \outputs.sample_rate.next_count[4] ;
 wire \outputs.sample_rate.next_count[5] ;
 wire \outputs.sample_rate.next_count[6] ;
 wire \outputs.sample_rate.next_count[7] ;
 wire \outputs.scaled_buffer[0] ;
 wire \outputs.scaled_buffer[1] ;
 wire \outputs.scaled_buffer[2] ;
 wire \outputs.scaled_buffer[3] ;
 wire \outputs.scaled_buffer[4] ;
 wire \outputs.scaled_buffer[5] ;
 wire \outputs.scaled_buffer[6] ;
 wire \outputs.scaled_buffer[7] ;
 wire \outputs.shaper.count[0] ;
 wire \outputs.shaper.count[10] ;
 wire \outputs.shaper.count[11] ;
 wire \outputs.shaper.count[12] ;
 wire \outputs.shaper.count[13] ;
 wire \outputs.shaper.count[14] ;
 wire \outputs.shaper.count[15] ;
 wire \outputs.shaper.count[16] ;
 wire \outputs.shaper.count[17] ;
 wire \outputs.shaper.count[1] ;
 wire \outputs.shaper.count[2] ;
 wire \outputs.shaper.count[3] ;
 wire \outputs.shaper.count[4] ;
 wire \outputs.shaper.count[5] ;
 wire \outputs.shaper.count[6] ;
 wire \outputs.shaper.count[7] ;
 wire \outputs.shaper.count[8] ;
 wire \outputs.shaper.count[9] ;
 wire \outputs.sig_gen.count[0] ;
 wire \outputs.sig_gen.count[10] ;
 wire \outputs.sig_gen.count[11] ;
 wire \outputs.sig_gen.count[12] ;
 wire \outputs.sig_gen.count[13] ;
 wire \outputs.sig_gen.count[14] ;
 wire \outputs.sig_gen.count[15] ;
 wire \outputs.sig_gen.count[16] ;
 wire \outputs.sig_gen.count[17] ;
 wire \outputs.sig_gen.count[1] ;
 wire \outputs.sig_gen.count[2] ;
 wire \outputs.sig_gen.count[3] ;
 wire \outputs.sig_gen.count[4] ;
 wire \outputs.sig_gen.count[5] ;
 wire \outputs.sig_gen.count[6] ;
 wire \outputs.sig_gen.count[7] ;
 wire \outputs.sig_gen.count[8] ;
 wire \outputs.sig_gen.count[9] ;
 wire \outputs.sig_gen.next_count[0] ;
 wire \outputs.sig_gen.next_count[10] ;
 wire \outputs.sig_gen.next_count[11] ;
 wire \outputs.sig_gen.next_count[12] ;
 wire \outputs.sig_gen.next_count[13] ;
 wire \outputs.sig_gen.next_count[14] ;
 wire \outputs.sig_gen.next_count[15] ;
 wire \outputs.sig_gen.next_count[16] ;
 wire \outputs.sig_gen.next_count[17] ;
 wire \outputs.sig_gen.next_count[1] ;
 wire \outputs.sig_gen.next_count[2] ;
 wire \outputs.sig_gen.next_count[3] ;
 wire \outputs.sig_gen.next_count[4] ;
 wire \outputs.sig_gen.next_count[5] ;
 wire \outputs.sig_gen.next_count[6] ;
 wire \outputs.sig_gen.next_count[7] ;
 wire \outputs.sig_gen.next_count[8] ;
 wire \outputs.sig_gen.next_count[9] ;
 wire \outputs.signal_buffer2[0] ;
 wire \outputs.signal_buffer2[10] ;
 wire \outputs.signal_buffer2[11] ;
 wire \outputs.signal_buffer2[12] ;
 wire \outputs.signal_buffer2[13] ;
 wire \outputs.signal_buffer2[14] ;
 wire \outputs.signal_buffer2[15] ;
 wire \outputs.signal_buffer2[16] ;
 wire \outputs.signal_buffer2[17] ;
 wire \outputs.signal_buffer2[1] ;
 wire \outputs.signal_buffer2[2] ;
 wire \outputs.signal_buffer2[3] ;
 wire \outputs.signal_buffer2[4] ;
 wire \outputs.signal_buffer2[5] ;
 wire \outputs.signal_buffer2[6] ;
 wire \outputs.signal_buffer2[7] ;
 wire \outputs.signal_buffer2[8] ;
 wire \outputs.signal_buffer2[9] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_96 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__and3_1 _1239_ (.A(\outputs.sample_rate.count[1] ),
    .B(\outputs.sample_rate.count[0] ),
    .C(\outputs.sample_rate.count[2] ),
    .X(_0906_));
 sky130_fd_sc_hd__and2_1 _1240_ (.A(\outputs.sample_rate.count[3] ),
    .B(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__and3_1 _1241_ (.A(\outputs.sample_rate.count[4] ),
    .B(\outputs.sample_rate.count[5] ),
    .C(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__and2_1 _1242_ (.A(\outputs.sample_rate.count[6] ),
    .B(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_4 _1243_ (.A(\outputs.sample_rate.count[7] ),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__a21o_1 _1244_ (.A1(\outputs.div.count[1] ),
    .A2(\outputs.div.count[0] ),
    .B1(\outputs.div.count[2] ),
    .X(_0911_));
 sky130_fd_sc_hd__inv_2 _1245_ (.A(\outputs.div.start ),
    .Y(_0912_));
 sky130_fd_sc_hd__a31o_1 _1246_ (.A1(\outputs.div.count[3] ),
    .A2(\outputs.div.count[4] ),
    .A3(_0911_),
    .B1(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__and2_1 _1247_ (.A(_0910_),
    .B(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_4 _1248_ (.A(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_4 _1249_ (.A(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__inv_2 _1250_ (.A(_0916_),
    .Y(\outputs.div.next_start ));
 sky130_fd_sc_hd__clkbuf_8 _1251_ (.A(net1),
    .X(_0917_));
 sky130_fd_sc_hd__and2b_1 _1252_ (.A_N(_0917_),
    .B(net2),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _1253_ (.A(_0918_),
    .X(\inputs.keypad[0] ));
 sky130_fd_sc_hd__and2b_1 _1254_ (.A_N(_0917_),
    .B(net10),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _1255_ (.A(_0919_),
    .X(\inputs.keypad[1] ));
 sky130_fd_sc_hd__and2b_1 _1256_ (.A_N(_0917_),
    .B(net11),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _1257_ (.A(_0920_),
    .X(\inputs.keypad[2] ));
 sky130_fd_sc_hd__and2b_1 _1258_ (.A_N(_0917_),
    .B(net12),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _1259_ (.A(_0921_),
    .X(\inputs.keypad[3] ));
 sky130_fd_sc_hd__and2b_1 _1260_ (.A_N(_0917_),
    .B(net13),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _1261_ (.A(_0922_),
    .X(\inputs.keypad[4] ));
 sky130_fd_sc_hd__and2b_1 _1262_ (.A_N(_0917_),
    .B(net14),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(_0923_),
    .X(\inputs.keypad[5] ));
 sky130_fd_sc_hd__and2b_1 _1264_ (.A_N(_0917_),
    .B(net15),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _1265_ (.A(_0924_),
    .X(\inputs.keypad[6] ));
 sky130_fd_sc_hd__and2b_1 _1266_ (.A_N(_0917_),
    .B(net16),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _1267_ (.A(_0925_),
    .X(\inputs.keypad[7] ));
 sky130_fd_sc_hd__and2b_1 _1268_ (.A_N(_0917_),
    .B(net17),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _1269_ (.A(_0926_),
    .X(\inputs.keypad[8] ));
 sky130_fd_sc_hd__and2b_1 _1270_ (.A_N(_0917_),
    .B(net18),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _1271_ (.A(_0927_),
    .X(\inputs.keypad[9] ));
 sky130_fd_sc_hd__and2b_1 _1272_ (.A_N(net1),
    .B(net3),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _1273_ (.A(_0928_),
    .X(\inputs.keypad[10] ));
 sky130_fd_sc_hd__and2b_1 _1274_ (.A_N(net1),
    .B(net4),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_1 _1275_ (.A(_0929_),
    .X(\inputs.keypad[11] ));
 sky130_fd_sc_hd__and2b_1 _1276_ (.A_N(net1),
    .B(net5),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _1277_ (.A(_0930_),
    .X(\inputs.keypad[12] ));
 sky130_fd_sc_hd__and2b_1 _1278_ (.A_N(net1),
    .B(net9),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _1279_ (.A(_0931_),
    .X(\inputs.keypad[13] ));
 sky130_fd_sc_hd__and2b_1 _1280_ (.A_N(net1),
    .B(net6),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _1281_ (.A(_0932_),
    .X(\inputs.keypad[14] ));
 sky130_fd_sc_hd__and2b_1 _1282_ (.A_N(net1),
    .B(net7),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_1 _1283_ (.A(_0933_),
    .X(\inputs.keypad[15] ));
 sky130_fd_sc_hd__and2b_1 _1284_ (.A_N(net1),
    .B(net8),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _1285_ (.A(_0934_),
    .X(\inputs.keypad[16] ));
 sky130_fd_sc_hd__and2b_1 _1286_ (.A_N(net1),
    .B(\outputs.pwm_output ),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _1287_ (.A(_0935_),
    .X(net20));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(net169),
    .Y(\inputs.random_update_clock.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1289_ (.A(net214),
    .B(net169),
    .X(\inputs.random_update_clock.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1290_ (.A(\inputs.random_update_clock.count[1] ),
    .B(\inputs.random_update_clock.count[0] ),
    .C(\inputs.random_update_clock.count[2] ),
    .X(_0936_));
 sky130_fd_sc_hd__a21oi_1 _1291_ (.A1(\inputs.random_update_clock.count[1] ),
    .A2(\inputs.random_update_clock.count[0] ),
    .B1(net202),
    .Y(_0937_));
 sky130_fd_sc_hd__nor2_1 _1292_ (.A(_0936_),
    .B(net203),
    .Y(\inputs.random_update_clock.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1293_ (.A(\inputs.random_update_clock.count[3] ),
    .B(_0936_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _1294_ (.A(net212),
    .B(_0936_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_1 _1295_ (.A(_0938_),
    .B(_0939_),
    .Y(\inputs.random_update_clock.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1296_ (.A(net200),
    .B(_0938_),
    .X(\inputs.random_update_clock.next_count[4] ));
 sky130_fd_sc_hd__a21oi_1 _1297_ (.A1(\inputs.random_update_clock.count[4] ),
    .A2(_0938_),
    .B1(net296),
    .Y(_0940_));
 sky130_fd_sc_hd__and3_1 _1298_ (.A(\inputs.random_update_clock.count[4] ),
    .B(\inputs.random_update_clock.count[5] ),
    .C(_0938_),
    .X(_0941_));
 sky130_fd_sc_hd__or4bb_1 _1299_ (.A(\inputs.random_update_clock.count[4] ),
    .B(\inputs.random_update_clock.count[6] ),
    .C_N(\inputs.random_update_clock.count[7] ),
    .D_N(\inputs.random_update_clock.count[5] ),
    .X(_0942_));
 sky130_fd_sc_hd__or4_1 _1300_ (.A(\inputs.random_update_clock.count[1] ),
    .B(\inputs.random_update_clock.count[0] ),
    .C(\inputs.random_update_clock.count[3] ),
    .D(\inputs.random_update_clock.count[2] ),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_1 _1301_ (.A(_0942_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__or4b_1 _1302_ (.A(\inputs.random_update_clock.count[12] ),
    .B(\inputs.random_update_clock.count[15] ),
    .C(\inputs.random_update_clock.count[14] ),
    .D_N(\inputs.random_update_clock.count[13] ),
    .X(_0945_));
 sky130_fd_sc_hd__or4bb_1 _1303_ (.A(\inputs.random_update_clock.count[9] ),
    .B(\inputs.random_update_clock.count[11] ),
    .C_N(\inputs.random_update_clock.count[10] ),
    .D_N(\inputs.random_update_clock.count[8] ),
    .X(_0946_));
 sky130_fd_sc_hd__nor2_1 _1304_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__and4bb_1 _1305_ (.A_N(\inputs.random_update_clock.count[16] ),
    .B_N(\inputs.random_update_clock.count[19] ),
    .C(\inputs.random_update_clock.count[18] ),
    .D(\inputs.random_update_clock.count[17] ),
    .X(_0948_));
 sky130_fd_sc_hd__nor3b_1 _1306_ (.A(\inputs.random_update_clock.count[20] ),
    .B(\inputs.random_update_clock.count[22] ),
    .C_N(\inputs.random_update_clock.count[21] ),
    .Y(_0949_));
 sky130_fd_sc_hd__and4_1 _1307_ (.A(_0944_),
    .B(_0947_),
    .C(_0948_),
    .D(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__clkbuf_4 _1308_ (.A(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__nor3_1 _1309_ (.A(_0940_),
    .B(_0941_),
    .C(_0951_),
    .Y(\inputs.random_update_clock.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _1310_ (.A(\inputs.random_update_clock.count[6] ),
    .B(_0941_),
    .X(_0952_));
 sky130_fd_sc_hd__nor2_1 _1311_ (.A(net237),
    .B(_0941_),
    .Y(_0953_));
 sky130_fd_sc_hd__nor2_1 _1312_ (.A(_0952_),
    .B(_0953_),
    .Y(\inputs.random_update_clock.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _1313_ (.A(\inputs.random_update_clock.count[6] ),
    .B(\inputs.random_update_clock.count[7] ),
    .C(_0941_),
    .X(_0954_));
 sky130_fd_sc_hd__nand4_2 _1314_ (.A(_0944_),
    .B(_0947_),
    .C(_0948_),
    .D(_0949_),
    .Y(_0955_));
 sky130_fd_sc_hd__o21ai_1 _1315_ (.A1(net247),
    .A2(_0952_),
    .B1(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__nor2_1 _1316_ (.A(_0954_),
    .B(_0956_),
    .Y(\inputs.random_update_clock.next_count[7] ));
 sky130_fd_sc_hd__nor2_1 _1317_ (.A(\inputs.random_update_clock.count[8] ),
    .B(_0954_),
    .Y(_0957_));
 sky130_fd_sc_hd__and2_1 _1318_ (.A(\inputs.random_update_clock.count[8] ),
    .B(_0954_),
    .X(_0958_));
 sky130_fd_sc_hd__nor3_1 _1319_ (.A(_0951_),
    .B(_0957_),
    .C(_0958_),
    .Y(\inputs.random_update_clock.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _1320_ (.A(\inputs.random_update_clock.count[9] ),
    .B(\inputs.random_update_clock.count[8] ),
    .C(_0954_),
    .X(_0959_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(net213),
    .B(_0958_),
    .Y(_0960_));
 sky130_fd_sc_hd__nor2_1 _1322_ (.A(_0959_),
    .B(_0960_),
    .Y(\inputs.random_update_clock.next_count[9] ));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(\inputs.random_update_clock.count[10] ),
    .B(_0959_),
    .Y(_0961_));
 sky130_fd_sc_hd__or2_1 _1324_ (.A(\inputs.random_update_clock.count[10] ),
    .B(_0959_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_1 _1325_ (.A(_0955_),
    .B(_0961_),
    .C(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_1 _1326_ (.A(_0963_),
    .X(\inputs.random_update_clock.next_count[10] ));
 sky130_fd_sc_hd__xnor2_1 _1327_ (.A(net221),
    .B(_0961_),
    .Y(\inputs.random_update_clock.next_count[11] ));
 sky130_fd_sc_hd__and4_1 _1328_ (.A(\inputs.random_update_clock.count[11] ),
    .B(\inputs.random_update_clock.count[10] ),
    .C(\inputs.random_update_clock.count[12] ),
    .D(_0959_),
    .X(_0964_));
 sky130_fd_sc_hd__a31o_1 _1329_ (.A1(\inputs.random_update_clock.count[11] ),
    .A2(\inputs.random_update_clock.count[10] ),
    .A3(_0959_),
    .B1(\inputs.random_update_clock.count[12] ),
    .X(_0965_));
 sky130_fd_sc_hd__and2b_1 _1330_ (.A_N(_0964_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_1 _1331_ (.A(_0966_),
    .X(\inputs.random_update_clock.next_count[12] ));
 sky130_fd_sc_hd__or2_1 _1332_ (.A(\inputs.random_update_clock.count[13] ),
    .B(_0964_),
    .X(_0967_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(\inputs.random_update_clock.count[13] ),
    .B(_0964_),
    .Y(_0968_));
 sky130_fd_sc_hd__and3_1 _1334_ (.A(_0955_),
    .B(_0967_),
    .C(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_1 _1335_ (.A(_0969_),
    .X(\inputs.random_update_clock.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _1336_ (.A(\inputs.random_update_clock.count[13] ),
    .B(\inputs.random_update_clock.count[14] ),
    .C(_0964_),
    .X(_0970_));
 sky130_fd_sc_hd__a21oi_1 _1337_ (.A1(\inputs.random_update_clock.count[13] ),
    .A2(_0964_),
    .B1(net185),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_1 _1338_ (.A(_0970_),
    .B(net186),
    .Y(\inputs.random_update_clock.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _1339_ (.A(\inputs.random_update_clock.count[15] ),
    .B(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_1 _1340_ (.A(net227),
    .B(_0970_),
    .Y(_0973_));
 sky130_fd_sc_hd__nor2_1 _1341_ (.A(_0972_),
    .B(_0973_),
    .Y(\inputs.random_update_clock.next_count[15] ));
 sky130_fd_sc_hd__xor2_1 _1342_ (.A(net206),
    .B(_0972_),
    .X(\inputs.random_update_clock.next_count[16] ));
 sky130_fd_sc_hd__a21oi_1 _1343_ (.A1(\inputs.random_update_clock.count[16] ),
    .A2(_0972_),
    .B1(net293),
    .Y(_0974_));
 sky130_fd_sc_hd__and3_1 _1344_ (.A(\inputs.random_update_clock.count[16] ),
    .B(\inputs.random_update_clock.count[17] ),
    .C(_0972_),
    .X(_0975_));
 sky130_fd_sc_hd__nor3_1 _1345_ (.A(_0951_),
    .B(_0974_),
    .C(_0975_),
    .Y(\inputs.random_update_clock.next_count[17] ));
 sky130_fd_sc_hd__nor2_1 _1346_ (.A(\inputs.random_update_clock.count[18] ),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__and2_1 _1347_ (.A(\inputs.random_update_clock.count[18] ),
    .B(_0975_),
    .X(_0977_));
 sky130_fd_sc_hd__nor3_1 _1348_ (.A(_0951_),
    .B(_0976_),
    .C(_0977_),
    .Y(\inputs.random_update_clock.next_count[18] ));
 sky130_fd_sc_hd__xor2_1 _1349_ (.A(net218),
    .B(_0977_),
    .X(\inputs.random_update_clock.next_count[19] ));
 sky130_fd_sc_hd__and3_1 _1350_ (.A(\inputs.random_update_clock.count[19] ),
    .B(\inputs.random_update_clock.count[20] ),
    .C(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__a21oi_1 _1351_ (.A1(net218),
    .A2(_0977_),
    .B1(net226),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_1 _1352_ (.A(_0978_),
    .B(_0979_),
    .Y(\inputs.random_update_clock.next_count[20] ));
 sky130_fd_sc_hd__or2_1 _1353_ (.A(\inputs.random_update_clock.count[21] ),
    .B(_0978_),
    .X(_0980_));
 sky130_fd_sc_hd__nand2_1 _1354_ (.A(\inputs.random_update_clock.count[21] ),
    .B(_0978_),
    .Y(_0981_));
 sky130_fd_sc_hd__and3_1 _1355_ (.A(_0955_),
    .B(_0980_),
    .C(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__clkbuf_1 _1356_ (.A(_0982_),
    .X(\inputs.random_update_clock.next_count[21] ));
 sky130_fd_sc_hd__xnor2_1 _1357_ (.A(net118),
    .B(_0981_),
    .Y(\inputs.random_update_clock.next_count[22] ));
 sky130_fd_sc_hd__nor3b_1 _1358_ (.A(net146),
    .B(net92),
    .C_N(\inputs.key_encoder.sync_keys[14] ),
    .Y(\inputs.key_encoder.mode_key ));
 sky130_fd_sc_hd__and2b_1 _1359_ (.A_N(\inputs.key_encoder.octave_key_up ),
    .B(\inputs.key_encoder.sync_keys[15] ),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _1360_ (.A(_0983_),
    .X(\inputs.down.in ));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(net100),
    .Y(\outputs.output_gen.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1362_ (.A(net153),
    .B(net100),
    .X(\outputs.output_gen.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _1363_ (.A(\outputs.output_gen.count[2] ),
    .B(\outputs.output_gen.count[1] ),
    .C(\outputs.output_gen.count[0] ),
    .X(_0984_));
 sky130_fd_sc_hd__a21oi_1 _1364_ (.A1(\outputs.output_gen.count[1] ),
    .A2(net100),
    .B1(net241),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_1 _1365_ (.A(_0984_),
    .B(net242),
    .Y(\outputs.output_gen.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _1366_ (.A(\outputs.output_gen.count[3] ),
    .B(_0984_),
    .X(_0986_));
 sky130_fd_sc_hd__nor2_1 _1367_ (.A(net261),
    .B(_0984_),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_1 _1368_ (.A(_0986_),
    .B(_0987_),
    .Y(\outputs.output_gen.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1369_ (.A(net245),
    .B(_0986_),
    .X(\outputs.output_gen.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1370_ (.A(\outputs.output_gen.count[5] ),
    .B(\outputs.output_gen.count[4] ),
    .C(_0986_),
    .X(_0988_));
 sky130_fd_sc_hd__a21oi_1 _1371_ (.A1(\outputs.output_gen.count[4] ),
    .A2(_0986_),
    .B1(net249),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_0988_),
    .B(net250),
    .Y(\outputs.output_gen.next_count[5] ));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(\outputs.output_gen.count[6] ),
    .B(_0988_),
    .Y(_0990_));
 sky130_fd_sc_hd__or2_1 _1374_ (.A(\outputs.output_gen.count[6] ),
    .B(_0988_),
    .X(_0991_));
 sky130_fd_sc_hd__and2_1 _1375_ (.A(_0990_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(_0992_),
    .X(\outputs.output_gen.next_count[6] ));
 sky130_fd_sc_hd__xnor2_1 _1377_ (.A(net177),
    .B(_0990_),
    .Y(\outputs.output_gen.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _1378_ (.A(\outputs.sample_rate.count[6] ),
    .B(\outputs.sample_rate.count[7] ),
    .C(_0908_),
    .X(_0993_));
 sky130_fd_sc_hd__buf_4 _1379_ (.A(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nor2_1 _1380_ (.A(_0994_),
    .B(_0913_),
    .Y(_0995_));
 sky130_fd_sc_hd__clkbuf_4 _1381_ (.A(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_4 _1382_ (.A(_0996_),
    .X(\outputs.div.next_div ));
 sky130_fd_sc_hd__inv_2 _1383_ (.A(net133),
    .Y(\outputs.sample_rate.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _1384_ (.A(net148),
    .B(net133),
    .X(\outputs.sample_rate.next_count[1] ));
 sky130_fd_sc_hd__a21oi_1 _1385_ (.A1(net148),
    .A2(\outputs.sample_rate.count[0] ),
    .B1(net156),
    .Y(_0997_));
 sky130_fd_sc_hd__nor2_1 _1386_ (.A(_0906_),
    .B(net157),
    .Y(\outputs.sample_rate.next_count[2] ));
 sky130_fd_sc_hd__nor2_1 _1387_ (.A(net152),
    .B(_0906_),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _1388_ (.A(_0907_),
    .B(_0998_),
    .Y(\outputs.sample_rate.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _1389_ (.A(net145),
    .B(_0907_),
    .X(\outputs.sample_rate.next_count[4] ));
 sky130_fd_sc_hd__a21oi_1 _1390_ (.A1(\outputs.sample_rate.count[4] ),
    .A2(_0907_),
    .B1(net139),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _1391_ (.A(_0908_),
    .B(net140),
    .Y(\outputs.sample_rate.next_count[5] ));
 sky130_fd_sc_hd__nor2_1 _1392_ (.A(net223),
    .B(_0908_),
    .Y(_1000_));
 sky130_fd_sc_hd__nor2_1 _1393_ (.A(_0909_),
    .B(_1000_),
    .Y(\outputs.sample_rate.next_count[6] ));
 sky130_fd_sc_hd__buf_4 _1394_ (.A(_0994_),
    .X(_1001_));
 sky130_fd_sc_hd__nor2_1 _1395_ (.A(net303),
    .B(_0909_),
    .Y(_1002_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(_1001_),
    .B(_1002_),
    .Y(\outputs.sample_rate.next_count[7] ));
 sky130_fd_sc_hd__inv_2 _1397_ (.A(\outputs.divider_buffer[1] ),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(\outputs.sig_gen.count[13] ),
    .Y(_1004_));
 sky130_fd_sc_hd__a2bb2o_1 _1399_ (.A1_N(_1003_),
    .A2_N(\outputs.sig_gen.count[1] ),
    .B1(\outputs.divider_buffer[13] ),
    .B2(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__inv_2 _1400_ (.A(\outputs.divider_buffer[9] ),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_2 _1401_ (.A(\outputs.divider_buffer[17] ),
    .Y(_1007_));
 sky130_fd_sc_hd__xor2_1 _1402_ (.A(\outputs.divider_buffer[12] ),
    .B(\outputs.sig_gen.count[12] ),
    .X(_1008_));
 sky130_fd_sc_hd__a221o_1 _1403_ (.A1(_1006_),
    .A2(\outputs.sig_gen.count[9] ),
    .B1(_1007_),
    .B2(\outputs.sig_gen.count[17] ),
    .C1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__inv_2 _1404_ (.A(\outputs.sig_gen.count[3] ),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_2 _1405_ (.A(\outputs.sig_gen.count[9] ),
    .Y(_1011_));
 sky130_fd_sc_hd__xor2_1 _1406_ (.A(\outputs.divider_buffer[4] ),
    .B(\outputs.sig_gen.count[4] ),
    .X(_1012_));
 sky130_fd_sc_hd__a221o_1 _1407_ (.A1(\outputs.divider_buffer[3] ),
    .A2(_1010_),
    .B1(\outputs.divider_buffer[9] ),
    .B2(_1011_),
    .C1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__inv_2 _1408_ (.A(\outputs.divider_buffer[10] ),
    .Y(_1014_));
 sky130_fd_sc_hd__a2bb2o_1 _1409_ (.A1_N(_1014_),
    .A2_N(\outputs.sig_gen.count[10] ),
    .B1(_1003_),
    .B2(\outputs.sig_gen.count[1] ),
    .X(_1015_));
 sky130_fd_sc_hd__or4_1 _1410_ (.A(_1005_),
    .B(_1009_),
    .C(_1013_),
    .D(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__inv_2 _1411_ (.A(\outputs.divider_buffer[3] ),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_2 _1412_ (.A(\outputs.divider_buffer[15] ),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_2 _1413_ (.A(\outputs.divider_buffer[5] ),
    .Y(_1019_));
 sky130_fd_sc_hd__o22ai_1 _1414_ (.A1(_1019_),
    .A2(\outputs.sig_gen.count[5] ),
    .B1(_1007_),
    .B2(\outputs.sig_gen.count[17] ),
    .Y(_1020_));
 sky130_fd_sc_hd__a221o_1 _1415_ (.A1(_1017_),
    .A2(\outputs.sig_gen.count[3] ),
    .B1(_1018_),
    .B2(\outputs.sig_gen.count[15] ),
    .C1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(\outputs.divider_buffer[14] ),
    .Y(_1022_));
 sky130_fd_sc_hd__inv_2 _1417_ (.A(\outputs.sig_gen.count[16] ),
    .Y(_1023_));
 sky130_fd_sc_hd__xor2_1 _1418_ (.A(\outputs.divider_buffer[2] ),
    .B(\outputs.sig_gen.count[2] ),
    .X(_1024_));
 sky130_fd_sc_hd__a221o_1 _1419_ (.A1(_1022_),
    .A2(\outputs.sig_gen.count[14] ),
    .B1(\outputs.divider_buffer[16] ),
    .B2(_1023_),
    .C1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__inv_2 _1420_ (.A(\outputs.sig_gen.count[7] ),
    .Y(_1026_));
 sky130_fd_sc_hd__inv_2 _1421_ (.A(\outputs.sig_gen.count[11] ),
    .Y(_1027_));
 sky130_fd_sc_hd__xor2_1 _1422_ (.A(\outputs.divider_buffer[8] ),
    .B(\outputs.sig_gen.count[8] ),
    .X(_1028_));
 sky130_fd_sc_hd__a221o_1 _1423_ (.A1(\outputs.divider_buffer[7] ),
    .A2(_1026_),
    .B1(\outputs.divider_buffer[11] ),
    .B2(_1027_),
    .C1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__inv_2 _1424_ (.A(\outputs.divider_buffer[6] ),
    .Y(_1030_));
 sky130_fd_sc_hd__o22a_1 _1425_ (.A1(_1030_),
    .A2(\outputs.sig_gen.count[6] ),
    .B1(\outputs.divider_buffer[16] ),
    .B2(_1023_),
    .X(_1031_));
 sky130_fd_sc_hd__o221ai_1 _1426_ (.A1(\outputs.divider_buffer[13] ),
    .A2(_1004_),
    .B1(_1022_),
    .B2(\outputs.sig_gen.count[14] ),
    .C1(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__inv_2 _1427_ (.A(\outputs.divider_buffer[0] ),
    .Y(_1033_));
 sky130_fd_sc_hd__inv_2 _1428_ (.A(\outputs.divider_buffer[11] ),
    .Y(_1034_));
 sky130_fd_sc_hd__a2bb2o_1 _1429_ (.A1_N(_1033_),
    .A2_N(\outputs.sig_gen.count[0] ),
    .B1(_1019_),
    .B2(\outputs.sig_gen.count[5] ),
    .X(_1035_));
 sky130_fd_sc_hd__a221o_1 _1430_ (.A1(_1033_),
    .A2(\outputs.sig_gen.count[0] ),
    .B1(_1034_),
    .B2(\outputs.sig_gen.count[11] ),
    .C1(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__inv_2 _1431_ (.A(\outputs.divider_buffer[7] ),
    .Y(_1037_));
 sky130_fd_sc_hd__a2bb2o_1 _1432_ (.A1_N(_1018_),
    .A2_N(\outputs.sig_gen.count[15] ),
    .B1(_1030_),
    .B2(\outputs.sig_gen.count[6] ),
    .X(_1038_));
 sky130_fd_sc_hd__a221o_1 _1433_ (.A1(_1037_),
    .A2(\outputs.sig_gen.count[7] ),
    .B1(_1014_),
    .B2(\outputs.sig_gen.count[10] ),
    .C1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__or4_1 _1434_ (.A(_1029_),
    .B(_1032_),
    .C(_1036_),
    .D(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__or4_4 _1435_ (.A(_1016_),
    .B(_1021_),
    .C(_1025_),
    .D(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__buf_2 _1436_ (.A(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(net248),
    .B(_1042_),
    .Y(\outputs.sig_gen.next_count[0] ));
 sky130_fd_sc_hd__or2_1 _1438_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .X(_1043_));
 sky130_fd_sc_hd__nand2_1 _1439_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .Y(_1044_));
 sky130_fd_sc_hd__and3_1 _1440_ (.A(_1042_),
    .B(_1043_),
    .C(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_1 _1441_ (.A(_1045_),
    .X(\outputs.sig_gen.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _1442_ (.A1(\outputs.sig_gen.count[0] ),
    .A2(\outputs.sig_gen.count[1] ),
    .B1(\outputs.sig_gen.count[2] ),
    .X(_1046_));
 sky130_fd_sc_hd__nand3_1 _1443_ (.A(\outputs.sig_gen.count[0] ),
    .B(\outputs.sig_gen.count[1] ),
    .C(\outputs.sig_gen.count[2] ),
    .Y(_1047_));
 sky130_fd_sc_hd__and3_1 _1444_ (.A(_1041_),
    .B(_1046_),
    .C(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_1 _1445_ (.A(_1048_),
    .X(\outputs.sig_gen.next_count[2] ));
 sky130_fd_sc_hd__nor2_1 _1446_ (.A(_1010_),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__inv_2 _1447_ (.A(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2_1 _1448_ (.A(_1010_),
    .B(_1047_),
    .Y(_1051_));
 sky130_fd_sc_hd__and3_1 _1449_ (.A(_1041_),
    .B(_1050_),
    .C(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(_1052_),
    .X(\outputs.sig_gen.next_count[3] ));
 sky130_fd_sc_hd__and2_1 _1451_ (.A(\outputs.sig_gen.count[4] ),
    .B(_1049_),
    .X(_1053_));
 sky130_fd_sc_hd__o21ai_1 _1452_ (.A1(\outputs.sig_gen.count[4] ),
    .A2(_1049_),
    .B1(_1042_),
    .Y(_1054_));
 sky130_fd_sc_hd__nor2_1 _1453_ (.A(_1053_),
    .B(_1054_),
    .Y(\outputs.sig_gen.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _1454_ (.A(\outputs.sig_gen.count[4] ),
    .B(\outputs.sig_gen.count[5] ),
    .C(_1049_),
    .X(_1055_));
 sky130_fd_sc_hd__o21ai_1 _1455_ (.A1(net307),
    .A2(_1053_),
    .B1(_1042_),
    .Y(_1056_));
 sky130_fd_sc_hd__nor2_1 _1456_ (.A(_1055_),
    .B(_1056_),
    .Y(\outputs.sig_gen.next_count[5] ));
 sky130_fd_sc_hd__or2_1 _1457_ (.A(\outputs.sig_gen.count[6] ),
    .B(_1055_),
    .X(_1057_));
 sky130_fd_sc_hd__and2_1 _1458_ (.A(\outputs.sig_gen.count[6] ),
    .B(_1055_),
    .X(_1058_));
 sky130_fd_sc_hd__inv_2 _1459_ (.A(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__and3_1 _1460_ (.A(_1041_),
    .B(_1057_),
    .C(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _1461_ (.A(_1060_),
    .X(\outputs.sig_gen.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _1462_ (.A(\outputs.sig_gen.count[6] ),
    .B(\outputs.sig_gen.count[7] ),
    .C(_1055_),
    .X(_1061_));
 sky130_fd_sc_hd__o21ai_1 _1463_ (.A1(\outputs.sig_gen.count[7] ),
    .A2(_1058_),
    .B1(_1042_),
    .Y(_1062_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_1061_),
    .B(_1062_),
    .Y(\outputs.sig_gen.next_count[7] ));
 sky130_fd_sc_hd__or2_1 _1465_ (.A(\outputs.sig_gen.count[8] ),
    .B(_1061_),
    .X(_1063_));
 sky130_fd_sc_hd__and2_1 _1466_ (.A(\outputs.sig_gen.count[8] ),
    .B(_1061_),
    .X(_1064_));
 sky130_fd_sc_hd__inv_2 _1467_ (.A(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__and3_1 _1468_ (.A(_1041_),
    .B(_1063_),
    .C(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _1469_ (.A(_1066_),
    .X(\outputs.sig_gen.next_count[8] ));
 sky130_fd_sc_hd__or2_1 _1470_ (.A(\outputs.sig_gen.count[9] ),
    .B(_1064_),
    .X(_1067_));
 sky130_fd_sc_hd__o211a_1 _1471_ (.A1(_1011_),
    .A2(_1065_),
    .B1(_1067_),
    .C1(_1042_),
    .X(\outputs.sig_gen.next_count[9] ));
 sky130_fd_sc_hd__nor2_1 _1472_ (.A(_1011_),
    .B(_1065_),
    .Y(_1068_));
 sky130_fd_sc_hd__or2_1 _1473_ (.A(\outputs.sig_gen.count[10] ),
    .B(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(\outputs.sig_gen.count[10] ),
    .B(_1068_),
    .Y(_1070_));
 sky130_fd_sc_hd__and3_1 _1475_ (.A(_1041_),
    .B(_1069_),
    .C(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _1476_ (.A(_1071_),
    .X(\outputs.sig_gen.next_count[10] ));
 sky130_fd_sc_hd__nand2_1 _1477_ (.A(_1027_),
    .B(_1070_),
    .Y(_1072_));
 sky130_fd_sc_hd__o211a_1 _1478_ (.A1(_1027_),
    .A2(_1070_),
    .B1(_1072_),
    .C1(_1042_),
    .X(\outputs.sig_gen.next_count[11] ));
 sky130_fd_sc_hd__nor2_1 _1479_ (.A(_1027_),
    .B(_1070_),
    .Y(_1073_));
 sky130_fd_sc_hd__or2_1 _1480_ (.A(\outputs.sig_gen.count[12] ),
    .B(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _1481_ (.A(\outputs.sig_gen.count[12] ),
    .B(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__inv_2 _1482_ (.A(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__and3_1 _1483_ (.A(_1041_),
    .B(_1074_),
    .C(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _1484_ (.A(_1077_),
    .X(\outputs.sig_gen.next_count[12] ));
 sky130_fd_sc_hd__or2_1 _1485_ (.A(\outputs.sig_gen.count[13] ),
    .B(_1075_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(\outputs.sig_gen.count[13] ),
    .B(_1075_),
    .Y(_1079_));
 sky130_fd_sc_hd__and3_1 _1487_ (.A(_1041_),
    .B(_1078_),
    .C(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _1488_ (.A(_1080_),
    .X(\outputs.sig_gen.next_count[13] ));
 sky130_fd_sc_hd__inv_2 _1489_ (.A(\outputs.sig_gen.count[14] ),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(_1081_),
    .B(_1079_),
    .Y(_1082_));
 sky130_fd_sc_hd__o211a_1 _1491_ (.A1(_1081_),
    .A2(_1079_),
    .B1(_1082_),
    .C1(_1042_),
    .X(\outputs.sig_gen.next_count[14] ));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(_1081_),
    .B(_1079_),
    .Y(_1083_));
 sky130_fd_sc_hd__or2_1 _1493_ (.A(\outputs.sig_gen.count[15] ),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(\outputs.sig_gen.count[15] ),
    .B(_1083_),
    .Y(_1085_));
 sky130_fd_sc_hd__and3_1 _1495_ (.A(_1041_),
    .B(_1084_),
    .C(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_1086_),
    .X(\outputs.sig_gen.next_count[15] ));
 sky130_fd_sc_hd__nand2_1 _1497_ (.A(_1023_),
    .B(_1085_),
    .Y(_1087_));
 sky130_fd_sc_hd__o211a_1 _1498_ (.A1(_1023_),
    .A2(_1085_),
    .B1(_1087_),
    .C1(_1042_),
    .X(\outputs.sig_gen.next_count[16] ));
 sky130_fd_sc_hd__nor2_1 _1499_ (.A(_1023_),
    .B(_1085_),
    .Y(_1088_));
 sky130_fd_sc_hd__o21ai_1 _1500_ (.A1(net207),
    .A2(_1088_),
    .B1(_1042_),
    .Y(_1089_));
 sky130_fd_sc_hd__a21oi_1 _1501_ (.A1(net207),
    .A2(_1088_),
    .B1(_1089_),
    .Y(\outputs.sig_gen.next_count[17] ));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(net254),
    .Y(_1090_));
 sky130_fd_sc_hd__or2_1 _1503_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.mode_edge.det_edge ),
    .X(_1091_));
 sky130_fd_sc_hd__and2_1 _1504_ (.A(_1090_),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__clkbuf_1 _1505_ (.A(_1092_),
    .X(\inputs.wavetype_fsm.next_state[0] ));
 sky130_fd_sc_hd__xnor2_1 _1506_ (.A(\inputs.wavetype_fsm.state[1] ),
    .B(_1090_),
    .Y(\inputs.wavetype_fsm.next_state[1] ));
 sky130_fd_sc_hd__buf_2 _1507_ (.A(\inputs.random_note_generator.out[15] ),
    .X(_1093_));
 sky130_fd_sc_hd__xor2_1 _1508_ (.A(_1093_),
    .B(\inputs.random_note_generator.out[13] ),
    .X(_1094_));
 sky130_fd_sc_hd__xor2_1 _1509_ (.A(net88),
    .B(\inputs.random_note_generator.out[10] ),
    .X(_1095_));
 sky130_fd_sc_hd__xnor2_1 _1510_ (.A(_1094_),
    .B(_1095_),
    .Y(\inputs.random_note_generator.feedback ));
 sky130_fd_sc_hd__or2b_1 _1511_ (.A(net149),
    .B_N(\inputs.key_encoder.mode_key ),
    .X(_1096_));
 sky130_fd_sc_hd__inv_2 _1512_ (.A(_1096_),
    .Y(\inputs.mode_edge.ff_in ));
 sky130_fd_sc_hd__and2b_1 _1513_ (.A_N(\inputs.down.ff_out ),
    .B(\inputs.down.in ),
    .X(_1097_));
 sky130_fd_sc_hd__clkbuf_1 _1514_ (.A(_1097_),
    .X(\inputs.down.ff_in ));
 sky130_fd_sc_hd__and2b_1 _1515_ (.A_N(\inputs.up.ff_out ),
    .B(\inputs.key_encoder.octave_key_up ),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _1516_ (.A(_1098_),
    .X(\inputs.up.ff_in ));
 sky130_fd_sc_hd__or4_2 _1517_ (.A(\outputs.scaled_buffer[0] ),
    .B(\outputs.scaled_buffer[1] ),
    .C(\outputs.scaled_buffer[3] ),
    .D(\outputs.scaled_buffer[2] ),
    .X(_1099_));
 sky130_fd_sc_hd__and2_1 _1518_ (.A(_1022_),
    .B(\outputs.shaper.count[13] ),
    .X(_1100_));
 sky130_fd_sc_hd__inv_2 _1519_ (.A(\outputs.shaper.count[14] ),
    .Y(_1101_));
 sky130_fd_sc_hd__nor2_1 _1520_ (.A(\outputs.divider_buffer[15] ),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__inv_2 _1521_ (.A(\outputs.divider_buffer[16] ),
    .Y(_1103_));
 sky130_fd_sc_hd__a2bb2o_1 _1522_ (.A1_N(_1103_),
    .A2_N(\outputs.shaper.count[15] ),
    .B1(_1101_),
    .B2(\outputs.divider_buffer[15] ),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_1103_),
    .B(\outputs.shaper.count[15] ),
    .Y(_1105_));
 sky130_fd_sc_hd__or3b_1 _1524_ (.A(_1102_),
    .B(_1104_),
    .C_N(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__inv_2 _1525_ (.A(\outputs.shaper.count[9] ),
    .Y(_1107_));
 sky130_fd_sc_hd__a2bb2o_1 _1526_ (.A1_N(_1006_),
    .A2_N(\outputs.shaper.count[8] ),
    .B1(\outputs.divider_buffer[10] ),
    .B2(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a21o_1 _1527_ (.A1(_1006_),
    .A2(\outputs.shaper.count[8] ),
    .B1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__inv_2 _1528_ (.A(\outputs.shaper.count[12] ),
    .Y(_1110_));
 sky130_fd_sc_hd__a2bb2o_1 _1529_ (.A1_N(_1022_),
    .A2_N(\outputs.shaper.count[13] ),
    .B1(_1110_),
    .B2(\outputs.divider_buffer[13] ),
    .X(_1111_));
 sky130_fd_sc_hd__inv_2 _1530_ (.A(\outputs.shaper.count[11] ),
    .Y(_1112_));
 sky130_fd_sc_hd__inv_2 _1531_ (.A(\outputs.shaper.count[10] ),
    .Y(_1113_));
 sky130_fd_sc_hd__a22o_1 _1532_ (.A1(\outputs.divider_buffer[12] ),
    .A2(_1112_),
    .B1(_1113_),
    .B2(\outputs.divider_buffer[11] ),
    .X(_1114_));
 sky130_fd_sc_hd__nor2_1 _1533_ (.A(\outputs.divider_buffer[10] ),
    .B(_1107_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(\outputs.divider_buffer[11] ),
    .B(_1113_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(\outputs.divider_buffer[12] ),
    .B(_1112_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor2_1 _1536_ (.A(\outputs.divider_buffer[13] ),
    .B(_1110_),
    .Y(_1118_));
 sky130_fd_sc_hd__or4_1 _1537_ (.A(_1115_),
    .B(_1116_),
    .C(_1117_),
    .D(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__or4_1 _1538_ (.A(_1109_),
    .B(_1111_),
    .C(_1114_),
    .D(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__or3_1 _1539_ (.A(_1100_),
    .B(_1106_),
    .C(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__inv_2 _1540_ (.A(\outputs.shaper.count[7] ),
    .Y(_1122_));
 sky130_fd_sc_hd__or2_1 _1541_ (.A(\outputs.divider_buffer[8] ),
    .B(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__inv_2 _1542_ (.A(\outputs.shaper.count[3] ),
    .Y(_1124_));
 sky130_fd_sc_hd__inv_2 _1543_ (.A(\outputs.shaper.count[2] ),
    .Y(_1125_));
 sky130_fd_sc_hd__a22o_1 _1544_ (.A1(\outputs.divider_buffer[4] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\outputs.divider_buffer[3] ),
    .X(_1126_));
 sky130_fd_sc_hd__or2b_1 _1545_ (.A(\outputs.shaper.count[1] ),
    .B_N(\outputs.divider_buffer[2] ),
    .X(_1127_));
 sky130_fd_sc_hd__inv_2 _1546_ (.A(\outputs.shaper.count[0] ),
    .Y(_1128_));
 sky130_fd_sc_hd__or2b_1 _1547_ (.A(\outputs.divider_buffer[2] ),
    .B_N(\outputs.shaper.count[1] ),
    .X(_1129_));
 sky130_fd_sc_hd__o211ai_1 _1548_ (.A1(\outputs.divider_buffer[1] ),
    .A2(_1128_),
    .B1(_1127_),
    .C1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nor2_1 _1549_ (.A(\outputs.divider_buffer[3] ),
    .B(_1125_),
    .Y(_1131_));
 sky130_fd_sc_hd__a21oi_1 _1550_ (.A1(_1127_),
    .A2(_1130_),
    .B1(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__or2_1 _1551_ (.A(_1126_),
    .B(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or2_1 _1552_ (.A(\outputs.divider_buffer[4] ),
    .B(_1124_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _1553_ (.A(_1019_),
    .B(\outputs.shaper.count[4] ),
    .Y(_1135_));
 sky130_fd_sc_hd__o22ai_2 _1554_ (.A1(_1030_),
    .A2(\outputs.shaper.count[5] ),
    .B1(\outputs.shaper.count[4] ),
    .B2(_1019_),
    .Y(_1136_));
 sky130_fd_sc_hd__a31o_1 _1555_ (.A1(_1133_),
    .A2(_1134_),
    .A3(_1135_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__nand2_1 _1556_ (.A(_1030_),
    .B(\outputs.shaper.count[5] ),
    .Y(_1138_));
 sky130_fd_sc_hd__nand2_1 _1557_ (.A(_1037_),
    .B(\outputs.shaper.count[6] ),
    .Y(_1139_));
 sky130_fd_sc_hd__a2bb2o_1 _1558_ (.A1_N(_1037_),
    .A2_N(\outputs.shaper.count[6] ),
    .B1(\outputs.divider_buffer[8] ),
    .B2(_1122_),
    .X(_1140_));
 sky130_fd_sc_hd__a31o_1 _1559_ (.A1(_1137_),
    .A2(_1138_),
    .A3(_1139_),
    .B1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__and3b_1 _1560_ (.A_N(_1121_),
    .B(_1123_),
    .C(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__nor2_1 _1561_ (.A(_1115_),
    .B(_1116_),
    .Y(_1143_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(_1108_),
    .A2(_1143_),
    .B1(_1114_),
    .Y(_1144_));
 sky130_fd_sc_hd__inv_2 _1563_ (.A(_1111_),
    .Y(_1145_));
 sky130_fd_sc_hd__o31a_1 _1564_ (.A1(_1117_),
    .A2(_1118_),
    .A3(_1144_),
    .B1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__o2bb2a_1 _1565_ (.A1_N(_1104_),
    .A2_N(_1105_),
    .B1(_1007_),
    .B2(\outputs.shaper.count[16] ),
    .X(_1147_));
 sky130_fd_sc_hd__o31ai_2 _1566_ (.A1(_1100_),
    .A2(_1106_),
    .A3(_1146_),
    .B1(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__a21oi_1 _1567_ (.A1(_1007_),
    .A2(\outputs.shaper.count[16] ),
    .B1(\outputs.shaper.count[17] ),
    .Y(_1149_));
 sky130_fd_sc_hd__or4b_1 _1568_ (.A(_1140_),
    .B(_1136_),
    .C(_1126_),
    .D_N(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__o22a_1 _1569_ (.A1(_1007_),
    .A2(\outputs.shaper.count[16] ),
    .B1(\outputs.shaper.count[0] ),
    .B2(_1003_),
    .X(_1151_));
 sky130_fd_sc_hd__and4b_1 _1570_ (.A_N(_1131_),
    .B(_1134_),
    .C(_1139_),
    .D(_1123_),
    .X(_1152_));
 sky130_fd_sc_hd__and4_1 _1571_ (.A(_1135_),
    .B(_1138_),
    .C(_1151_),
    .D(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__or4b_1 _1572_ (.A(_1130_),
    .B(_1121_),
    .C(_1150_),
    .D_N(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__o211ai_2 _1573_ (.A1(_1142_),
    .A2(_1148_),
    .B1(_1149_),
    .C1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__a21oi_1 _1574_ (.A1(_1099_),
    .A2(net21),
    .B1(\outputs.scaled_buffer[4] ),
    .Y(_1156_));
 sky130_fd_sc_hd__nor2b_2 _1575_ (.A(\inputs.wavetype_fsm.state[1] ),
    .B_N(\inputs.wavetype_fsm.state[0] ),
    .Y(_1157_));
 sky130_fd_sc_hd__inv_2 _1576_ (.A(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__a31o_1 _1577_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1099_),
    .A3(net21),
    .B1(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__and2b_1 _1578_ (.A_N(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.wavetype_fsm.state[1] ),
    .X(_1160_));
 sky130_fd_sc_hd__buf_2 _1579_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_1 _1580_ (.A(\inputs.wavetype_fsm.state[0] ),
    .B(\inputs.wavetype_fsm.state[1] ),
    .Y(_1162_));
 sky130_fd_sc_hd__or3_1 _1581_ (.A(\outputs.scaled_buffer[5] ),
    .B(\outputs.scaled_buffer[4] ),
    .C(_1099_),
    .X(_1163_));
 sky130_fd_sc_hd__or4b_2 _1582_ (.A(\outputs.scaled_buffer[6] ),
    .B(_1158_),
    .C(_1163_),
    .D_N(\outputs.scaled_buffer[7] ),
    .X(_1164_));
 sky130_fd_sc_hd__o21ai_4 _1583_ (.A1(net21),
    .A2(_1162_),
    .B1(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21oi_1 _1584_ (.A1(\outputs.scaled_buffer[5] ),
    .A2(_1161_),
    .B1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__o21a_1 _1585_ (.A1(_1156_),
    .A2(_1159_),
    .B1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__o21ai_1 _1586_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .B1(net21),
    .Y(_1168_));
 sky130_fd_sc_hd__xnor2_1 _1587_ (.A(\outputs.scaled_buffer[2] ),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__a221oi_2 _1588_ (.A1(\outputs.scaled_buffer[3] ),
    .A2(_1161_),
    .B1(_1169_),
    .B2(_1157_),
    .C1(_1165_),
    .Y(_1170_));
 sky130_fd_sc_hd__a21oi_1 _1589_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(net21),
    .B1(\outputs.scaled_buffer[1] ),
    .Y(_1171_));
 sky130_fd_sc_hd__a31o_1 _1590_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .A3(net21),
    .B1(_1158_),
    .X(_1172_));
 sky130_fd_sc_hd__a21oi_1 _1591_ (.A1(\outputs.scaled_buffer[2] ),
    .A2(_1161_),
    .B1(_1165_),
    .Y(_1173_));
 sky130_fd_sc_hd__o21a_1 _1592_ (.A1(_1171_),
    .A2(_1172_),
    .B1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__a221oi_2 _1593_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(_1157_),
    .B1(_1161_),
    .B2(\outputs.scaled_buffer[1] ),
    .C1(_1165_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_1 _1594_ (.A(\outputs.output_gen.count[1] ),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__a21oi_1 _1595_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(_1161_),
    .B1(_1165_),
    .Y(_1177_));
 sky130_fd_sc_hd__a211o_1 _1596_ (.A1(\outputs.output_gen.count[1] ),
    .A2(_1175_),
    .B1(_1177_),
    .C1(\outputs.output_gen.count[0] ),
    .X(_1178_));
 sky130_fd_sc_hd__a22o_1 _1597_ (.A1(\outputs.output_gen.count[2] ),
    .A2(_1174_),
    .B1(_1176_),
    .B2(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__o221a_1 _1598_ (.A1(\outputs.output_gen.count[3] ),
    .A2(_1170_),
    .B1(_1174_),
    .B2(\outputs.output_gen.count[2] ),
    .C1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__o31a_1 _1599_ (.A1(\outputs.scaled_buffer[0] ),
    .A2(\outputs.scaled_buffer[1] ),
    .A3(\outputs.scaled_buffer[2] ),
    .B1(net21),
    .X(_1181_));
 sky130_fd_sc_hd__xor2_1 _1600_ (.A(\outputs.scaled_buffer[3] ),
    .B(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a221oi_2 _1601_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1161_),
    .B1(_1182_),
    .B2(_1157_),
    .C1(_1165_),
    .Y(_1183_));
 sky130_fd_sc_hd__a22o_1 _1602_ (.A1(\outputs.output_gen.count[4] ),
    .A2(_1183_),
    .B1(_1170_),
    .B2(\outputs.output_gen.count[3] ),
    .X(_1184_));
 sky130_fd_sc_hd__or2_1 _1603_ (.A(\outputs.output_gen.count[4] ),
    .B(_1183_),
    .X(_1185_));
 sky130_fd_sc_hd__o221a_1 _1604_ (.A1(\outputs.output_gen.count[5] ),
    .A2(_1167_),
    .B1(_1180_),
    .B2(_1184_),
    .C1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__o21ai_1 _1605_ (.A1(\outputs.scaled_buffer[4] ),
    .A2(_1099_),
    .B1(net21),
    .Y(_1187_));
 sky130_fd_sc_hd__xnor2_1 _1606_ (.A(\outputs.scaled_buffer[5] ),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__a221oi_1 _1607_ (.A1(\outputs.scaled_buffer[6] ),
    .A2(_1161_),
    .B1(_1188_),
    .B2(_1157_),
    .C1(_1165_),
    .Y(_1189_));
 sky130_fd_sc_hd__a22o_1 _1608_ (.A1(\outputs.output_gen.count[5] ),
    .A2(_1167_),
    .B1(_1189_),
    .B2(\outputs.output_gen.count[6] ),
    .X(_1190_));
 sky130_fd_sc_hd__a21oi_1 _1609_ (.A1(net21),
    .A2(_1163_),
    .B1(\outputs.scaled_buffer[6] ),
    .Y(_1191_));
 sky130_fd_sc_hd__a31o_1 _1610_ (.A1(\outputs.scaled_buffer[6] ),
    .A2(net21),
    .A3(_1163_),
    .B1(_1158_),
    .X(_1192_));
 sky130_fd_sc_hd__a21oi_1 _1611_ (.A1(\outputs.scaled_buffer[7] ),
    .A2(_1161_),
    .B1(_1165_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21a_1 _1612_ (.A1(_1191_),
    .A2(_1192_),
    .B1(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _1613_ (.A(\outputs.output_gen.count[6] ),
    .B(_1189_),
    .X(_1195_));
 sky130_fd_sc_hd__o221a_1 _1614_ (.A1(_1186_),
    .A2(_1190_),
    .B1(_1194_),
    .B2(\outputs.output_gen.count[7] ),
    .C1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__nand2_1 _1615_ (.A(\outputs.output_gen.count[7] ),
    .B(_1194_),
    .Y(_1197_));
 sky130_fd_sc_hd__nor3_2 _1616_ (.A(\inputs.key_encoder.sync_keys[14] ),
    .B(\inputs.key_encoder.sync_keys[15] ),
    .C(\inputs.key_encoder.octave_key_up ),
    .Y(_1198_));
 sky130_fd_sc_hd__or4_4 _1617_ (.A(\inputs.key_encoder.sync_keys[11] ),
    .B(\inputs.key_encoder.sync_keys[8] ),
    .C(\inputs.key_encoder.sync_keys[9] ),
    .D(\inputs.key_encoder.sync_keys[10] ),
    .X(_1199_));
 sky130_fd_sc_hd__or2_1 _1618_ (.A(\inputs.key_encoder.sync_keys[2] ),
    .B(\inputs.key_encoder.sync_keys[3] ),
    .X(_1200_));
 sky130_fd_sc_hd__or4_1 _1619_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(\inputs.key_encoder.sync_keys[1] ),
    .C(\inputs.key_encoder.sync_keys[0] ),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__or4_1 _1620_ (.A(\inputs.key_encoder.sync_keys[4] ),
    .B(\inputs.key_encoder.sync_keys[5] ),
    .C(\inputs.key_encoder.sync_keys[6] ),
    .D(\inputs.key_encoder.sync_keys[7] ),
    .X(_1202_));
 sky130_fd_sc_hd__or4_1 _1621_ (.A(\inputs.key_encoder.sync_keys[12] ),
    .B(_1199_),
    .C(_1201_),
    .D(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__and4b_1 _1622_ (.A_N(_1196_),
    .B(_1197_),
    .C(_1198_),
    .D(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _1623_ (.A(_1204_),
    .X(\outputs.output_gen.pwm_unff ));
 sky130_fd_sc_hd__nor2_1 _1624_ (.A(\inputs.octave_fsm.state[1] ),
    .B(\inputs.octave_fsm.state[0] ),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _1625_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__clkbuf_4 _1626_ (.A(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__buf_2 _1627_ (.A(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__or2b_1 _1628_ (.A(\inputs.octave_fsm.state[2] ),
    .B_N(\inputs.octave_fsm.state[1] ),
    .X(_1209_));
 sky130_fd_sc_hd__and2b_2 _1629_ (.A_N(\inputs.down.det_edge ),
    .B(\inputs.octave_fsm.octave_key_up ),
    .X(_1210_));
 sky130_fd_sc_hd__or2b_1 _1630_ (.A(\inputs.octave_fsm.octave_key_up ),
    .B_N(\inputs.down.det_edge ),
    .X(_1211_));
 sky130_fd_sc_hd__or2b_1 _1631_ (.A(_1210_),
    .B_N(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(_1208_),
    .A2(_1209_),
    .B1(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__nor2b_2 _1633_ (.A(\inputs.octave_fsm.state[2] ),
    .B_N(\inputs.octave_fsm.state[0] ),
    .Y(_1214_));
 sky130_fd_sc_hd__inv_2 _1634_ (.A(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(\inputs.octave_fsm.state[1] ),
    .B(_1210_),
    .Y(_1216_));
 sky130_fd_sc_hd__o32a_1 _1636_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .A3(_1216_),
    .B1(_1208_),
    .B2(_1210_),
    .X(_1217_));
 sky130_fd_sc_hd__o31a_1 _1637_ (.A1(\inputs.octave_fsm.state[1] ),
    .A2(_1212_),
    .A3(_1215_),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__xnor2_1 _1638_ (.A(_1213_),
    .B(_1218_),
    .Y(_0000_));
 sky130_fd_sc_hd__a21o_1 _1639_ (.A1(\inputs.octave_fsm.state[1] ),
    .A2(\inputs.octave_fsm.state[0] ),
    .B1(\inputs.octave_fsm.state[2] ),
    .X(_1219_));
 sky130_fd_sc_hd__and3b_1 _1640_ (.A_N(\inputs.octave_fsm.state[2] ),
    .B(\inputs.octave_fsm.state[0] ),
    .C(\inputs.octave_fsm.state[1] ),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(_1205_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(_1219_),
    .A1(_1221_),
    .S(_1210_),
    .X(_1222_));
 sky130_fd_sc_hd__o22a_1 _1643_ (.A1(_1212_),
    .A2(_1208_),
    .B1(_1213_),
    .B2(_1222_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1644_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_1205_),
    .X(_1223_));
 sky130_fd_sc_hd__buf_2 _1645_ (.A(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _1646_ (.A1(_1211_),
    .A2(_1224_),
    .B1(_1220_),
    .B2(_1210_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _1647_ (.A(_0996_),
    .X(_1225_));
 sky130_fd_sc_hd__nand2_1 _1648_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.q[26] ),
    .Y(_1226_));
 sky130_fd_sc_hd__or2_1 _1649_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.q[26] ),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_4 _1650_ (.A(_0915_),
    .X(_1228_));
 sky130_fd_sc_hd__a32o_1 _1651_ (.A1(_1225_),
    .A2(_1226_),
    .A3(_1227_),
    .B1(_1228_),
    .B2(net173),
    .X(_0003_));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(\outputs.div.a[25] ),
    .Y(_1229_));
 sky130_fd_sc_hd__a21o_1 _1653_ (.A1(\outputs.div.m[0] ),
    .A2(_1229_),
    .B1(\outputs.div.m[1] ),
    .X(_1230_));
 sky130_fd_sc_hd__nand3_1 _1654_ (.A(\outputs.div.m[0] ),
    .B(\outputs.div.m[1] ),
    .C(_1229_),
    .Y(_1231_));
 sky130_fd_sc_hd__and3_1 _1655_ (.A(\outputs.div.a[0] ),
    .B(_1230_),
    .C(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__a21oi_1 _1656_ (.A1(_1230_),
    .A2(_1231_),
    .B1(\outputs.div.a[0] ),
    .Y(_1233_));
 sky130_fd_sc_hd__or2_1 _1657_ (.A(_1232_),
    .B(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__xor2_1 _1658_ (.A(_1226_),
    .B(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a22o_1 _1659_ (.A1(net210),
    .A2(_0916_),
    .B1(\outputs.div.next_div ),
    .B2(_1235_),
    .X(_0004_));
 sky130_fd_sc_hd__o21ba_1 _1660_ (.A1(_1226_),
    .A2(_1233_),
    .B1_N(_1232_),
    .X(_1236_));
 sky130_fd_sc_hd__inv_2 _1661_ (.A(\outputs.div.a[1] ),
    .Y(_1237_));
 sky130_fd_sc_hd__o21ba_1 _1662_ (.A1(\outputs.div.m[0] ),
    .A2(\outputs.div.m[1] ),
    .B1_N(\outputs.div.a[25] ),
    .X(_1238_));
 sky130_fd_sc_hd__xnor2_1 _1663_ (.A(\outputs.div.m[2] ),
    .B(_1238_),
    .Y(_0191_));
 sky130_fd_sc_hd__or2_1 _1664_ (.A(_1237_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _1665_ (.A(_1237_),
    .B(_0191_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _1666_ (.A(_0192_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _1667_ (.A(_1236_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__or2_1 _1668_ (.A(_1236_),
    .B(_0194_),
    .X(_0196_));
 sky130_fd_sc_hd__a32o_1 _1669_ (.A1(_1225_),
    .A2(_0195_),
    .A3(_0196_),
    .B1(_1228_),
    .B2(net231),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _1670_ (.A(_0192_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__a21o_1 _1671_ (.A1(\outputs.div.m[2] ),
    .A2(_1229_),
    .B1(_1238_),
    .X(_0198_));
 sky130_fd_sc_hd__xor2_1 _1672_ (.A(\outputs.div.m[3] ),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_1 _1673_ (.A(\outputs.div.a[2] ),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__nor2_1 _1674_ (.A(\outputs.div.a[2] ),
    .B(_0199_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor2_1 _1675_ (.A(_0200_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(_0197_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__o21a_1 _1677_ (.A1(_0197_),
    .A2(_0202_),
    .B1(_0996_),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _1678_ (.A1(net278),
    .A2(_0916_),
    .B1(_0203_),
    .B2(_0204_),
    .X(_0006_));
 sky130_fd_sc_hd__clkbuf_4 _1679_ (.A(_0996_),
    .X(_0205_));
 sky130_fd_sc_hd__nand2_1 _1680_ (.A(\outputs.div.a[2] ),
    .B(_0199_),
    .Y(_0206_));
 sky130_fd_sc_hd__o211a_1 _1681_ (.A1(_1236_),
    .A2(_0194_),
    .B1(_0206_),
    .C1(_0192_),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_1 _1682_ (.A(_0201_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__or4_2 _1683_ (.A(\outputs.div.m[3] ),
    .B(\outputs.div.m[2] ),
    .C(\outputs.div.m[0] ),
    .D(\outputs.div.m[1] ),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(_1229_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_2 _1685_ (.A(\outputs.div.m[4] ),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_1 _1686_ (.A(\outputs.div.a[3] ),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2_1 _1687_ (.A(_0208_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__or2_1 _1688_ (.A(_0208_),
    .B(_0212_),
    .X(_0214_));
 sky130_fd_sc_hd__a32o_1 _1689_ (.A1(_0205_),
    .A2(_0213_),
    .A3(_0214_),
    .B1(_1228_),
    .B2(net182),
    .X(_0007_));
 sky130_fd_sc_hd__inv_2 _1690_ (.A(\outputs.div.a[3] ),
    .Y(_0215_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_0215_),
    .B(_0211_),
    .X(_0216_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(\outputs.div.a[4] ),
    .Y(_0217_));
 sky130_fd_sc_hd__o21a_1 _1693_ (.A1(\outputs.div.m[4] ),
    .A2(_0209_),
    .B1(_1229_),
    .X(_0218_));
 sky130_fd_sc_hd__xnor2_2 _1694_ (.A(\outputs.div.m[5] ),
    .B(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__xnor2_1 _1695_ (.A(_0217_),
    .B(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__a21o_1 _1696_ (.A1(_0216_),
    .A2(_0213_),
    .B1(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__nand3_1 _1697_ (.A(_0216_),
    .B(_0213_),
    .C(_0220_),
    .Y(_0222_));
 sky130_fd_sc_hd__a32o_1 _1698_ (.A1(_0205_),
    .A2(_0221_),
    .A3(_0222_),
    .B1(_1228_),
    .B2(net191),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _1699_ (.A(\outputs.div.a[5] ),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _1700_ (.A(\outputs.div.m[5] ),
    .B(\outputs.div.m[4] ),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_1 _1701_ (.A1(_0209_),
    .A2(_0224_),
    .B1(_1229_),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_1 _1702_ (.A(\outputs.div.m[6] ),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__or2_1 _1703_ (.A(_0223_),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_1 _1704_ (.A(_0223_),
    .B(_0226_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(_0215_),
    .B(_0211_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _1707_ (.A(_0216_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__o22a_1 _1708_ (.A1(_0215_),
    .A2(_0211_),
    .B1(_0219_),
    .B2(_0217_),
    .X(_0232_));
 sky130_fd_sc_hd__a21o_1 _1709_ (.A1(_0217_),
    .A2(_0219_),
    .B1(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__o41a_1 _1710_ (.A1(_0201_),
    .A2(_0207_),
    .A3(_0231_),
    .A4(_0220_),
    .B1(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _1711_ (.A(_0229_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_0229_),
    .B(_0234_),
    .Y(_0236_));
 sky130_fd_sc_hd__a32o_1 _1713_ (.A1(_0205_),
    .A2(_0235_),
    .A3(_0236_),
    .B1(_1228_),
    .B2(net190),
    .X(_0009_));
 sky130_fd_sc_hd__inv_2 _1714_ (.A(\outputs.div.a[6] ),
    .Y(_0237_));
 sky130_fd_sc_hd__o31a_1 _1715_ (.A1(\outputs.div.m[6] ),
    .A2(_0209_),
    .A3(_0224_),
    .B1(_1229_),
    .X(_0238_));
 sky130_fd_sc_hd__xnor2_1 _1716_ (.A(\outputs.div.m[7] ),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _1717_ (.A(_0237_),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(_0237_),
    .B(_0239_),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _1719_ (.A(_0240_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__o21a_1 _1720_ (.A1(_0229_),
    .A2(_0234_),
    .B1(_0227_),
    .X(_0243_));
 sky130_fd_sc_hd__xor2_1 _1721_ (.A(_0242_),
    .B(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _1722_ (.A1(net211),
    .A2(_0916_),
    .B1(\outputs.div.next_div ),
    .B2(_0244_),
    .X(_0010_));
 sky130_fd_sc_hd__o21a_1 _1723_ (.A1(_0237_),
    .A2(_0239_),
    .B1(_0227_),
    .X(_0245_));
 sky130_fd_sc_hd__o32a_2 _1724_ (.A1(_0229_),
    .A2(_0234_),
    .A3(_0242_),
    .B1(_0245_),
    .B2(_0241_),
    .X(_0246_));
 sky130_fd_sc_hd__inv_2 _1725_ (.A(\outputs.div.a[7] ),
    .Y(_0247_));
 sky130_fd_sc_hd__buf_2 _1726_ (.A(_1229_),
    .X(_0248_));
 sky130_fd_sc_hd__or4_2 _1727_ (.A(\outputs.div.m[7] ),
    .B(\outputs.div.m[6] ),
    .C(_0209_),
    .D(_0224_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _1728_ (.A(_0248_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__xor2_1 _1729_ (.A(\outputs.div.m[8] ),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_1 _1730_ (.A(_0247_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__and2_1 _1731_ (.A(_0247_),
    .B(_0251_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_2 _1732_ (.A(_0252_),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_1 _1733_ (.A(_0246_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21bo_1 _1734_ (.A1(_0246_),
    .A2(_0254_),
    .B1_N(_0996_),
    .X(_0256_));
 sky130_fd_sc_hd__a2bb2o_1 _1735_ (.A1_N(_0255_),
    .A2_N(_0256_),
    .B1(net192),
    .B2(_0916_),
    .X(_0011_));
 sky130_fd_sc_hd__o21a_1 _1736_ (.A1(\outputs.div.m[8] ),
    .A2(_0249_),
    .B1(_1229_),
    .X(_0257_));
 sky130_fd_sc_hd__xor2_1 _1737_ (.A(\outputs.div.m[9] ),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__and2_1 _1738_ (.A(\outputs.div.a[8] ),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _1739_ (.A(\outputs.div.a[8] ),
    .B(_0258_),
    .X(_0260_));
 sky130_fd_sc_hd__and2b_1 _1740_ (.A_N(_0259_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__o21ai_1 _1741_ (.A1(_0252_),
    .A2(_0255_),
    .B1(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__o31a_1 _1742_ (.A1(_0252_),
    .A2(_0255_),
    .A3(_0261_),
    .B1(_0996_),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _1743_ (.A1(net268),
    .A2(_0916_),
    .B1(_0262_),
    .B2(_0263_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _1744_ (.A(\outputs.div.m[9] ),
    .B(\outputs.div.m[8] ),
    .X(_0264_));
 sky130_fd_sc_hd__o21a_1 _1745_ (.A1(_0249_),
    .A2(_0264_),
    .B1(_0248_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_2 _1746_ (.A(\outputs.div.m[10] ),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__xnor2_2 _1747_ (.A(\outputs.div.a[9] ),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _1748_ (.A(_0261_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_1 _1749_ (.A1(_0252_),
    .A2(_0259_),
    .B1(_0260_),
    .Y(_0269_));
 sky130_fd_sc_hd__o31ai_4 _1750_ (.A1(_0246_),
    .A2(_0254_),
    .A3(_0268_),
    .B1(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _1751_ (.A(_0267_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__or2_1 _1752_ (.A(_0267_),
    .B(_0270_),
    .X(_0272_));
 sky130_fd_sc_hd__a32o_1 _1753_ (.A1(_0205_),
    .A2(_0271_),
    .A3(_0272_),
    .B1(_1228_),
    .B2(net180),
    .X(_0013_));
 sky130_fd_sc_hd__o31a_1 _1754_ (.A1(\outputs.div.m[10] ),
    .A2(_0249_),
    .A3(_0264_),
    .B1(_0248_),
    .X(_0273_));
 sky130_fd_sc_hd__xnor2_1 _1755_ (.A(\outputs.div.m[11] ),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _1756_ (.A(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_2 _1757_ (.A(\outputs.div.a[10] ),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(\outputs.div.a[10] ),
    .B(_0275_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _1759_ (.A(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _1760_ (.A(_0276_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _1761_ (.A(\outputs.div.a[9] ),
    .Y(_0280_));
 sky130_fd_sc_hd__or2_1 _1762_ (.A(_0280_),
    .B(_0266_),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_0281_),
    .B(_0271_),
    .Y(_0282_));
 sky130_fd_sc_hd__xnor2_1 _1764_ (.A(_0279_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__a22o_1 _1765_ (.A1(net225),
    .A2(_0916_),
    .B1(\outputs.div.next_div ),
    .B2(_0283_),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _1766_ (.A(\outputs.div.a[11] ),
    .Y(_0284_));
 sky130_fd_sc_hd__or4_2 _1767_ (.A(\outputs.div.m[11] ),
    .B(\outputs.div.m[10] ),
    .C(_0249_),
    .D(_0264_),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_1 _1768_ (.A(_0248_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__xor2_1 _1769_ (.A(\outputs.div.m[12] ),
    .B(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _1770_ (.A(_0284_),
    .B(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(_0284_),
    .B(_0287_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _1772_ (.A(_0288_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21oi_1 _1773_ (.A1(_0281_),
    .A2(_0276_),
    .B1(_0277_),
    .Y(_0291_));
 sky130_fd_sc_hd__a41oi_4 _1774_ (.A1(_0267_),
    .A2(_0270_),
    .A3(_0276_),
    .A4(_0278_),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__or2_1 _1775_ (.A(_0290_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(_0290_),
    .B(_0292_),
    .Y(_0294_));
 sky130_fd_sc_hd__a32o_1 _1777_ (.A1(_0205_),
    .A2(_0293_),
    .A3(_0294_),
    .B1(_1228_),
    .B2(net181),
    .X(_0015_));
 sky130_fd_sc_hd__inv_2 _1778_ (.A(\outputs.div.a[12] ),
    .Y(_0295_));
 sky130_fd_sc_hd__o21a_1 _1779_ (.A1(\outputs.div.m[12] ),
    .A2(_0285_),
    .B1(_0248_),
    .X(_0296_));
 sky130_fd_sc_hd__xnor2_1 _1780_ (.A(\outputs.div.m[13] ),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _1781_ (.A(_0295_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__and2_1 _1782_ (.A(_0295_),
    .B(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _1783_ (.A(_0298_),
    .B(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__o21ai_1 _1784_ (.A1(_0290_),
    .A2(_0292_),
    .B1(_0288_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_1 _1785_ (.A(_0300_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__a22o_1 _1786_ (.A1(net224),
    .A2(_0916_),
    .B1(\outputs.div.next_div ),
    .B2(_0302_),
    .X(_0016_));
 sky130_fd_sc_hd__inv_2 _1787_ (.A(\outputs.div.a[13] ),
    .Y(_0303_));
 sky130_fd_sc_hd__o31a_1 _1788_ (.A1(\outputs.div.m[13] ),
    .A2(\outputs.div.m[12] ),
    .A3(_0285_),
    .B1(_0248_),
    .X(_0304_));
 sky130_fd_sc_hd__xnor2_1 _1789_ (.A(\outputs.div.m[14] ),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__or2_1 _1790_ (.A(_0303_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(_0303_),
    .B(_0305_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2_1 _1792_ (.A(_0306_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _1793_ (.A(_0298_),
    .Y(_0309_));
 sky130_fd_sc_hd__a21o_1 _1794_ (.A1(_0288_),
    .A2(_0309_),
    .B1(_0299_),
    .X(_0310_));
 sky130_fd_sc_hd__o31a_1 _1795_ (.A1(_0290_),
    .A2(_0292_),
    .A3(_0300_),
    .B1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _1796_ (.A(_0308_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(_0308_),
    .B(_0311_),
    .Y(_0313_));
 sky130_fd_sc_hd__a32o_1 _1798_ (.A1(_0205_),
    .A2(_0312_),
    .A3(_0313_),
    .B1(_1228_),
    .B2(net166),
    .X(_0017_));
 sky130_fd_sc_hd__or4_2 _1799_ (.A(\outputs.div.m[14] ),
    .B(\outputs.div.m[13] ),
    .C(\outputs.div.m[12] ),
    .D(_0285_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _1800_ (.A(_0248_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__xor2_1 _1801_ (.A(\outputs.div.m[15] ),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__inv_2 _1802_ (.A(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(\outputs.div.a[14] ),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__or2_1 _1804_ (.A(\outputs.div.a[14] ),
    .B(_0317_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(_0318_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_1 _1806_ (.A1(_0308_),
    .A2(_0311_),
    .B1(_0306_),
    .Y(_0321_));
 sky130_fd_sc_hd__xnor2_1 _1807_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__a22o_1 _1808_ (.A1(net228),
    .A2(_0916_),
    .B1(\outputs.div.next_div ),
    .B2(_0322_),
    .X(_0018_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(\outputs.div.a[15] ),
    .Y(_0323_));
 sky130_fd_sc_hd__o21a_1 _1810_ (.A1(\outputs.div.m[15] ),
    .A2(_0314_),
    .B1(_0248_),
    .X(_0324_));
 sky130_fd_sc_hd__xnor2_1 _1811_ (.A(\outputs.div.m[16] ),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__or2_1 _1812_ (.A(_0323_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _1813_ (.A(_0323_),
    .B(_0325_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _1814_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__a21bo_1 _1815_ (.A1(_0306_),
    .A2(_0318_),
    .B1_N(_0319_),
    .X(_0329_));
 sky130_fd_sc_hd__o31a_2 _1816_ (.A1(_0308_),
    .A2(_0311_),
    .A3(_0320_),
    .B1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _1817_ (.A(_0328_),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _1818_ (.A(_0328_),
    .B(_0330_),
    .Y(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _1819_ (.A(_0914_),
    .X(_0333_));
 sky130_fd_sc_hd__a32o_1 _1820_ (.A1(_0205_),
    .A2(_0331_),
    .A3(_0332_),
    .B1(_0333_),
    .B2(net172),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _1821_ (.A(_0915_),
    .X(_0334_));
 sky130_fd_sc_hd__inv_2 _1822_ (.A(\outputs.div.a[16] ),
    .Y(_0335_));
 sky130_fd_sc_hd__or3_1 _1823_ (.A(\outputs.div.m[16] ),
    .B(\outputs.div.m[15] ),
    .C(_0314_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _1824_ (.A(_0248_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__xnor2_2 _1825_ (.A(\outputs.div.m[17] ),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_1 _1826_ (.A(_0335_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_1 _1827_ (.A1(_0328_),
    .A2(_0330_),
    .B1(_0326_),
    .Y(_0340_));
 sky130_fd_sc_hd__xnor2_1 _1828_ (.A(_0339_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__a22o_1 _1829_ (.A1(net229),
    .A2(_0334_),
    .B1(\outputs.div.next_div ),
    .B2(_0341_),
    .X(_0020_));
 sky130_fd_sc_hd__o21a_2 _1830_ (.A1(\outputs.div.m[17] ),
    .A2(_0336_),
    .B1(_0248_),
    .X(_0342_));
 sky130_fd_sc_hd__nand2_1 _1831_ (.A(\outputs.div.a[17] ),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__or2_1 _1832_ (.A(\outputs.div.a[17] ),
    .B(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__nand2_1 _1833_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__or2_1 _1834_ (.A(_0328_),
    .B(_0339_),
    .X(_0346_));
 sky130_fd_sc_hd__o21a_1 _1835_ (.A1(_0335_),
    .A2(_0338_),
    .B1(_0326_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_1 _1836_ (.A1(_0335_),
    .A2(_0338_),
    .B1(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__o21ba_1 _1837_ (.A1(_0330_),
    .A2(_0346_),
    .B1_N(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__xor2_1 _1838_ (.A(_0345_),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _1839_ (.A1(net266),
    .A2(_0334_),
    .B1(\outputs.div.next_div ),
    .B2(_0350_),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _1840_ (.A(\outputs.div.a[18] ),
    .B(_0342_),
    .Y(_0351_));
 sky130_fd_sc_hd__o21ai_1 _1841_ (.A1(_0345_),
    .A2(_0349_),
    .B1(_0343_),
    .Y(_0352_));
 sky130_fd_sc_hd__xnor2_1 _1842_ (.A(_0351_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__a22o_1 _1843_ (.A1(net251),
    .A2(_0334_),
    .B1(\outputs.div.next_div ),
    .B2(_0353_),
    .X(_0022_));
 sky130_fd_sc_hd__or3_1 _1844_ (.A(_0345_),
    .B(_0346_),
    .C(_0351_),
    .X(_0354_));
 sky130_fd_sc_hd__buf_2 _1845_ (.A(_0342_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_1 _1846_ (.A(_0345_),
    .B(_0351_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(_0343_),
    .Y(_0357_));
 sky130_fd_sc_hd__a221o_1 _1848_ (.A1(\outputs.div.a[18] ),
    .A2(_0355_),
    .B1(_0348_),
    .B2(_0356_),
    .C1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__o21ba_1 _1849_ (.A1(_0330_),
    .A2(_0354_),
    .B1_N(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_2 _1850_ (.A(\outputs.div.a[19] ),
    .B(_0342_),
    .Y(_0360_));
 sky130_fd_sc_hd__or2_1 _1851_ (.A(\outputs.div.a[19] ),
    .B(_0342_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _1852_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__or2_1 _1853_ (.A(_0359_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _1854_ (.A(_0359_),
    .B(_0362_),
    .Y(_0364_));
 sky130_fd_sc_hd__a32o_1 _1855_ (.A1(_0205_),
    .A2(_0363_),
    .A3(_0364_),
    .B1(_0333_),
    .B2(net236),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _1856_ (.A(\outputs.div.a[20] ),
    .B(_0355_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _1857_ (.A(\outputs.div.a[20] ),
    .B(_0342_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _1858_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__a21o_1 _1859_ (.A1(_0360_),
    .A2(_0363_),
    .B1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__nand3_1 _1860_ (.A(_0360_),
    .B(_0363_),
    .C(_0367_),
    .Y(_0369_));
 sky130_fd_sc_hd__a32o_1 _1861_ (.A1(_0205_),
    .A2(_0368_),
    .A3(_0369_),
    .B1(_0333_),
    .B2(net238),
    .X(_0024_));
 sky130_fd_sc_hd__or2_1 _1862_ (.A(_0362_),
    .B(_0367_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _1863_ (.A(_0359_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _1864_ (.A(\outputs.div.a[21] ),
    .B(_0355_),
    .Y(_0372_));
 sky130_fd_sc_hd__or2_1 _1865_ (.A(\outputs.div.a[21] ),
    .B(_0355_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_1 _1866_ (.A(_0372_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__a31o_1 _1867_ (.A1(_0360_),
    .A2(_0365_),
    .A3(_0371_),
    .B1(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__nand4_1 _1868_ (.A(_0360_),
    .B(_0365_),
    .C(_0374_),
    .D(_0371_),
    .Y(_0376_));
 sky130_fd_sc_hd__a32o_1 _1869_ (.A1(_0205_),
    .A2(_0375_),
    .A3(_0376_),
    .B1(_0333_),
    .B2(net243),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_4 _1870_ (.A(_0995_),
    .X(_0377_));
 sky130_fd_sc_hd__xnor2_1 _1871_ (.A(\outputs.div.a[22] ),
    .B(_0355_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _1872_ (.A1(_0372_),
    .A2(_0375_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__nand3_1 _1873_ (.A(_0372_),
    .B(_0375_),
    .C(_0378_),
    .Y(_0380_));
 sky130_fd_sc_hd__a32o_1 _1874_ (.A1(_0377_),
    .A2(_0379_),
    .A3(_0380_),
    .B1(_0333_),
    .B2(net188),
    .X(_0026_));
 sky130_fd_sc_hd__or4_1 _1875_ (.A(_0359_),
    .B(_0374_),
    .C(_0370_),
    .D(_0378_),
    .X(_0381_));
 sky130_fd_sc_hd__o41ai_1 _1876_ (.A1(\outputs.div.a[22] ),
    .A2(\outputs.div.a[21] ),
    .A3(\outputs.div.a[20] ),
    .A4(\outputs.div.a[19] ),
    .B1(_0355_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _1877_ (.A(\outputs.div.a[23] ),
    .B(_0355_),
    .Y(_0383_));
 sky130_fd_sc_hd__or2_1 _1878_ (.A(\outputs.div.a[23] ),
    .B(_0355_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _1879_ (.A(_0383_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _1880_ (.A(_0381_),
    .B(_0382_),
    .C(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a21o_1 _1881_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0385_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _1882_ (.A(_0996_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__a2bb2o_1 _1883_ (.A1_N(_0386_),
    .A2_N(_0388_),
    .B1(net215),
    .B2(_0916_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(\outputs.div.a[24] ),
    .B(_0355_),
    .Y(_0389_));
 sky130_fd_sc_hd__or2_1 _1885_ (.A(\outputs.div.a[24] ),
    .B(_0355_),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _1886_ (.A(_0389_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a21o_1 _1887_ (.A1(_0383_),
    .A2(_0387_),
    .B1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__nand3_1 _1888_ (.A(_0383_),
    .B(_0387_),
    .C(_0391_),
    .Y(_0393_));
 sky130_fd_sc_hd__a32o_1 _1889_ (.A1(_0377_),
    .A2(_0392_),
    .A3(_0393_),
    .B1(_0333_),
    .B2(net302),
    .X(_0028_));
 sky130_fd_sc_hd__o311a_1 _1890_ (.A1(\outputs.div.m[17] ),
    .A2(\outputs.div.a[25] ),
    .A3(_0336_),
    .B1(_0383_),
    .C1(_0389_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _1891_ (.A1(_0387_),
    .A2(_0391_),
    .B1(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a22o_1 _1892_ (.A1(net257),
    .A2(_0334_),
    .B1(\outputs.div.next_div ),
    .B2(_0395_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _1893_ (.A1(net244),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net257),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _1894_ (.A1(net233),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net244),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _1895_ (.A1(\outputs.div.q[3] ),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net233),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _1896_ (.A1(\outputs.div.q[4] ),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net252),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _1897_ (.A1(net258),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net260),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _1898_ (.A1(\outputs.div.q[6] ),
    .A2(_0334_),
    .B1(_1225_),
    .B2(net258),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _1899_ (.A1(\outputs.div.q[7] ),
    .A2(_1228_),
    .B1(_1225_),
    .B2(net262),
    .X(_0036_));
 sky130_fd_sc_hd__buf_4 _1900_ (.A(_0994_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _1901_ (.A(\outputs.div.oscillator_out[0] ),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _1902_ (.A1(net195),
    .A2(_0333_),
    .B1(_0377_),
    .B2(net271),
    .C1(_0397_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _1903_ (.A(_0994_),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _1904_ (.A(\outputs.div.oscillator_out[1] ),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__a221o_1 _1905_ (.A1(net189),
    .A2(_0333_),
    .B1(_0377_),
    .B2(net195),
    .C1(_0399_),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_4 _1906_ (.A(_0914_),
    .X(_0400_));
 sky130_fd_sc_hd__and2_1 _1907_ (.A(net315),
    .B(_0398_),
    .X(_0401_));
 sky130_fd_sc_hd__a221o_1 _1908_ (.A1(net183),
    .A2(_0400_),
    .B1(_0377_),
    .B2(net189),
    .C1(_0401_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _1909_ (.A(\outputs.div.oscillator_out[3] ),
    .B(_0398_),
    .X(_0402_));
 sky130_fd_sc_hd__a221o_1 _1910_ (.A1(net98),
    .A2(_0400_),
    .B1(_0377_),
    .B2(net183),
    .C1(_0402_),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _1911_ (.A(\outputs.div.oscillator_out[4] ),
    .B(_0398_),
    .X(_0403_));
 sky130_fd_sc_hd__a221o_1 _1912_ (.A1(\outputs.div.q[12] ),
    .A2(_0400_),
    .B1(_0377_),
    .B2(net98),
    .C1(_0403_),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _1913_ (.A(\outputs.div.oscillator_out[5] ),
    .B(_0398_),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _1914_ (.A1(net167),
    .A2(_0400_),
    .B1(_0377_),
    .B2(net208),
    .C1(_0404_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _1915_ (.A(_0995_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _1916_ (.A(\outputs.div.oscillator_out[6] ),
    .B(_0398_),
    .X(_0406_));
 sky130_fd_sc_hd__a221o_1 _1917_ (.A1(\outputs.div.q[14] ),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net167),
    .C1(_0406_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _1918_ (.A(\outputs.div.oscillator_out[7] ),
    .B(_0398_),
    .X(_0407_));
 sky130_fd_sc_hd__a221o_1 _1919_ (.A1(net150),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net196),
    .C1(_0407_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _1920_ (.A(\outputs.div.oscillator_out[8] ),
    .B(_0398_),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _1921_ (.A1(net137),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net150),
    .C1(_0408_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _1922_ (.A(\outputs.div.oscillator_out[9] ),
    .B(_0398_),
    .X(_0409_));
 sky130_fd_sc_hd__a221o_1 _1923_ (.A1(\outputs.div.q[17] ),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net137),
    .C1(_0409_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _1924_ (.A(\outputs.div.oscillator_out[10] ),
    .B(_0398_),
    .X(_0410_));
 sky130_fd_sc_hd__a221o_1 _1925_ (.A1(\outputs.div.q[18] ),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net143),
    .C1(_0410_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _1926_ (.A(_0994_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _1927_ (.A(\outputs.div.oscillator_out[11] ),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__a221o_1 _1928_ (.A1(net187),
    .A2(_0400_),
    .B1(_0405_),
    .B2(net193),
    .C1(_0412_),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _1929_ (.A(net314),
    .B(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__a221o_1 _1930_ (.A1(net141),
    .A2(_0915_),
    .B1(_0405_),
    .B2(net187),
    .C1(_0413_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _1931_ (.A(\outputs.div.oscillator_out[13] ),
    .B(_0411_),
    .X(_0414_));
 sky130_fd_sc_hd__a221o_1 _1932_ (.A1(\outputs.div.q[21] ),
    .A2(_0915_),
    .B1(_0405_),
    .B2(net141),
    .C1(_0414_),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _1933_ (.A(\outputs.div.oscillator_out[14] ),
    .B(_0411_),
    .X(_0415_));
 sky130_fd_sc_hd__a221o_1 _1934_ (.A1(\outputs.div.q[22] ),
    .A2(_0915_),
    .B1(_0405_),
    .B2(net178),
    .C1(_0415_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _1935_ (.A(net313),
    .B(_0411_),
    .X(_0416_));
 sky130_fd_sc_hd__a221o_1 _1936_ (.A1(net96),
    .A2(_0915_),
    .B1(_0405_),
    .B2(net201),
    .C1(_0416_),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _1937_ (.A(\outputs.div.oscillator_out[16] ),
    .B(_0411_),
    .X(_0417_));
 sky130_fd_sc_hd__a221o_1 _1938_ (.A1(\outputs.div.q[24] ),
    .A2(_0915_),
    .B1(_0996_),
    .B2(net96),
    .C1(_0417_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _1939_ (.A(\outputs.div.oscillator_out[17] ),
    .B(_0411_),
    .X(_0418_));
 sky130_fd_sc_hd__a221o_1 _1940_ (.A1(\outputs.div.q[25] ),
    .A2(_0915_),
    .B1(_0996_),
    .B2(net204),
    .C1(_0418_),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _1941_ (.A1(net216),
    .A2(_1228_),
    .B1(_1225_),
    .B2(\outputs.div.q[25] ),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(_0996_),
    .A1(_0915_),
    .S(\outputs.div.count[0] ),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1943_ (.A(_0419_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _1944_ (.A(\outputs.div.count[1] ),
    .B(\outputs.div.count[0] ),
    .Y(_0420_));
 sky130_fd_sc_hd__or2_1 _1945_ (.A(\outputs.div.count[1] ),
    .B(\outputs.div.count[0] ),
    .X(_0421_));
 sky130_fd_sc_hd__a32o_1 _1946_ (.A1(_0420_),
    .A2(_0377_),
    .A3(_0421_),
    .B1(_0333_),
    .B2(net246),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _1947_ (.A(\outputs.div.count[2] ),
    .B(\outputs.div.count[1] ),
    .C(\outputs.div.count[0] ),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _1948_ (.A(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a32o_1 _1949_ (.A1(_0911_),
    .A2(_0377_),
    .A3(_0423_),
    .B1(_0333_),
    .B2(net176),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _1950_ (.A(\outputs.div.count[3] ),
    .Y(_0424_));
 sky130_fd_sc_hd__or3_1 _1951_ (.A(_0424_),
    .B(_0913_),
    .C(_0423_),
    .X(_0425_));
 sky130_fd_sc_hd__a21o_1 _1952_ (.A1(\outputs.div.start ),
    .A2(_0422_),
    .B1(\outputs.div.count[3] ),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _1953_ (.A(_0910_),
    .B(_0425_),
    .C(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _1954_ (.A(_0427_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _1955_ (.A(net235),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_1 _1956_ (.A1(_0428_),
    .A2(_0425_),
    .B1(_1001_),
    .Y(_0060_));
 sky130_fd_sc_hd__mux2_1 _1957_ (.A0(\outputs.scaled_buffer[0] ),
    .A1(net164),
    .S(_1001_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1958_ (.A(_0429_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1959_ (.A0(\outputs.scaled_buffer[1] ),
    .A1(net154),
    .S(_1001_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1960_ (.A(_0430_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1961_ (.A0(\outputs.scaled_buffer[2] ),
    .A1(net160),
    .S(_1001_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1962_ (.A(_0431_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(\outputs.scaled_buffer[3] ),
    .A1(net170),
    .S(_1001_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1964_ (.A(_0432_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1965_ (.A0(\outputs.scaled_buffer[4] ),
    .A1(net174),
    .S(_1001_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _1966_ (.A(_0433_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1967_ (.A0(\outputs.scaled_buffer[5] ),
    .A1(net162),
    .S(_1001_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1968_ (.A(_0434_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(\outputs.scaled_buffer[6] ),
    .A1(\outputs.div.q_out[6] ),
    .S(_1001_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1970_ (.A(_0435_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_4 _1971_ (.A(_0411_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _1972_ (.A0(net308),
    .A1(net219),
    .S(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1973_ (.A(_0437_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _1974_ (.A(\outputs.div.div ),
    .B(_0910_),
    .C(_0913_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_4 _1975_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or3b_1 _1976_ (.A(\outputs.div.q[7] ),
    .B(\outputs.div.q[6] ),
    .C_N(\outputs.div.q[8] ),
    .X(_0440_));
 sky130_fd_sc_hd__or4_1 _1977_ (.A(\outputs.div.q[3] ),
    .B(\outputs.div.q[2] ),
    .C(\outputs.div.q[5] ),
    .D(\outputs.div.q[4] ),
    .X(_0441_));
 sky130_fd_sc_hd__or4_1 _1978_ (.A(\outputs.div.q[1] ),
    .B(\outputs.div.q[0] ),
    .C(_0440_),
    .D(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_2 _1979_ (.A(_0439_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__o22a_1 _1980_ (.A1(net164),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[0] ),
    .X(_0069_));
 sky130_fd_sc_hd__o22a_1 _1981_ (.A1(net154),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[1] ),
    .X(_0070_));
 sky130_fd_sc_hd__o22a_1 _1982_ (.A1(net160),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[2] ),
    .X(_0071_));
 sky130_fd_sc_hd__o22a_1 _1983_ (.A1(net170),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[3] ),
    .X(_0072_));
 sky130_fd_sc_hd__o22a_1 _1984_ (.A1(net174),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[4] ),
    .X(_0073_));
 sky130_fd_sc_hd__o22a_1 _1985_ (.A1(net162),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[5] ),
    .X(_0074_));
 sky130_fd_sc_hd__o22a_1 _1986_ (.A1(net198),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[6] ),
    .X(_0075_));
 sky130_fd_sc_hd__o22a_1 _1987_ (.A1(net219),
    .A2(_0439_),
    .B1(_0443_),
    .B2(\outputs.div.q[7] ),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1988_ (.A0(\outputs.div.m[0] ),
    .A1(net283),
    .S(_0436_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _1989_ (.A(_0444_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1990_ (.A0(\outputs.div.m[1] ),
    .A1(net280),
    .S(_0436_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _1991_ (.A(_0445_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(\outputs.div.m[2] ),
    .A1(net222),
    .S(_0436_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _1993_ (.A(_0446_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(\outputs.div.m[3] ),
    .A1(net240),
    .S(_0436_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _1995_ (.A(_0447_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1996_ (.A0(\outputs.div.m[4] ),
    .A1(net273),
    .S(_0436_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1997_ (.A(_0448_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1998_ (.A0(\outputs.div.m[5] ),
    .A1(net294),
    .S(_0436_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _1999_ (.A(_0449_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2000_ (.A0(\outputs.div.m[6] ),
    .A1(net159),
    .S(_0436_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _2001_ (.A(_0450_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(\outputs.div.m[7] ),
    .A1(net282),
    .S(_0436_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _2003_ (.A(_0451_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2004_ (.A0(\outputs.div.m[8] ),
    .A1(net292),
    .S(_0436_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _2005_ (.A(_0452_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_4 _2006_ (.A(_0411_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _2007_ (.A0(\outputs.div.m[9] ),
    .A1(net295),
    .S(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _2008_ (.A(_0454_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2009_ (.A0(\outputs.div.m[10] ),
    .A1(net285),
    .S(_0453_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _2010_ (.A(_0455_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2011_ (.A0(\outputs.div.m[11] ),
    .A1(net288),
    .S(_0453_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_0456_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2013_ (.A0(\outputs.div.m[12] ),
    .A1(net256),
    .S(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _2014_ (.A(_0457_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(\outputs.div.m[13] ),
    .A1(net286),
    .S(_0453_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _2016_ (.A(_0458_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(\outputs.div.m[14] ),
    .A1(net230),
    .S(_0453_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _2018_ (.A(_0459_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(\outputs.div.m[15] ),
    .A1(net239),
    .S(_0453_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _2020_ (.A(_0460_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(\outputs.div.m[16] ),
    .A1(net232),
    .S(_0453_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _2022_ (.A(_0461_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(\outputs.div.m[17] ),
    .A1(net122),
    .S(_0453_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _2024_ (.A(_0462_),
    .X(_0094_));
 sky130_fd_sc_hd__nand2_1 _2025_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(_1198_),
    .Y(_0463_));
 sky130_fd_sc_hd__clkbuf_4 _2026_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_4 _2027_ (.A(\inputs.frequency_lut.rng[2] ),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_4 _2028_ (.A(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _2029_ (.A(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _2030_ (.A(\inputs.frequency_lut.rng[0] ),
    .Y(_0468_));
 sky130_fd_sc_hd__or2_1 _2031_ (.A(_0468_),
    .B(\inputs.frequency_lut.rng[1] ),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _2032_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_2 _2033_ (.A(_0468_),
    .B(\inputs.frequency_lut.rng[1] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_2 _2034_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__clkbuf_4 _2035_ (.A(\inputs.frequency_lut.rng[1] ),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _2036_ (.A(_0473_),
    .B(_0465_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21a_1 _2037_ (.A1(_0467_),
    .A2(_0472_),
    .B1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _2038_ (.A(_0468_),
    .B(\inputs.frequency_lut.rng[1] ),
    .X(_0476_));
 sky130_fd_sc_hd__nor2_4 _2039_ (.A(_0465_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__and3_1 _2040_ (.A(\inputs.frequency_lut.rng[2] ),
    .B(_0469_),
    .C(_0471_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_2 _2041_ (.A(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_2 _2042_ (.A(_0477_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__buf_2 _2043_ (.A(\inputs.frequency_lut.rng[3] ),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_4 _2044_ (.A(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(_0475_),
    .A1(_0480_),
    .S(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(\inputs.frequency_lut.rng[3] ),
    .Y(_0484_));
 sky130_fd_sc_hd__clkbuf_4 _2047_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _2048_ (.A(\inputs.frequency_lut.rng[0] ),
    .X(_0486_));
 sky130_fd_sc_hd__a21o_1 _2049_ (.A1(_0486_),
    .A2(_0473_),
    .B1(_0466_),
    .X(_0487_));
 sky130_fd_sc_hd__nor2_2 _2050_ (.A(_0486_),
    .B(_0473_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_2 _2051_ (.A(_0467_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _2052_ (.A1(_0485_),
    .A2(_0487_),
    .B1(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__buf_2 _2053_ (.A(_0481_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_4 _2054_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _2055_ (.A(_0465_),
    .B(_0470_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_4 _2056_ (.A(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_1 _2057_ (.A(_0466_),
    .B(_0472_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2_1 _2058_ (.A(_0494_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_2 _2059_ (.A(_0467_),
    .B(_0470_),
    .Y(_0497_));
 sky130_fd_sc_hd__buf_2 _2060_ (.A(\inputs.frequency_lut.rng[3] ),
    .X(_0498_));
 sky130_fd_sc_hd__buf_2 _2061_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a21oi_1 _2062_ (.A1(_0494_),
    .A2(_0497_),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a21oi_1 _2063_ (.A1(_0492_),
    .A2(_0496_),
    .B1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_2 _2064_ (.A(_0473_),
    .B(_0466_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_1 _2065_ (.A(_0486_),
    .B(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21oi_1 _2066_ (.A1(_0492_),
    .A2(_0477_),
    .B1(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _2067_ (.A(\inputs.frequency_lut.rng[4] ),
    .Y(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _2068_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__inv_2 _2069_ (.A(\inputs.frequency_lut.rng[5] ),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_4 _2070_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__mux4_1 _2071_ (.A0(_0483_),
    .A1(_0490_),
    .A2(_0501_),
    .A3(_0504_),
    .S0(_0506_),
    .S1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__inv_2 _2072_ (.A(\inputs.key_encoder.sync_keys[2] ),
    .Y(_0510_));
 sky130_fd_sc_hd__a21oi_1 _2073_ (.A1(\inputs.key_encoder.sync_keys[1] ),
    .A2(_0510_),
    .B1(\inputs.key_encoder.sync_keys[3] ),
    .Y(_0511_));
 sky130_fd_sc_hd__o21ba_1 _2074_ (.A1(\inputs.key_encoder.sync_keys[4] ),
    .A2(_0511_),
    .B1_N(\inputs.key_encoder.sync_keys[5] ),
    .X(_0512_));
 sky130_fd_sc_hd__o21ba_1 _2075_ (.A1(\inputs.key_encoder.sync_keys[6] ),
    .A2(_0512_),
    .B1_N(\inputs.key_encoder.sync_keys[7] ),
    .X(_0513_));
 sky130_fd_sc_hd__o21ba_1 _2076_ (.A1(\inputs.key_encoder.sync_keys[8] ),
    .A2(_0513_),
    .B1_N(\inputs.key_encoder.sync_keys[9] ),
    .X(_0514_));
 sky130_fd_sc_hd__o21bai_4 _2077_ (.A1(\inputs.key_encoder.sync_keys[10] ),
    .A2(_0514_),
    .B1_N(\inputs.key_encoder.sync_keys[11] ),
    .Y(_0515_));
 sky130_fd_sc_hd__and2b_1 _2078_ (.A_N(\inputs.key_encoder.sync_keys[13] ),
    .B(_1198_),
    .X(_0516_));
 sky130_fd_sc_hd__o31a_1 _2079_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_1199_),
    .A3(_1202_),
    .B1(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__nor2_1 _2080_ (.A(\inputs.key_encoder.sync_keys[8] ),
    .B(\inputs.key_encoder.sync_keys[9] ),
    .Y(_0518_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(\inputs.key_encoder.sync_keys[4] ),
    .B(\inputs.key_encoder.sync_keys[5] ),
    .Y(_0519_));
 sky130_fd_sc_hd__a211o_1 _2082_ (.A1(_1200_),
    .A2(_0519_),
    .B1(\inputs.key_encoder.sync_keys[6] ),
    .C1(\inputs.key_encoder.sync_keys[7] ),
    .X(_0520_));
 sky130_fd_sc_hd__a211o_2 _2083_ (.A1(_0518_),
    .A2(_0520_),
    .B1(\inputs.key_encoder.sync_keys[11] ),
    .C1(\inputs.key_encoder.sync_keys[10] ),
    .X(_0521_));
 sky130_fd_sc_hd__nor2b_2 _2084_ (.A(\inputs.key_encoder.sync_keys[12] ),
    .B_N(_0516_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _2085_ (.A(_0521_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_1 _2086_ (.A(_0517_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__inv_2 _2087_ (.A(_1199_),
    .Y(_0525_));
 sky130_fd_sc_hd__and2_1 _2088_ (.A(_0525_),
    .B(_1202_),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_2 _2089_ (.A(_0526_),
    .B(_0522_),
    .Y(_0527_));
 sky130_fd_sc_hd__or2_2 _2090_ (.A(_0521_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or3_1 _2091_ (.A(_0525_),
    .B(_0515_),
    .C(_0523_),
    .X(_0529_));
 sky130_fd_sc_hd__nand2_1 _2092_ (.A(_0515_),
    .B(_0522_),
    .Y(_0530_));
 sky130_fd_sc_hd__or3_4 _2093_ (.A(_0517_),
    .B(_0521_),
    .C(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__o2111ai_2 _2094_ (.A1(_0515_),
    .A2(_0524_),
    .B1(_0528_),
    .C1(_0529_),
    .D1(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__and2_2 _2095_ (.A(\inputs.key_encoder.sync_keys[13] ),
    .B(_1198_),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _2096_ (.A(_0533_),
    .B(_0517_),
    .X(_0534_));
 sky130_fd_sc_hd__nand2_1 _2097_ (.A(_0530_),
    .B(_0523_),
    .Y(_0535_));
 sky130_fd_sc_hd__or2_1 _2098_ (.A(_0534_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__o211a_1 _2099_ (.A1(_0530_),
    .A2(_0528_),
    .B1(_0536_),
    .C1(_0531_),
    .X(_0537_));
 sky130_fd_sc_hd__or3b_1 _2100_ (.A(_0525_),
    .B(_0515_),
    .C_N(_0522_),
    .X(_0538_));
 sky130_fd_sc_hd__nand2b_2 _2101_ (.A_N(_0524_),
    .B(_0515_),
    .Y(_0539_));
 sky130_fd_sc_hd__and3_1 _2102_ (.A(_0537_),
    .B(_0538_),
    .C(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_4 _2103_ (.A(_1214_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(_0532_),
    .A1(_0540_),
    .S(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__o21a_1 _2105_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_0526_),
    .B1(_0516_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(_0543_),
    .B(_0528_),
    .Y(_0544_));
 sky130_fd_sc_hd__and2_1 _2107_ (.A(_0531_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or3_1 _2108_ (.A(_0525_),
    .B(_0521_),
    .C(_0530_),
    .X(_0546_));
 sky130_fd_sc_hd__and3_1 _2109_ (.A(_0529_),
    .B(_0544_),
    .C(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__inv_2 _2110_ (.A(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _2111_ (.A(_0521_),
    .B(_0538_),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _2112_ (.A(_0515_),
    .B(_0528_),
    .Y(_0550_));
 sky130_fd_sc_hd__or4b_1 _2113_ (.A(_0548_),
    .B(_0549_),
    .C(_0550_),
    .D_N(_0534_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(_0545_),
    .A1(_0551_),
    .S(_1215_),
    .X(_0552_));
 sky130_fd_sc_hd__a21o_1 _2115_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .B1(\inputs.octave_fsm.state[1] ),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_4 _2116_ (.A(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(_0542_),
    .A1(_0552_),
    .S(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__a21oi_4 _2118_ (.A1(\inputs.octave_fsm.state[0] ),
    .A2(\inputs.octave_fsm.state[2] ),
    .B1(\inputs.octave_fsm.state[1] ),
    .Y(_0556_));
 sky130_fd_sc_hd__or2b_1 _2119_ (.A(_0530_),
    .B_N(_0521_),
    .X(_0557_));
 sky130_fd_sc_hd__nor2_1 _2120_ (.A(_0534_),
    .B(_0535_),
    .Y(_0558_));
 sky130_fd_sc_hd__a311o_1 _2121_ (.A1(_0526_),
    .A2(_0522_),
    .A3(_0557_),
    .B1(_0549_),
    .C1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__nor2_1 _2122_ (.A(_0527_),
    .B(_0557_),
    .Y(_0560_));
 sky130_fd_sc_hd__or2_1 _2123_ (.A(_0515_),
    .B(_0528_),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_1 _2124_ (.A(_0524_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__or3_1 _2125_ (.A(_0558_),
    .B(_0560_),
    .C(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(_0559_),
    .A1(_0563_),
    .S(_1215_),
    .X(_0564_));
 sky130_fd_sc_hd__inv_2 _2127_ (.A(_0531_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _2128_ (.A(_0539_),
    .B(_0561_),
    .Y(_0566_));
 sky130_fd_sc_hd__a31o_1 _2129_ (.A1(_0526_),
    .A2(_0521_),
    .A3(_0522_),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__or3b_1 _2130_ (.A(_0565_),
    .B(_0567_),
    .C_N(_0546_),
    .X(_0568_));
 sky130_fd_sc_hd__a31oi_1 _2131_ (.A1(_0537_),
    .A2(_0539_),
    .A3(_0544_),
    .B1(_0541_),
    .Y(_0569_));
 sky130_fd_sc_hd__a211o_1 _2132_ (.A1(_0541_),
    .A2(_0568_),
    .B1(_0569_),
    .C1(_0554_),
    .X(_0570_));
 sky130_fd_sc_hd__o211a_1 _2133_ (.A1(_0556_),
    .A2(_0564_),
    .B1(_0570_),
    .C1(_1207_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_4 _2134_ (.A(_0533_),
    .X(_0572_));
 sky130_fd_sc_hd__a211o_1 _2135_ (.A1(_1224_),
    .A2(_0555_),
    .B1(_0571_),
    .C1(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__o21ai_1 _2136_ (.A1(_0464_),
    .A2(_0509_),
    .B1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(net283),
    .A1(_0574_),
    .S(_0453_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _2138_ (.A(_0575_),
    .X(_0095_));
 sky130_fd_sc_hd__o21ai_1 _2139_ (.A1(_0484_),
    .A2(_0488_),
    .B1(_0470_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_2 _2140_ (.A(_0481_),
    .B(_0474_),
    .Y(_0577_));
 sky130_fd_sc_hd__o22a_1 _2141_ (.A1(_0477_),
    .A2(_0576_),
    .B1(_0577_),
    .B2(_0468_),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_4 _2142_ (.A(_0466_),
    .B(_0488_),
    .Y(_0579_));
 sky130_fd_sc_hd__or2b_1 _2143_ (.A(_0465_),
    .B_N(_0473_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_2 _2144_ (.A(_0465_),
    .B(_0471_),
    .Y(_0581_));
 sky130_fd_sc_hd__and2_1 _2145_ (.A(_0580_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _2146_ (.A(_0491_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__o31a_1 _2147_ (.A1(_0491_),
    .A2(_0479_),
    .A3(_0579_),
    .B1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__and3_4 _2148_ (.A(\inputs.frequency_lut.rng[0] ),
    .B(\inputs.frequency_lut.rng[1] ),
    .C(\inputs.frequency_lut.rng[2] ),
    .X(_0585_));
 sky130_fd_sc_hd__a21oi_4 _2149_ (.A1(_0486_),
    .A2(\inputs.frequency_lut.rng[1] ),
    .B1(\inputs.frequency_lut.rng[2] ),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _2150_ (.A(_0481_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__and2b_1 _2151_ (.A_N(_0465_),
    .B(_0473_),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_1 _2152_ (.A(_0484_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__o32a_1 _2153_ (.A1(_0579_),
    .A2(_0585_),
    .A3(_0587_),
    .B1(_0589_),
    .B2(_0468_),
    .X(_0590_));
 sky130_fd_sc_hd__nor2_2 _2154_ (.A(_0486_),
    .B(_0465_),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _2155_ (.A(_0481_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__a21oi_1 _2156_ (.A1(_0494_),
    .A2(_0497_),
    .B1(_0485_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_1 _2157_ (.A1(_0495_),
    .A2(_0592_),
    .B1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__mux4_1 _2158_ (.A0(_0578_),
    .A1(_0584_),
    .A2(_0590_),
    .A3(_0594_),
    .S0(_0506_),
    .S1(_0508_),
    .X(_0595_));
 sky130_fd_sc_hd__a31o_1 _2159_ (.A1(_0528_),
    .A2(_0529_),
    .A3(_0546_),
    .B1(_0562_),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _2160_ (.A(_0531_),
    .B(_0536_),
    .C(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _2161_ (.A0(_0545_),
    .A1(_0597_),
    .S(_1214_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(_0540_),
    .A1(_0551_),
    .S(_0541_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _2163_ (.A0(_0598_),
    .A1(_0599_),
    .S(_0556_),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _2164_ (.A(_1207_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__mux4_1 _2165_ (.A0(_0532_),
    .A1(_0559_),
    .A2(_0563_),
    .A3(_0568_),
    .S0(_1215_),
    .S1(_0556_),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_4 _2166_ (.A(_0463_),
    .X(_0603_));
 sky130_fd_sc_hd__o21ai_1 _2167_ (.A1(_1224_),
    .A2(_0602_),
    .B1(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__o22a_1 _2168_ (.A1(_0464_),
    .A2(_0595_),
    .B1(_0601_),
    .B2(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_4 _2169_ (.A(_0411_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(net280),
    .A1(_0605_),
    .S(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_1 _2171_ (.A(_0607_),
    .X(_0096_));
 sky130_fd_sc_hd__and4_1 _2172_ (.A(_0531_),
    .B(_0528_),
    .C(_0539_),
    .D(_0547_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(_0597_),
    .A1(_0608_),
    .S(_1214_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(_0552_),
    .A1(_0609_),
    .S(_0554_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _2175_ (.A0(_0542_),
    .A1(_0564_),
    .S(_0556_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(_0610_),
    .A1(_0611_),
    .S(_1207_),
    .X(_0612_));
 sky130_fd_sc_hd__nor2_1 _2177_ (.A(_0485_),
    .B(_0475_),
    .Y(_0613_));
 sky130_fd_sc_hd__a21o_1 _2178_ (.A1(_0489_),
    .A2(_0587_),
    .B1(_0506_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_4 _2179_ (.A(\inputs.frequency_lut.rng[4] ),
    .X(_0615_));
 sky130_fd_sc_hd__clkbuf_4 _2180_ (.A(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__a211o_1 _2181_ (.A1(_0499_),
    .A2(_0489_),
    .B1(_0496_),
    .C1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__o211a_1 _2182_ (.A1(_0613_),
    .A2(_0614_),
    .B1(_0617_),
    .C1(_0508_),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _2183_ (.A(_0616_),
    .B(_0576_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _2184_ (.A(_0468_),
    .B(_0466_),
    .Y(_0620_));
 sky130_fd_sc_hd__nor2_1 _2185_ (.A(_0498_),
    .B(_0471_),
    .Y(_0621_));
 sky130_fd_sc_hd__a31o_1 _2186_ (.A1(_0482_),
    .A2(_0494_),
    .A3(_0620_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o32a_1 _2187_ (.A1(_0586_),
    .A2(_0585_),
    .A3(_0619_),
    .B1(_0622_),
    .B2(_0616_),
    .X(_0623_));
 sky130_fd_sc_hd__o21ai_1 _2188_ (.A1(_0508_),
    .A2(_0623_),
    .B1(_0533_),
    .Y(_0624_));
 sky130_fd_sc_hd__o2bb2a_1 _2189_ (.A1_N(_0464_),
    .A2_N(_0612_),
    .B1(_0618_),
    .B2(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(net222),
    .A1(_0625_),
    .S(_0606_),
    .X(_0626_));
 sky130_fd_sc_hd__clkbuf_1 _2191_ (.A(_0626_),
    .X(_0097_));
 sky130_fd_sc_hd__o221a_1 _2192_ (.A1(\inputs.key_encoder.sync_keys[12] ),
    .A2(_1199_),
    .B1(_0526_),
    .B2(_0523_),
    .C1(_0516_),
    .X(_0627_));
 sky130_fd_sc_hd__or3_1 _2193_ (.A(_0565_),
    .B(_0550_),
    .C(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2194_ (.A0(_0608_),
    .A1(_0628_),
    .S(_1214_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _2195_ (.A0(_0598_),
    .A1(_0629_),
    .S(_0553_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2196_ (.A0(_0532_),
    .A1(_0559_),
    .S(_1215_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(_0599_),
    .A1(_0631_),
    .S(_0556_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(_0630_),
    .A1(_0632_),
    .S(_1207_),
    .X(_0633_));
 sky130_fd_sc_hd__inv_2 _2199_ (.A(_0585_),
    .Y(_0634_));
 sky130_fd_sc_hd__a31o_1 _2200_ (.A1(_0491_),
    .A2(_0494_),
    .A3(_0634_),
    .B1(_0592_),
    .X(_0635_));
 sky130_fd_sc_hd__or2b_1 _2201_ (.A(\inputs.frequency_lut.rng[1] ),
    .B_N(\inputs.frequency_lut.rng[2] ),
    .X(_0636_));
 sky130_fd_sc_hd__nor2_1 _2202_ (.A(_0484_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a31oi_1 _2203_ (.A1(_0580_),
    .A2(_0592_),
    .A3(_0636_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__and2_1 _2204_ (.A(_0468_),
    .B(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__nor3_1 _2205_ (.A(_0579_),
    .B(_0585_),
    .C(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__o22a_1 _2206_ (.A1(_0503_),
    .A2(_0577_),
    .B1(_0582_),
    .B2(_0491_),
    .X(_0641_));
 sky130_fd_sc_hd__mux4_1 _2207_ (.A0(_0635_),
    .A1(_0638_),
    .A2(_0640_),
    .A3(_0641_),
    .S0(_0615_),
    .S1(_0507_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _2208_ (.A(_0603_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__o21ai_1 _2209_ (.A1(_0572_),
    .A2(_0633_),
    .B1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__mux2_1 _2210_ (.A0(net240),
    .A1(_0644_),
    .S(_0606_),
    .X(_0645_));
 sky130_fd_sc_hd__clkbuf_1 _2211_ (.A(_0645_),
    .X(_0098_));
 sky130_fd_sc_hd__nor2_1 _2212_ (.A(_0616_),
    .B(_0480_),
    .Y(_0646_));
 sky130_fd_sc_hd__and3b_2 _2213_ (.A_N(_0473_),
    .B(_0465_),
    .C(_0486_),
    .X(_0647_));
 sky130_fd_sc_hd__nand3_1 _2214_ (.A(_0484_),
    .B(_0494_),
    .C(_0620_),
    .Y(_0648_));
 sky130_fd_sc_hd__o21a_1 _2215_ (.A1(_0485_),
    .A2(_0647_),
    .B1(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__buf_2 _2216_ (.A(\inputs.frequency_lut.rng[5] ),
    .X(_0650_));
 sky130_fd_sc_hd__a21oi_1 _2217_ (.A1(_0646_),
    .A2(_0649_),
    .B1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__o21a_1 _2218_ (.A1(_0646_),
    .A2(_0649_),
    .B1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__a21oi_2 _2219_ (.A1(_0469_),
    .A2(_0471_),
    .B1(_0465_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21a_1 _2220_ (.A1(_0479_),
    .A2(_0653_),
    .B1(_0499_),
    .X(_0654_));
 sky130_fd_sc_hd__o21a_1 _2221_ (.A1(_0502_),
    .A2(_0647_),
    .B1(_0484_),
    .X(_0655_));
 sky130_fd_sc_hd__a21oi_1 _2222_ (.A1(_0491_),
    .A2(_0588_),
    .B1(_0615_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21bo_1 _2223_ (.A1(_0497_),
    .A2(_0587_),
    .B1_N(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_4 _2224_ (.A(_0650_),
    .X(_0658_));
 sky130_fd_sc_hd__o311a_1 _2225_ (.A1(_0506_),
    .A2(_0654_),
    .A3(_0655_),
    .B1(_0657_),
    .C1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _2226_ (.A(_0521_),
    .B(_0527_),
    .Y(_0660_));
 sky130_fd_sc_hd__o21a_1 _2227_ (.A1(_0515_),
    .A2(_0527_),
    .B1(_0546_),
    .X(_0661_));
 sky130_fd_sc_hd__o21ai_1 _2228_ (.A1(_0660_),
    .A2(_0661_),
    .B1(_0534_),
    .Y(_0662_));
 sky130_fd_sc_hd__mux2_1 _2229_ (.A0(_0628_),
    .A1(_0662_),
    .S(_0541_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(_0609_),
    .A1(_0663_),
    .S(_0554_),
    .X(_0664_));
 sky130_fd_sc_hd__nor2_1 _2231_ (.A(_1207_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__o21ai_1 _2232_ (.A1(_1224_),
    .A2(_0555_),
    .B1(_0603_),
    .Y(_0666_));
 sky130_fd_sc_hd__o32a_1 _2233_ (.A1(_0603_),
    .A2(_0652_),
    .A3(_0659_),
    .B1(_0665_),
    .B2(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(net273),
    .A1(_0667_),
    .S(_0606_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_0668_),
    .X(_0099_));
 sky130_fd_sc_hd__or2_1 _2236_ (.A(_0486_),
    .B(_0467_),
    .X(_0669_));
 sky130_fd_sc_hd__a31o_1 _2237_ (.A1(_0498_),
    .A2(_0468_),
    .A3(_0588_),
    .B1(_0592_),
    .X(_0670_));
 sky130_fd_sc_hd__a211o_1 _2238_ (.A1(_0669_),
    .A2(_0582_),
    .B1(_0670_),
    .C1(_0505_),
    .X(_0671_));
 sky130_fd_sc_hd__nor2_1 _2239_ (.A(_0491_),
    .B(_0636_),
    .Y(_0672_));
 sky130_fd_sc_hd__a211o_1 _2240_ (.A1(_0499_),
    .A2(_0496_),
    .B1(_0672_),
    .C1(_0616_),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _2241_ (.A(_0481_),
    .B(_0477_),
    .Y(_0674_));
 sky130_fd_sc_hd__o2bb2a_1 _2242_ (.A1_N(_0495_),
    .A2_N(_0674_),
    .B1(_0485_),
    .B2(_0591_),
    .X(_0675_));
 sky130_fd_sc_hd__or2_1 _2243_ (.A(\inputs.frequency_lut.rng[3] ),
    .B(_0585_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _2244_ (.A(_0577_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__a31o_1 _2245_ (.A1(_0615_),
    .A2(_0494_),
    .A3(_0677_),
    .B1(_0650_),
    .X(_0678_));
 sky130_fd_sc_hd__o21ba_1 _2246_ (.A1(_0616_),
    .A2(_0675_),
    .B1_N(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__a31o_1 _2247_ (.A1(_0658_),
    .A2(_0671_),
    .A3(_0673_),
    .B1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _2248_ (.A(_1208_),
    .B(_0600_),
    .Y(_0681_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(_0548_),
    .A1(_0662_),
    .S(_1215_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(_0629_),
    .A1(_0682_),
    .S(_0554_),
    .X(_0683_));
 sky130_fd_sc_hd__a21oi_1 _2251_ (.A1(_1224_),
    .A2(_0683_),
    .B1(_0533_),
    .Y(_0684_));
 sky130_fd_sc_hd__a22o_1 _2252_ (.A1(_0572_),
    .A2(_0680_),
    .B1(_0681_),
    .B2(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _2253_ (.A0(net294),
    .A1(_0685_),
    .S(_0606_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _2254_ (.A(_0686_),
    .X(_0100_));
 sky130_fd_sc_hd__o21a_1 _2255_ (.A1(_0515_),
    .A2(_0523_),
    .B1(_0527_),
    .X(_0687_));
 sky130_fd_sc_hd__a31o_1 _2256_ (.A1(_0543_),
    .A2(_0535_),
    .A3(_0557_),
    .B1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__and2_1 _2257_ (.A(_0536_),
    .B(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(_0547_),
    .A1(_0689_),
    .S(_0541_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _2259_ (.A(_0556_),
    .B(_0663_),
    .Y(_0691_));
 sky130_fd_sc_hd__o21a_1 _2260_ (.A1(_0556_),
    .A2(_0690_),
    .B1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__nand2_1 _2261_ (.A(_1208_),
    .B(_0610_),
    .Y(_0693_));
 sky130_fd_sc_hd__o211a_1 _2262_ (.A1(_1208_),
    .A2(_0692_),
    .B1(_0693_),
    .C1(_0464_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_1 _2263_ (.A(\inputs.frequency_lut.rng[0] ),
    .B(\inputs.frequency_lut.rng[2] ),
    .X(_0695_));
 sky130_fd_sc_hd__or3_1 _2264_ (.A(_0498_),
    .B(_0653_),
    .C(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _2265_ (.A(_0498_),
    .B(_0467_),
    .Y(_0697_));
 sky130_fd_sc_hd__or2_1 _2266_ (.A(_0472_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_4 _2267_ (.A(_0615_),
    .X(_0699_));
 sky130_fd_sc_hd__a41o_1 _2268_ (.A1(_0699_),
    .A2(_0489_),
    .A3(_0494_),
    .A4(_0583_),
    .B1(_0508_),
    .X(_0700_));
 sky130_fd_sc_hd__a31o_1 _2269_ (.A1(_0506_),
    .A2(_0696_),
    .A3(_0698_),
    .B1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__o21a_1 _2270_ (.A1(_0502_),
    .A2(_0647_),
    .B1(_0499_),
    .X(_0702_));
 sky130_fd_sc_hd__or3b_1 _2271_ (.A(_0702_),
    .B(_0506_),
    .C_N(_0589_),
    .X(_0703_));
 sky130_fd_sc_hd__a311o_1 _2272_ (.A1(_0492_),
    .A2(_0487_),
    .A3(_0497_),
    .B1(_0647_),
    .C1(_0699_),
    .X(_0704_));
 sky130_fd_sc_hd__a21o_1 _2273_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0658_),
    .X(_0705_));
 sky130_fd_sc_hd__a31o_1 _2274_ (.A1(_0572_),
    .A2(_0701_),
    .A3(_0705_),
    .B1(_0910_),
    .X(_0706_));
 sky130_fd_sc_hd__o22a_1 _2275_ (.A1(net159),
    .A2(_1001_),
    .B1(_0694_),
    .B2(_0706_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _2276_ (.A(_0466_),
    .B(_0470_),
    .X(_0707_));
 sky130_fd_sc_hd__o32a_1 _2277_ (.A1(_0491_),
    .A2(_0707_),
    .A3(_0653_),
    .B1(_0579_),
    .B2(_0577_),
    .X(_0708_));
 sky130_fd_sc_hd__nand2_1 _2278_ (.A(_0491_),
    .B(_0470_),
    .Y(_0709_));
 sky130_fd_sc_hd__a22oi_1 _2279_ (.A1(_0482_),
    .A2(_0695_),
    .B1(_0709_),
    .B2(_0581_),
    .Y(_0710_));
 sky130_fd_sc_hd__a21oi_1 _2280_ (.A1(_0493_),
    .A2(_0634_),
    .B1(_0498_),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _2281_ (.A(_0637_),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__o21ba_1 _2282_ (.A1(_0482_),
    .A2(_0472_),
    .B1_N(_0591_),
    .X(_0713_));
 sky130_fd_sc_hd__mux4_1 _2283_ (.A0(_0708_),
    .A1(_0710_),
    .A2(_0712_),
    .A3(_0713_),
    .S0(_0616_),
    .S1(_0508_),
    .X(_0714_));
 sky130_fd_sc_hd__a311o_1 _2284_ (.A1(_1199_),
    .A2(_0522_),
    .A3(_0557_),
    .B1(_0566_),
    .C1(_0558_),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _2285_ (.A(_0541_),
    .B(_0689_),
    .X(_0716_));
 sky130_fd_sc_hd__o21ai_1 _2286_ (.A1(_1215_),
    .A2(_0715_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(_0682_),
    .A1(_0717_),
    .S(_0554_),
    .X(_0718_));
 sky130_fd_sc_hd__and2_1 _2288_ (.A(_1206_),
    .B(_0630_),
    .X(_0719_));
 sky130_fd_sc_hd__a21oi_1 _2289_ (.A1(_1224_),
    .A2(_0718_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(_0714_),
    .A1(_0720_),
    .S(_0603_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(net282),
    .A1(_0721_),
    .S(_0606_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_1 _2292_ (.A(_0722_),
    .X(_0102_));
 sky130_fd_sc_hd__o21a_1 _2293_ (.A1(_0653_),
    .A2(_0695_),
    .B1(_0481_),
    .X(_0723_));
 sky130_fd_sc_hd__or2_1 _2294_ (.A(_0655_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _2295_ (.A(_0498_),
    .B(_0479_),
    .Y(_0725_));
 sky130_fd_sc_hd__a31o_1 _2296_ (.A1(_0482_),
    .A2(_0489_),
    .A3(_0494_),
    .B1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__nand3_1 _2297_ (.A(_0481_),
    .B(_0466_),
    .C(_0470_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _2298_ (.A(_0589_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a21o_1 _2299_ (.A1(_0482_),
    .A2(_0477_),
    .B1(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__a21o_1 _2300_ (.A1(_0470_),
    .A2(_0477_),
    .B1(_0695_),
    .X(_0730_));
 sky130_fd_sc_hd__and2_1 _2301_ (.A(_0484_),
    .B(_0474_),
    .X(_0731_));
 sky130_fd_sc_hd__a21o_1 _2302_ (.A1(_0482_),
    .A2(_0730_),
    .B1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__mux4_1 _2303_ (.A0(_0724_),
    .A1(_0726_),
    .A2(_0729_),
    .A3(_0732_),
    .S0(_0616_),
    .S1(_0650_),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _2304_ (.A(_1208_),
    .B(_0664_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _2305_ (.A(_0527_),
    .B(_0539_),
    .Y(_0735_));
 sky130_fd_sc_hd__mux2_1 _2306_ (.A0(_0715_),
    .A1(_0735_),
    .S(_0541_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _2307_ (.A0(_0690_),
    .A1(_0736_),
    .S(_0554_),
    .X(_0737_));
 sky130_fd_sc_hd__o21a_1 _2308_ (.A1(_1207_),
    .A2(_0737_),
    .B1(_0603_),
    .X(_0738_));
 sky130_fd_sc_hd__a22o_1 _2309_ (.A1(_0572_),
    .A2(_0733_),
    .B1(_0734_),
    .B2(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _2310_ (.A0(net292),
    .A1(_0739_),
    .S(_0606_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_1 _2311_ (.A(_0740_),
    .X(_0103_));
 sky130_fd_sc_hd__or3_1 _2312_ (.A(_0498_),
    .B(_0479_),
    .C(_0591_),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _2313_ (.A(_0468_),
    .B(_0466_),
    .X(_0742_));
 sky130_fd_sc_hd__o21ai_1 _2314_ (.A1(_0477_),
    .A2(_0742_),
    .B1(_0499_),
    .Y(_0743_));
 sky130_fd_sc_hd__a21o_1 _2315_ (.A1(_0741_),
    .A2(_0743_),
    .B1(_0507_),
    .X(_0744_));
 sky130_fd_sc_hd__inv_2 _2316_ (.A(_0579_),
    .Y(_0745_));
 sky130_fd_sc_hd__a221o_1 _2317_ (.A1(_0492_),
    .A2(_0581_),
    .B1(_0731_),
    .B2(_0745_),
    .C1(_0650_),
    .X(_0746_));
 sky130_fd_sc_hd__and3_1 _2318_ (.A(_0699_),
    .B(_0744_),
    .C(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__inv_2 _2319_ (.A(_0653_),
    .Y(_0748_));
 sky130_fd_sc_hd__or3_1 _2320_ (.A(_0498_),
    .B(_0479_),
    .C(_0502_),
    .X(_0749_));
 sky130_fd_sc_hd__a311o_1 _2321_ (.A1(_0497_),
    .A2(_0748_),
    .A3(_0749_),
    .B1(_0621_),
    .C1(_0650_),
    .X(_0750_));
 sky130_fd_sc_hd__or3_1 _2322_ (.A(_0485_),
    .B(_0479_),
    .C(_0502_),
    .X(_0751_));
 sky130_fd_sc_hd__o211ai_1 _2323_ (.A1(_0492_),
    .A2(_0494_),
    .B1(_0751_),
    .C1(_0658_),
    .Y(_0752_));
 sky130_fd_sc_hd__a31o_1 _2324_ (.A1(_0506_),
    .A2(_0750_),
    .A3(_0752_),
    .B1(_0603_),
    .X(_0753_));
 sky130_fd_sc_hd__o211a_2 _2325_ (.A1(_0515_),
    .A2(_0524_),
    .B1(_0536_),
    .C1(_0531_),
    .X(_0754_));
 sky130_fd_sc_hd__o21ai_1 _2326_ (.A1(_0541_),
    .A2(_0735_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(_0717_),
    .A1(_0755_),
    .S(_0554_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(_0683_),
    .A1(_0756_),
    .S(_1224_),
    .X(_0757_));
 sky130_fd_sc_hd__o22ai_1 _2329_ (.A1(_0747_),
    .A2(_0753_),
    .B1(_0757_),
    .B2(_0572_),
    .Y(_0758_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(net295),
    .A1(_0758_),
    .S(_0606_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_0759_),
    .X(_0104_));
 sky130_fd_sc_hd__xnor2_1 _2332_ (.A(_1215_),
    .B(_0754_),
    .Y(_0760_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(_0736_),
    .A1(_0760_),
    .S(_0554_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(_0692_),
    .A1(_0761_),
    .S(_1224_),
    .X(_0762_));
 sky130_fd_sc_hd__o21a_1 _2335_ (.A1(_0586_),
    .A2(_0695_),
    .B1(\inputs.frequency_lut.rng[3] ),
    .X(_0763_));
 sky130_fd_sc_hd__a31o_1 _2336_ (.A1(_0470_),
    .A2(_0471_),
    .A3(_0731_),
    .B1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__a31o_1 _2337_ (.A1(_0481_),
    .A2(_0581_),
    .A3(_0748_),
    .B1(_0615_),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _2338_ (.A(_0491_),
    .B(_0730_),
    .Y(_0766_));
 sky130_fd_sc_hd__o2bb2a_1 _2339_ (.A1_N(_0615_),
    .A2_N(_0764_),
    .B1(_0765_),
    .B2(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__o21ai_1 _2340_ (.A1(_0477_),
    .A2(_0707_),
    .B1(_0485_),
    .Y(_0768_));
 sky130_fd_sc_hd__a32o_1 _2341_ (.A1(_0615_),
    .A2(_0577_),
    .A3(_0768_),
    .B1(_0656_),
    .B2(_0648_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(_0767_),
    .A1(_0769_),
    .S(_0508_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2_1 _2343_ (.A(_0603_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a21o_1 _2344_ (.A1(_0464_),
    .A2(_0762_),
    .B1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(net285),
    .A1(_0772_),
    .S(_0606_),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_1 _2346_ (.A(_0773_),
    .X(_0105_));
 sky130_fd_sc_hd__nor2_1 _2347_ (.A(_0587_),
    .B(_0742_),
    .Y(_0774_));
 sky130_fd_sc_hd__or3_1 _2348_ (.A(_0484_),
    .B(_0579_),
    .C(_0585_),
    .X(_0775_));
 sky130_fd_sc_hd__o21a_1 _2349_ (.A1(_0499_),
    .A2(_0480_),
    .B1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__o21ai_1 _2350_ (.A1(_0479_),
    .A2(_0591_),
    .B1(_0492_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_1 _2351_ (.A(_0749_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21oi_1 _2352_ (.A1(_0492_),
    .A2(_0470_),
    .B1(_0467_),
    .Y(_0779_));
 sky130_fd_sc_hd__mux4_1 _2353_ (.A0(_0774_),
    .A1(_0776_),
    .A2(_0778_),
    .A3(_0779_),
    .S0(_0506_),
    .S1(_0508_),
    .X(_0780_));
 sky130_fd_sc_hd__or3_1 _2354_ (.A(_0541_),
    .B(_0556_),
    .C(_0754_),
    .X(_0781_));
 sky130_fd_sc_hd__o21ai_1 _2355_ (.A1(_0554_),
    .A2(_0755_),
    .B1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__nor2_1 _2356_ (.A(_1207_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__a211o_1 _2357_ (.A1(_1207_),
    .A2(_0718_),
    .B1(_0783_),
    .C1(_0572_),
    .X(_0784_));
 sky130_fd_sc_hd__o21ai_1 _2358_ (.A1(_0464_),
    .A2(_0780_),
    .B1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(net288),
    .A1(_0785_),
    .S(_0606_),
    .X(_0786_));
 sky130_fd_sc_hd__clkbuf_1 _2360_ (.A(_0786_),
    .X(_0106_));
 sky130_fd_sc_hd__and2_1 _2361_ (.A(_0581_),
    .B(_0748_),
    .X(_0787_));
 sky130_fd_sc_hd__o22ai_1 _2362_ (.A1(_0472_),
    .A2(_0577_),
    .B1(_0787_),
    .B2(_0492_),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_1 _2363_ (.A(_0615_),
    .B(_0676_),
    .Y(_0789_));
 sky130_fd_sc_hd__a311o_1 _2364_ (.A1(_0506_),
    .A2(_0499_),
    .A3(_0730_),
    .B1(_0789_),
    .C1(_0650_),
    .X(_0790_));
 sky130_fd_sc_hd__a21o_1 _2365_ (.A1(_0699_),
    .A2(_0788_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _2366_ (.A(_0485_),
    .B(_0586_),
    .Y(_0792_));
 sky130_fd_sc_hd__o311a_1 _2367_ (.A1(_0482_),
    .A2(_0586_),
    .A3(_0585_),
    .B1(_0697_),
    .C1(_0505_),
    .X(_0793_));
 sky130_fd_sc_hd__a311o_1 _2368_ (.A1(_0699_),
    .A2(_0727_),
    .A3(_0792_),
    .B1(_0793_),
    .C1(_0508_),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _2369_ (.A(_1206_),
    .B(_0754_),
    .X(_0795_));
 sky130_fd_sc_hd__o211a_1 _2370_ (.A1(_1224_),
    .A2(_0737_),
    .B1(_0795_),
    .C1(_0463_),
    .X(_0796_));
 sky130_fd_sc_hd__a31o_1 _2371_ (.A1(_0572_),
    .A2(_0791_),
    .A3(_0794_),
    .B1(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_4 _2372_ (.A(_0994_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(net256),
    .A1(_0797_),
    .S(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_1 _2374_ (.A(_0799_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(_0754_),
    .A1(_0756_),
    .S(_1207_),
    .X(_0800_));
 sky130_fd_sc_hd__a31o_1 _2376_ (.A1(_0699_),
    .A2(_0698_),
    .A3(_0792_),
    .B1(_0789_),
    .X(_0801_));
 sky130_fd_sc_hd__o211ai_1 _2377_ (.A1(_0485_),
    .A2(_0480_),
    .B1(_0741_),
    .C1(_0506_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _2378_ (.A1(_0498_),
    .A2(_0487_),
    .B1(_0505_),
    .Y(_0803_));
 sky130_fd_sc_hd__o21ai_1 _2379_ (.A1(_0579_),
    .A2(_0676_),
    .B1(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__a21oi_1 _2380_ (.A1(_0802_),
    .A2(_0804_),
    .B1(_0658_),
    .Y(_0805_));
 sky130_fd_sc_hd__a211o_1 _2381_ (.A1(_0658_),
    .A2(_0801_),
    .B1(_0805_),
    .C1(_0603_),
    .X(_0806_));
 sky130_fd_sc_hd__o21ai_1 _2382_ (.A1(_0572_),
    .A2(_0800_),
    .B1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(net286),
    .A1(_0807_),
    .S(_0798_),
    .X(_0808_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_0808_),
    .X(_0108_));
 sky130_fd_sc_hd__a41o_1 _2385_ (.A1(_0481_),
    .A2(_0486_),
    .A3(_0473_),
    .A4(_0466_),
    .B1(_0615_),
    .X(_0809_));
 sky130_fd_sc_hd__a21oi_1 _2386_ (.A1(_0482_),
    .A2(_0586_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__o21a_1 _2387_ (.A1(_0482_),
    .A2(_0467_),
    .B1(_0803_),
    .X(_0811_));
 sky130_fd_sc_hd__a21oi_1 _2388_ (.A1(_0696_),
    .A2(_0810_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__a41o_1 _2389_ (.A1(_0616_),
    .A2(_0499_),
    .A3(_0467_),
    .A4(_0476_),
    .B1(_0507_),
    .X(_0813_));
 sky130_fd_sc_hd__o221a_1 _2390_ (.A1(_0658_),
    .A2(_0812_),
    .B1(_0813_),
    .B2(_0789_),
    .C1(_0533_),
    .X(_0814_));
 sky130_fd_sc_hd__a31o_1 _2391_ (.A1(_1208_),
    .A2(_0464_),
    .A3(_0761_),
    .B1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(net230),
    .A1(_0815_),
    .S(_0798_),
    .X(_0816_));
 sky130_fd_sc_hd__clkbuf_1 _2393_ (.A(_0816_),
    .X(_0109_));
 sky130_fd_sc_hd__and4_1 _2394_ (.A(_0650_),
    .B(_0616_),
    .C(_0499_),
    .D(_0647_),
    .X(_0817_));
 sky130_fd_sc_hd__o211a_1 _2395_ (.A1(_0585_),
    .A2(_0731_),
    .B1(_0505_),
    .C1(_0487_),
    .X(_0818_));
 sky130_fd_sc_hd__o21a_1 _2396_ (.A1(_0803_),
    .A2(_0818_),
    .B1(_0508_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_1 _2397_ (.A1(_0817_),
    .A2(_0819_),
    .B1(_0533_),
    .X(_0820_));
 sky130_fd_sc_hd__a31o_1 _2398_ (.A1(_1208_),
    .A2(_0464_),
    .A3(_0782_),
    .B1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(net239),
    .A1(_0821_),
    .S(_0798_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(_0822_),
    .X(_0110_));
 sky130_fd_sc_hd__nand2_1 _2401_ (.A(_0650_),
    .B(_0639_),
    .Y(_0823_));
 sky130_fd_sc_hd__a21o_1 _2402_ (.A1(_0485_),
    .A2(_0586_),
    .B1(_0809_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(_0650_),
    .A1(_0823_),
    .S(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nor2_1 _2404_ (.A(_0603_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a41o_1 _2405_ (.A1(_1208_),
    .A2(_0464_),
    .A3(_0556_),
    .A4(_0760_),
    .B1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(net232),
    .A1(_0827_),
    .S(_0798_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _2407_ (.A(_0828_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _2408_ (.A(_0910_),
    .X(_0829_));
 sky130_fd_sc_hd__or3b_1 _2409_ (.A(\inputs.octave_fsm.state[2] ),
    .B(_0754_),
    .C_N(_1205_),
    .X(_0830_));
 sky130_fd_sc_hd__or4_1 _2410_ (.A(_0658_),
    .B(_0699_),
    .C(_0464_),
    .D(_0792_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_4 _2411_ (.A(_0910_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_1 _2412_ (.A1(_0830_),
    .A2(_0831_),
    .B1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a21o_1 _2413_ (.A1(net122),
    .A2(_0829_),
    .B1(_0833_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2414_ (.A0(net311),
    .A1(\outputs.div.m[0] ),
    .S(_0798_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _2415_ (.A(_0834_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(\outputs.divider_buffer[1] ),
    .A1(\outputs.div.m[1] ),
    .S(_0798_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_1 _2417_ (.A(_0835_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(\outputs.divider_buffer[2] ),
    .A1(\outputs.div.m[2] ),
    .S(_0798_),
    .X(_0836_));
 sky130_fd_sc_hd__clkbuf_1 _2419_ (.A(_0836_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(\outputs.divider_buffer[3] ),
    .A1(\outputs.div.m[3] ),
    .S(_0798_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _2421_ (.A(_0837_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(\outputs.divider_buffer[4] ),
    .A1(\outputs.div.m[4] ),
    .S(_0798_),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_1 _2423_ (.A(_0838_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _2424_ (.A(_0994_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(\outputs.divider_buffer[5] ),
    .A1(\outputs.div.m[5] ),
    .S(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _2426_ (.A(_0840_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(net309),
    .A1(net297),
    .S(_0839_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _2428_ (.A(_0841_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(\outputs.divider_buffer[7] ),
    .A1(\outputs.div.m[7] ),
    .S(_0839_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(_0842_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(\outputs.divider_buffer[8] ),
    .A1(\outputs.div.m[8] ),
    .S(_0839_),
    .X(_0843_));
 sky130_fd_sc_hd__clkbuf_1 _2432_ (.A(_0843_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(\outputs.divider_buffer[9] ),
    .A1(\outputs.div.m[9] ),
    .S(_0839_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _2434_ (.A(_0844_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(\outputs.divider_buffer[10] ),
    .A1(\outputs.div.m[10] ),
    .S(_0839_),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _2436_ (.A(_0845_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2437_ (.A0(\outputs.divider_buffer[11] ),
    .A1(\outputs.div.m[11] ),
    .S(_0839_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _2438_ (.A(_0846_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(\outputs.divider_buffer[12] ),
    .A1(\outputs.div.m[12] ),
    .S(_0839_),
    .X(_0847_));
 sky130_fd_sc_hd__clkbuf_1 _2440_ (.A(_0847_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(\outputs.divider_buffer[13] ),
    .A1(\outputs.div.m[13] ),
    .S(_0839_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_1 _2442_ (.A(_0848_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(net310),
    .A1(\outputs.div.m[14] ),
    .S(_0839_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_1 _2444_ (.A(_0849_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_4 _2445_ (.A(_0994_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _2446_ (.A0(\outputs.divider_buffer[15] ),
    .A1(\outputs.div.m[15] ),
    .S(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__clkbuf_1 _2447_ (.A(_0851_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(\outputs.divider_buffer[16] ),
    .A1(\outputs.div.m[16] ),
    .S(_0850_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_1 _2449_ (.A(_0852_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(net312),
    .A1(\outputs.div.m[17] ),
    .S(_0850_),
    .X(_0853_));
 sky130_fd_sc_hd__clkbuf_1 _2451_ (.A(_0853_),
    .X(_0130_));
 sky130_fd_sc_hd__a21o_1 _2452_ (.A1(net128),
    .A2(_0829_),
    .B1(_0397_),
    .X(_0131_));
 sky130_fd_sc_hd__a21o_1 _2453_ (.A1(net125),
    .A2(_0829_),
    .B1(_0399_),
    .X(_0132_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(net110),
    .A2(_0829_),
    .B1(_0401_),
    .X(_0133_));
 sky130_fd_sc_hd__a21o_1 _2455_ (.A1(net108),
    .A2(_0829_),
    .B1(_0402_),
    .X(_0134_));
 sky130_fd_sc_hd__a21o_1 _2456_ (.A1(net105),
    .A2(_0829_),
    .B1(_0403_),
    .X(_0135_));
 sky130_fd_sc_hd__a21o_1 _2457_ (.A1(net123),
    .A2(_0829_),
    .B1(_0404_),
    .X(_0136_));
 sky130_fd_sc_hd__a21o_1 _2458_ (.A1(net101),
    .A2(_0829_),
    .B1(_0406_),
    .X(_0137_));
 sky130_fd_sc_hd__a21o_1 _2459_ (.A1(net120),
    .A2(_0829_),
    .B1(_0407_),
    .X(_0138_));
 sky130_fd_sc_hd__a21o_1 _2460_ (.A1(net129),
    .A2(_0829_),
    .B1(_0408_),
    .X(_0139_));
 sky130_fd_sc_hd__a21o_1 _2461_ (.A1(net116),
    .A2(_0832_),
    .B1(_0409_),
    .X(_0140_));
 sky130_fd_sc_hd__a21o_1 _2462_ (.A1(net131),
    .A2(_0832_),
    .B1(_0410_),
    .X(_0141_));
 sky130_fd_sc_hd__a21o_1 _2463_ (.A1(net112),
    .A2(_0832_),
    .B1(_0412_),
    .X(_0142_));
 sky130_fd_sc_hd__a21o_1 _2464_ (.A1(net103),
    .A2(_0832_),
    .B1(_0413_),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _2465_ (.A1(net114),
    .A2(_0832_),
    .B1(_0414_),
    .X(_0144_));
 sky130_fd_sc_hd__a21o_1 _2466_ (.A1(net106),
    .A2(_0832_),
    .B1(_0415_),
    .X(_0145_));
 sky130_fd_sc_hd__a21o_1 _2467_ (.A1(net135),
    .A2(_0832_),
    .B1(_0416_),
    .X(_0146_));
 sky130_fd_sc_hd__a21o_1 _2468_ (.A1(net126),
    .A2(_0832_),
    .B1(_0417_),
    .X(_0147_));
 sky130_fd_sc_hd__a21o_1 _2469_ (.A1(net111),
    .A2(_0832_),
    .B1(_0418_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2470_ (.A0(net265),
    .A1(\outputs.sig_gen.count[0] ),
    .S(_0850_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_1 _2471_ (.A(_0854_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2472_ (.A0(net281),
    .A1(\outputs.sig_gen.count[1] ),
    .S(_0850_),
    .X(_0855_));
 sky130_fd_sc_hd__clkbuf_1 _2473_ (.A(_0855_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(net279),
    .A1(\outputs.sig_gen.count[2] ),
    .S(_0850_),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_1 _2475_ (.A(_0856_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(net267),
    .A1(\outputs.sig_gen.count[3] ),
    .S(_0850_),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_1 _2477_ (.A(_0857_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(net274),
    .A1(\outputs.sig_gen.count[4] ),
    .S(_0850_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_1 _2479_ (.A(_0858_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(net270),
    .A1(\outputs.sig_gen.count[5] ),
    .S(_0850_),
    .X(_0859_));
 sky130_fd_sc_hd__clkbuf_1 _2481_ (.A(_0859_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(net264),
    .A1(\outputs.sig_gen.count[6] ),
    .S(_0850_),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_1 _2483_ (.A(_0860_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_4 _2484_ (.A(_0994_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(net277),
    .A1(\outputs.sig_gen.count[7] ),
    .S(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_0862_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(net269),
    .A1(\outputs.sig_gen.count[8] ),
    .S(_0861_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_0863_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2489_ (.A0(net272),
    .A1(\outputs.sig_gen.count[9] ),
    .S(_0861_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_1 _2490_ (.A(_0864_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2491_ (.A0(net276),
    .A1(\outputs.sig_gen.count[10] ),
    .S(_0861_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _2492_ (.A(_0865_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(net275),
    .A1(\outputs.sig_gen.count[11] ),
    .S(_0861_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(_0866_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2495_ (.A0(net289),
    .A1(\outputs.sig_gen.count[12] ),
    .S(_0861_),
    .X(_0867_));
 sky130_fd_sc_hd__clkbuf_1 _2496_ (.A(_0867_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(net306),
    .A1(\outputs.sig_gen.count[13] ),
    .S(_0861_),
    .X(_0868_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(_0868_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(net284),
    .A1(\outputs.sig_gen.count[14] ),
    .S(_0861_),
    .X(_0869_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_0869_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(net287),
    .A1(\outputs.sig_gen.count[15] ),
    .S(_0861_),
    .X(_0870_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_0870_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(net291),
    .A1(\outputs.sig_gen.count[16] ),
    .S(_0861_),
    .X(_0871_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(_0871_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_4 _2505_ (.A(_0994_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(net290),
    .A1(\outputs.sig_gen.count[17] ),
    .S(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_0873_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(\outputs.shaper.count[0] ),
    .A1(net128),
    .S(_0872_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(_0874_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(net300),
    .A1(net125),
    .S(_0872_),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_0875_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\outputs.shaper.count[2] ),
    .A1(net110),
    .S(_0872_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_0876_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\outputs.shaper.count[3] ),
    .A1(net108),
    .S(_0872_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_0877_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(\outputs.shaper.count[4] ),
    .A1(net105),
    .S(_0872_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_0878_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(\outputs.shaper.count[5] ),
    .A1(net123),
    .S(_0872_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_0879_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\outputs.shaper.count[6] ),
    .A1(net101),
    .S(_0872_),
    .X(_0880_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_0880_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net304),
    .A1(net120),
    .S(_0872_),
    .X(_0881_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_0881_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net301),
    .A1(net129),
    .S(_0872_),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(_0882_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\outputs.shaper.count[9] ),
    .A1(net116),
    .S(_0396_),
    .X(_0883_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_0883_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(\outputs.shaper.count[10] ),
    .A1(net131),
    .S(_0396_),
    .X(_0884_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(_0884_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net298),
    .A1(net112),
    .S(_0396_),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(_0885_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net299),
    .A1(net103),
    .S(_0396_),
    .X(_0886_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(_0886_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\outputs.shaper.count[13] ),
    .A1(net114),
    .S(_0396_),
    .X(_0887_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_0887_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\outputs.shaper.count[14] ),
    .A1(net106),
    .S(_0396_),
    .X(_0888_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(_0888_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\outputs.shaper.count[15] ),
    .A1(net135),
    .S(_0396_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_0889_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\outputs.shaper.count[16] ),
    .A1(net126),
    .S(_0396_),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(_0890_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(net305),
    .A1(net111),
    .S(_0396_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_0891_),
    .X(_0184_));
 sky130_fd_sc_hd__xnor2_1 _2544_ (.A(_0658_),
    .B(_0699_),
    .Y(_0892_));
 sky130_fd_sc_hd__xnor2_1 _2545_ (.A(_0492_),
    .B(_1093_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_1 _2546_ (.A(_0892_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_4 _2547_ (.A(_0951_),
    .B(_0572_),
    .Y(_0895_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(_0894_),
    .A1(_0486_),
    .S(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0896_),
    .X(_0185_));
 sky130_fd_sc_hd__xor2_1 _2550_ (.A(_0486_),
    .B(_1093_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(_0897_),
    .A1(_0473_),
    .S(_0895_),
    .X(_0898_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_0898_),
    .X(_0186_));
 sky130_fd_sc_hd__xor2_1 _2553_ (.A(_0473_),
    .B(_1093_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(_0899_),
    .A1(_0467_),
    .S(_0895_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_1 _2555_ (.A(_0900_),
    .X(_0187_));
 sky130_fd_sc_hd__xor2_1 _2556_ (.A(_0467_),
    .B(_1093_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(_0901_),
    .A1(_0492_),
    .S(_0895_),
    .X(_0902_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_0902_),
    .X(_0188_));
 sky130_fd_sc_hd__nand2_1 _2559_ (.A(_0699_),
    .B(_0895_),
    .Y(_0903_));
 sky130_fd_sc_hd__o21ai_1 _2560_ (.A1(_0895_),
    .A2(_0893_),
    .B1(_0903_),
    .Y(_0189_));
 sky130_fd_sc_hd__xor2_1 _2561_ (.A(_0699_),
    .B(_1093_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(_0904_),
    .A1(_0658_),
    .S(_0895_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(_0905_),
    .X(_0190_));
 sky130_fd_sc_hd__dfrtp_1 _2564_ (.CLK(clknet_leaf_27_clk),
    .D(\outputs.sample_rate.next_count[0] ),
    .RESET_B(net31),
    .Q(\outputs.sample_rate.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2565_ (.CLK(clknet_leaf_26_clk),
    .D(\outputs.sample_rate.next_count[1] ),
    .RESET_B(net31),
    .Q(\outputs.sample_rate.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2566_ (.CLK(clknet_leaf_27_clk),
    .D(net158),
    .RESET_B(net31),
    .Q(\outputs.sample_rate.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2567_ (.CLK(clknet_leaf_27_clk),
    .D(\outputs.sample_rate.next_count[3] ),
    .RESET_B(net30),
    .Q(\outputs.sample_rate.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2568_ (.CLK(clknet_leaf_28_clk),
    .D(\outputs.sample_rate.next_count[4] ),
    .RESET_B(net30),
    .Q(\outputs.sample_rate.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2569_ (.CLK(clknet_leaf_27_clk),
    .D(\outputs.sample_rate.next_count[5] ),
    .RESET_B(net30),
    .Q(\outputs.sample_rate.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2570_ (.CLK(clknet_leaf_25_clk),
    .D(\outputs.sample_rate.next_count[6] ),
    .RESET_B(net30),
    .Q(\outputs.sample_rate.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2571_ (.CLK(clknet_leaf_22_clk),
    .D(\outputs.sample_rate.next_count[7] ),
    .RESET_B(net34),
    .Q(\outputs.sample_rate.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2572_ (.CLK(clknet_leaf_24_clk),
    .D(\inputs.wavetype_fsm.next_state[0] ),
    .RESET_B(net30),
    .Q(\inputs.wavetype_fsm.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2573_ (.CLK(clknet_leaf_24_clk),
    .D(net255),
    .RESET_B(net34),
    .Q(\inputs.wavetype_fsm.state[1] ));
 sky130_fd_sc_hd__dfstp_1 _2574_ (.CLK(clknet_leaf_36_clk),
    .D(\inputs.random_note_generator.feedback ),
    .SET_B(net24),
    .Q(\inputs.random_note_generator.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2575_ (.CLK(clknet_leaf_36_clk),
    .D(net87),
    .RESET_B(net24),
    .Q(\inputs.random_note_generator.out[1] ));
 sky130_fd_sc_hd__dfstp_1 _2576_ (.CLK(clknet_leaf_36_clk),
    .D(net81),
    .SET_B(net24),
    .Q(\inputs.random_note_generator.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2577_ (.CLK(clknet_leaf_36_clk),
    .D(net85),
    .RESET_B(net24),
    .Q(\inputs.random_note_generator.out[3] ));
 sky130_fd_sc_hd__dfstp_1 _2578_ (.CLK(clknet_leaf_36_clk),
    .D(net79),
    .SET_B(net24),
    .Q(\inputs.random_note_generator.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2579_ (.CLK(clknet_leaf_36_clk),
    .D(net84),
    .RESET_B(net26),
    .Q(\inputs.random_note_generator.out[5] ));
 sky130_fd_sc_hd__dfstp_1 _2580_ (.CLK(clknet_leaf_0_clk),
    .D(net69),
    .SET_B(net26),
    .Q(\inputs.random_note_generator.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2581_ (.CLK(clknet_leaf_36_clk),
    .D(net83),
    .RESET_B(net25),
    .Q(\inputs.random_note_generator.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2582_ (.CLK(clknet_leaf_0_clk),
    .D(net68),
    .RESET_B(net25),
    .Q(\inputs.random_note_generator.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2583_ (.CLK(clknet_leaf_36_clk),
    .D(net70),
    .RESET_B(net24),
    .Q(\inputs.random_note_generator.out[9] ));
 sky130_fd_sc_hd__dfstp_1 _2584_ (.CLK(clknet_leaf_36_clk),
    .D(net80),
    .SET_B(net24),
    .Q(\inputs.random_note_generator.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2585_ (.CLK(clknet_leaf_36_clk),
    .D(net93),
    .RESET_B(net24),
    .Q(\inputs.random_note_generator.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2586_ (.CLK(clknet_leaf_36_clk),
    .D(net77),
    .RESET_B(net24),
    .Q(\inputs.random_note_generator.out[12] ));
 sky130_fd_sc_hd__dfstp_1 _2587_ (.CLK(clknet_leaf_35_clk),
    .D(net88),
    .SET_B(net24),
    .Q(\inputs.random_note_generator.out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2588_ (.CLK(clknet_leaf_35_clk),
    .D(net91),
    .RESET_B(net22),
    .Q(\inputs.random_note_generator.out[14] ));
 sky130_fd_sc_hd__dfstp_1 _2589_ (.CLK(clknet_leaf_35_clk),
    .D(net74),
    .SET_B(net22),
    .Q(\inputs.random_note_generator.out[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2590_ (.CLK(clknet_leaf_29_clk),
    .D(_0000_),
    .RESET_B(net32),
    .Q(\inputs.octave_fsm.state[0] ));
 sky130_fd_sc_hd__dfstp_2 _2591_ (.CLK(clknet_leaf_33_clk),
    .D(_0001_),
    .SET_B(net23),
    .Q(\inputs.octave_fsm.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2592_ (.CLK(clknet_leaf_29_clk),
    .D(_0002_),
    .RESET_B(net32),
    .Q(\inputs.octave_fsm.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _2593_ (.CLK(clknet_leaf_14_clk),
    .D(\inputs.random_update_clock.next_count[0] ),
    .SET_B(net60),
    .Q(\inputs.random_update_clock.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2594_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[1] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2595_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[2] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2596_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[3] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2597_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[4] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2598_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[5] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2599_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[6] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2600_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[7] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2601_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[8] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2602_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[9] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2603_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[10] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2604_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[11] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2605_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.random_update_clock.next_count[12] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2606_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.random_update_clock.next_count[13] ),
    .RESET_B(net60),
    .Q(\inputs.random_update_clock.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2607_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.random_update_clock.next_count[14] ),
    .RESET_B(net61),
    .Q(\inputs.random_update_clock.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2608_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.random_update_clock.next_count[15] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2609_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[16] ),
    .RESET_B(net55),
    .Q(\inputs.random_update_clock.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2610_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[17] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2611_ (.CLK(clknet_leaf_17_clk),
    .D(\inputs.random_update_clock.next_count[18] ),
    .RESET_B(net55),
    .Q(\inputs.random_update_clock.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2612_ (.CLK(clknet_leaf_18_clk),
    .D(\inputs.random_update_clock.next_count[19] ),
    .RESET_B(net55),
    .Q(\inputs.random_update_clock.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2613_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.random_update_clock.next_count[20] ),
    .RESET_B(net59),
    .Q(\inputs.random_update_clock.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2614_ (.CLK(clknet_leaf_16_clk),
    .D(\inputs.random_update_clock.next_count[21] ),
    .RESET_B(net61),
    .Q(\inputs.random_update_clock.count[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2615_ (.CLK(clknet_leaf_16_clk),
    .D(net119),
    .RESET_B(net61),
    .Q(\inputs.random_update_clock.count[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2616_ (.CLK(clknet_leaf_25_clk),
    .D(net147),
    .RESET_B(net30),
    .Q(\inputs.mode_edge.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2617_ (.CLK(clknet_leaf_25_clk),
    .D(\inputs.mode_edge.ff_in ),
    .RESET_B(net30),
    .Q(\inputs.mode_edge.det_edge ));
 sky130_fd_sc_hd__dfrtp_1 _2618_ (.CLK(clknet_leaf_27_clk),
    .D(\inputs.down.in ),
    .RESET_B(net31),
    .Q(\inputs.down.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2619_ (.CLK(clknet_leaf_28_clk),
    .D(\inputs.down.ff_in ),
    .RESET_B(net32),
    .Q(\inputs.down.det_edge ));
 sky130_fd_sc_hd__dfrtp_1 _2620_ (.CLK(clknet_leaf_28_clk),
    .D(net92),
    .RESET_B(net30),
    .Q(\inputs.up.ff_out ));
 sky130_fd_sc_hd__dfrtp_1 _2621_ (.CLK(clknet_leaf_28_clk),
    .D(\inputs.up.ff_in ),
    .RESET_B(net31),
    .Q(\inputs.octave_fsm.octave_key_up ));
 sky130_fd_sc_hd__dfrtp_1 _2622_ (.CLK(clknet_leaf_25_clk),
    .D(net94),
    .RESET_B(net30),
    .Q(\inputs.key_encoder.sync_keys[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2623_ (.CLK(clknet_leaf_29_clk),
    .D(net82),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2624_ (.CLK(clknet_leaf_28_clk),
    .D(net72),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2625_ (.CLK(clknet_leaf_29_clk),
    .D(net66),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2626_ (.CLK(clknet_leaf_14_clk),
    .D(net78),
    .RESET_B(net58),
    .Q(\inputs.key_encoder.sync_keys[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2627_ (.CLK(clknet_leaf_24_clk),
    .D(net65),
    .RESET_B(net34),
    .Q(\inputs.key_encoder.sync_keys[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2628_ (.CLK(clknet_leaf_36_clk),
    .D(net90),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2629_ (.CLK(clknet_leaf_15_clk),
    .D(net64),
    .RESET_B(net58),
    .Q(\inputs.key_encoder.sync_keys[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2630_ (.CLK(clknet_leaf_29_clk),
    .D(net76),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2631_ (.CLK(clknet_leaf_36_clk),
    .D(net71),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2632_ (.CLK(clknet_leaf_30_clk),
    .D(net95),
    .RESET_B(net33),
    .Q(\inputs.key_encoder.sync_keys[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2633_ (.CLK(clknet_leaf_35_clk),
    .D(net73),
    .RESET_B(net22),
    .Q(\inputs.key_encoder.sync_keys[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2634_ (.CLK(clknet_leaf_0_clk),
    .D(net63),
    .RESET_B(net25),
    .Q(\inputs.key_encoder.sync_keys[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2635_ (.CLK(clknet_leaf_33_clk),
    .D(net86),
    .RESET_B(net23),
    .Q(\inputs.key_encoder.sync_keys[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2636_ (.CLK(clknet_leaf_25_clk),
    .D(net67),
    .RESET_B(net30),
    .Q(\inputs.key_encoder.sync_keys[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2637_ (.CLK(clknet_leaf_30_clk),
    .D(net134),
    .RESET_B(net32),
    .Q(\inputs.key_encoder.sync_keys[15] ));
 sky130_fd_sc_hd__dfrtp_2 _2638_ (.CLK(clknet_leaf_26_clk),
    .D(net89),
    .RESET_B(net31),
    .Q(\inputs.key_encoder.octave_key_up ));
 sky130_fd_sc_hd__dfrtp_1 _2639_ (.CLK(clknet_leaf_15_clk),
    .D(\inputs.keypad[0] ),
    .RESET_B(net60),
    .Q(\inputs.keypad_synchronizer.half_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2640_ (.CLK(clknet_leaf_34_clk),
    .D(\inputs.keypad[1] ),
    .RESET_B(net22),
    .Q(\inputs.keypad_synchronizer.half_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2641_ (.CLK(clknet_leaf_27_clk),
    .D(\inputs.keypad[2] ),
    .RESET_B(net31),
    .Q(\inputs.keypad_synchronizer.half_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2642_ (.CLK(clknet_leaf_33_clk),
    .D(\inputs.keypad[3] ),
    .RESET_B(net23),
    .Q(\inputs.keypad_synchronizer.half_sync[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2643_ (.CLK(clknet_leaf_8_clk),
    .D(\inputs.keypad[4] ),
    .RESET_B(net49),
    .Q(\inputs.keypad_synchronizer.half_sync[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2644_ (.CLK(clknet_leaf_23_clk),
    .D(\inputs.keypad[5] ),
    .RESET_B(net36),
    .Q(\inputs.keypad_synchronizer.half_sync[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2645_ (.CLK(clknet_leaf_6_clk),
    .D(\inputs.keypad[6] ),
    .RESET_B(net45),
    .Q(\inputs.keypad_synchronizer.half_sync[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2646_ (.CLK(clknet_leaf_14_clk),
    .D(\inputs.keypad[7] ),
    .RESET_B(net58),
    .Q(\inputs.keypad_synchronizer.half_sync[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2647_ (.CLK(clknet_leaf_29_clk),
    .D(\inputs.keypad[8] ),
    .RESET_B(net32),
    .Q(\inputs.keypad_synchronizer.half_sync[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2648_ (.CLK(clknet_leaf_3_clk),
    .D(\inputs.keypad[9] ),
    .RESET_B(net39),
    .Q(\inputs.keypad_synchronizer.half_sync[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2649_ (.CLK(clknet_leaf_13_clk),
    .D(\inputs.keypad[10] ),
    .RESET_B(net58),
    .Q(\inputs.keypad_synchronizer.half_sync[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2650_ (.CLK(clknet_leaf_35_clk),
    .D(\inputs.keypad[11] ),
    .RESET_B(net22),
    .Q(\inputs.keypad_synchronizer.half_sync[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2651_ (.CLK(clknet_leaf_37_clk),
    .D(\inputs.keypad[12] ),
    .RESET_B(net25),
    .Q(\inputs.keypad_synchronizer.half_sync[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2652_ (.CLK(clknet_leaf_34_clk),
    .D(\inputs.keypad[13] ),
    .RESET_B(net22),
    .Q(\inputs.keypad_synchronizer.half_sync[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2653_ (.CLK(clknet_leaf_26_clk),
    .D(\inputs.keypad[14] ),
    .RESET_B(net31),
    .Q(\inputs.keypad_synchronizer.half_sync[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2654_ (.CLK(clknet_leaf_5_clk),
    .D(\inputs.keypad[15] ),
    .RESET_B(net44),
    .Q(\inputs.keypad_synchronizer.half_sync[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2655_ (.CLK(clknet_leaf_18_clk),
    .D(\inputs.keypad[16] ),
    .RESET_B(net55),
    .Q(\inputs.keypad_synchronizer.half_sync[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2656_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.pwm_unff ),
    .RESET_B(net34),
    .Q(\outputs.output_gen.pwm_ff ));
 sky130_fd_sc_hd__dfrtp_1 _2657_ (.CLK(clknet_leaf_20_clk),
    .D(_0003_),
    .RESET_B(net53),
    .Q(\outputs.div.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2658_ (.CLK(clknet_leaf_23_clk),
    .D(_0004_),
    .RESET_B(net36),
    .Q(\outputs.div.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2659_ (.CLK(clknet_leaf_22_clk),
    .D(_0005_),
    .RESET_B(net36),
    .Q(\outputs.div.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2660_ (.CLK(clknet_leaf_22_clk),
    .D(_0006_),
    .RESET_B(net34),
    .Q(\outputs.div.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2661_ (.CLK(clknet_leaf_22_clk),
    .D(_0007_),
    .RESET_B(net34),
    .Q(\outputs.div.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2662_ (.CLK(clknet_leaf_22_clk),
    .D(_0008_),
    .RESET_B(net33),
    .Q(\outputs.div.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2663_ (.CLK(clknet_leaf_30_clk),
    .D(_0009_),
    .RESET_B(net33),
    .Q(\outputs.div.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2664_ (.CLK(clknet_leaf_21_clk),
    .D(_0010_),
    .RESET_B(net33),
    .Q(\outputs.div.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2665_ (.CLK(clknet_leaf_31_clk),
    .D(_0011_),
    .RESET_B(net33),
    .Q(\outputs.div.a[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2666_ (.CLK(clknet_leaf_21_clk),
    .D(_0012_),
    .RESET_B(net33),
    .Q(\outputs.div.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2667_ (.CLK(clknet_leaf_21_clk),
    .D(_0013_),
    .RESET_B(net33),
    .Q(\outputs.div.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2668_ (.CLK(clknet_leaf_19_clk),
    .D(_0014_),
    .RESET_B(net51),
    .Q(\outputs.div.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2669_ (.CLK(clknet_leaf_20_clk),
    .D(_0015_),
    .RESET_B(net51),
    .Q(\outputs.div.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2670_ (.CLK(clknet_leaf_19_clk),
    .D(_0016_),
    .RESET_B(net51),
    .Q(\outputs.div.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2671_ (.CLK(clknet_leaf_20_clk),
    .D(_0017_),
    .RESET_B(net51),
    .Q(\outputs.div.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2672_ (.CLK(clknet_leaf_19_clk),
    .D(_0018_),
    .RESET_B(net53),
    .Q(\outputs.div.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2673_ (.CLK(clknet_leaf_20_clk),
    .D(_0019_),
    .RESET_B(net51),
    .Q(\outputs.div.a[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2674_ (.CLK(clknet_leaf_19_clk),
    .D(_0020_),
    .RESET_B(net55),
    .Q(\outputs.div.a[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2675_ (.CLK(clknet_leaf_17_clk),
    .D(_0021_),
    .RESET_B(net55),
    .Q(\outputs.div.a[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2676_ (.CLK(clknet_leaf_17_clk),
    .D(_0022_),
    .RESET_B(net59),
    .Q(\outputs.div.a[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2677_ (.CLK(clknet_leaf_14_clk),
    .D(_0023_),
    .RESET_B(net57),
    .Q(\outputs.div.a[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2678_ (.CLK(clknet_leaf_14_clk),
    .D(_0024_),
    .RESET_B(net57),
    .Q(\outputs.div.a[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2679_ (.CLK(clknet_leaf_13_clk),
    .D(_0025_),
    .RESET_B(net57),
    .Q(\outputs.div.a[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2680_ (.CLK(clknet_leaf_12_clk),
    .D(_0026_),
    .RESET_B(net57),
    .Q(\outputs.div.a[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2681_ (.CLK(clknet_leaf_12_clk),
    .D(_0027_),
    .RESET_B(net51),
    .Q(\outputs.div.a[24] ));
 sky130_fd_sc_hd__dfrtp_2 _2682_ (.CLK(clknet_leaf_12_clk),
    .D(_0028_),
    .RESET_B(net51),
    .Q(\outputs.div.a[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2683_ (.CLK(clknet_leaf_17_clk),
    .D(_0029_),
    .RESET_B(net55),
    .Q(\outputs.div.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2684_ (.CLK(clknet_leaf_17_clk),
    .D(_0030_),
    .RESET_B(net55),
    .Q(\outputs.div.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2685_ (.CLK(clknet_leaf_17_clk),
    .D(_0031_),
    .RESET_B(net55),
    .Q(\outputs.div.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2686_ (.CLK(clknet_leaf_19_clk),
    .D(net234),
    .RESET_B(net53),
    .Q(\outputs.div.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2687_ (.CLK(clknet_leaf_19_clk),
    .D(net253),
    .RESET_B(net53),
    .Q(\outputs.div.q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2688_ (.CLK(clknet_leaf_19_clk),
    .D(_0034_),
    .RESET_B(net53),
    .Q(\outputs.div.q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2689_ (.CLK(clknet_leaf_19_clk),
    .D(net259),
    .RESET_B(net53),
    .Q(\outputs.div.q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2690_ (.CLK(clknet_leaf_19_clk),
    .D(net263),
    .RESET_B(net53),
    .Q(\outputs.div.q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2691_ (.CLK(clknet_leaf_12_clk),
    .D(_0037_),
    .RESET_B(net52),
    .Q(\outputs.div.q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2692_ (.CLK(clknet_leaf_12_clk),
    .D(_0038_),
    .RESET_B(net52),
    .Q(\outputs.div.q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2693_ (.CLK(clknet_leaf_12_clk),
    .D(_0039_),
    .RESET_B(net52),
    .Q(\outputs.div.q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2694_ (.CLK(clknet_leaf_12_clk),
    .D(net184),
    .RESET_B(net52),
    .Q(\outputs.div.q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2695_ (.CLK(clknet_leaf_13_clk),
    .D(net99),
    .RESET_B(net57),
    .Q(\outputs.div.q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2696_ (.CLK(clknet_leaf_13_clk),
    .D(net209),
    .RESET_B(net57),
    .Q(\outputs.div.q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2697_ (.CLK(clknet_leaf_9_clk),
    .D(net168),
    .RESET_B(net46),
    .Q(\outputs.div.q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2698_ (.CLK(clknet_leaf_9_clk),
    .D(net197),
    .RESET_B(net46),
    .Q(\outputs.div.q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2699_ (.CLK(clknet_leaf_7_clk),
    .D(net151),
    .RESET_B(net46),
    .Q(\outputs.div.q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2700_ (.CLK(clknet_leaf_6_clk),
    .D(net138),
    .RESET_B(net44),
    .Q(\outputs.div.q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2701_ (.CLK(clknet_leaf_7_clk),
    .D(net144),
    .RESET_B(net45),
    .Q(\outputs.div.q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2702_ (.CLK(clknet_leaf_7_clk),
    .D(net194),
    .RESET_B(net48),
    .Q(\outputs.div.q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2703_ (.CLK(clknet_leaf_7_clk),
    .D(_0049_),
    .RESET_B(net48),
    .Q(\outputs.div.q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2704_ (.CLK(clknet_leaf_8_clk),
    .D(net142),
    .RESET_B(net48),
    .Q(\outputs.div.q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2705_ (.CLK(clknet_leaf_8_clk),
    .D(net179),
    .RESET_B(net49),
    .Q(\outputs.div.q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2706_ (.CLK(clknet_leaf_8_clk),
    .D(_0052_),
    .RESET_B(net49),
    .Q(\outputs.div.q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2707_ (.CLK(clknet_leaf_13_clk),
    .D(net97),
    .RESET_B(net58),
    .Q(\outputs.div.q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _2708_ (.CLK(clknet_leaf_13_clk),
    .D(net205),
    .RESET_B(net57),
    .Q(\outputs.div.q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2709_ (.CLK(clknet_leaf_20_clk),
    .D(net217),
    .RESET_B(net53),
    .Q(\outputs.div.q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _2710_ (.CLK(clknet_leaf_13_clk),
    .D(_0056_),
    .RESET_B(net58),
    .Q(\outputs.div.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2711_ (.CLK(clknet_leaf_13_clk),
    .D(_0057_),
    .RESET_B(net57),
    .Q(\outputs.div.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2712_ (.CLK(clknet_leaf_13_clk),
    .D(_0058_),
    .RESET_B(net57),
    .Q(\outputs.div.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2713_ (.CLK(clknet_leaf_13_clk),
    .D(_0059_),
    .RESET_B(net57),
    .Q(\outputs.div.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2714_ (.CLK(clknet_leaf_12_clk),
    .D(_0060_),
    .RESET_B(net52),
    .Q(\outputs.div.count[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2715_ (.CLK(clknet_leaf_18_clk),
    .D(_0061_),
    .RESET_B(net55),
    .Q(\outputs.scaled_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2716_ (.CLK(clknet_leaf_18_clk),
    .D(_0062_),
    .RESET_B(net56),
    .Q(\outputs.scaled_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2717_ (.CLK(clknet_leaf_18_clk),
    .D(_0063_),
    .RESET_B(net54),
    .Q(\outputs.scaled_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2718_ (.CLK(clknet_leaf_18_clk),
    .D(_0064_),
    .RESET_B(net54),
    .Q(\outputs.scaled_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2719_ (.CLK(clknet_leaf_19_clk),
    .D(_0065_),
    .RESET_B(net54),
    .Q(\outputs.scaled_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2720_ (.CLK(clknet_leaf_23_clk),
    .D(_0066_),
    .RESET_B(net54),
    .Q(\outputs.scaled_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2721_ (.CLK(clknet_leaf_23_clk),
    .D(_0067_),
    .RESET_B(net36),
    .Q(\outputs.scaled_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2722_ (.CLK(clknet_leaf_22_clk),
    .D(_0068_),
    .RESET_B(net36),
    .Q(\outputs.scaled_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2723_ (.CLK(clknet_leaf_17_clk),
    .D(net165),
    .RESET_B(net56),
    .Q(\outputs.div.q_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2724_ (.CLK(clknet_leaf_18_clk),
    .D(net155),
    .RESET_B(net56),
    .Q(\outputs.div.q_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2725_ (.CLK(clknet_leaf_18_clk),
    .D(net161),
    .RESET_B(net54),
    .Q(\outputs.div.q_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2726_ (.CLK(clknet_leaf_18_clk),
    .D(net171),
    .RESET_B(net54),
    .Q(\outputs.div.q_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2727_ (.CLK(clknet_leaf_19_clk),
    .D(net175),
    .RESET_B(net54),
    .Q(\outputs.div.q_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2728_ (.CLK(clknet_leaf_19_clk),
    .D(net163),
    .RESET_B(net54),
    .Q(\outputs.div.q_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2729_ (.CLK(clknet_leaf_19_clk),
    .D(net199),
    .RESET_B(net53),
    .Q(\outputs.div.q_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2730_ (.CLK(clknet_leaf_19_clk),
    .D(net220),
    .RESET_B(net53),
    .Q(\outputs.div.q_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2731_ (.CLK(clknet_leaf_17_clk),
    .D(\outputs.div.next_div ),
    .RESET_B(net59),
    .Q(\outputs.div.div ));
 sky130_fd_sc_hd__dfrtp_1 _2732_ (.CLK(clknet_leaf_12_clk),
    .D(\outputs.div.next_start ),
    .RESET_B(net52),
    .Q(\outputs.div.start ));
 sky130_fd_sc_hd__dfrtp_1 _2733_ (.CLK(clknet_leaf_25_clk),
    .D(\outputs.output_gen.next_count[0] ),
    .RESET_B(net34),
    .Q(\outputs.output_gen.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2734_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.next_count[1] ),
    .RESET_B(net34),
    .Q(\outputs.output_gen.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2735_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.next_count[2] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2736_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.next_count[3] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2737_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.next_count[4] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2738_ (.CLK(clknet_leaf_24_clk),
    .D(\outputs.output_gen.next_count[5] ),
    .RESET_B(net35),
    .Q(\outputs.output_gen.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2739_ (.CLK(clknet_leaf_22_clk),
    .D(\outputs.output_gen.next_count[6] ),
    .RESET_B(net34),
    .Q(\outputs.output_gen.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2740_ (.CLK(clknet_leaf_22_clk),
    .D(\outputs.output_gen.next_count[7] ),
    .RESET_B(net34),
    .Q(\outputs.output_gen.count[7] ));
 sky130_fd_sc_hd__dfstp_2 _2741_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[0] ),
    .SET_B(net39),
    .Q(\outputs.sig_gen.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2742_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[1] ),
    .RESET_B(net39),
    .Q(\outputs.sig_gen.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2743_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[2] ),
    .RESET_B(net39),
    .Q(\outputs.sig_gen.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2744_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[3] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2745_ (.CLK(clknet_leaf_3_clk),
    .D(\outputs.sig_gen.next_count[4] ),
    .RESET_B(net39),
    .Q(\outputs.sig_gen.count[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2746_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[5] ),
    .RESET_B(net39),
    .Q(\outputs.sig_gen.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2747_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[6] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[6] ));
 sky130_fd_sc_hd__dfrtp_4 _2748_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[7] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2749_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[8] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2750_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[9] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2751_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[10] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2752_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[11] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2753_ (.CLK(clknet_leaf_4_clk),
    .D(\outputs.sig_gen.next_count[12] ),
    .RESET_B(net40),
    .Q(\outputs.sig_gen.count[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2754_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[13] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2755_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[14] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2756_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[15] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2757_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[16] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2758_ (.CLK(clknet_leaf_5_clk),
    .D(\outputs.sig_gen.next_count[17] ),
    .RESET_B(net44),
    .Q(\outputs.sig_gen.count[17] ));
 sky130_fd_sc_hd__dfrtp_4 _2759_ (.CLK(clknet_leaf_1_clk),
    .D(_0077_),
    .RESET_B(net28),
    .Q(\outputs.div.m[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2760_ (.CLK(clknet_leaf_31_clk),
    .D(_0078_),
    .RESET_B(net28),
    .Q(\outputs.div.m[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2761_ (.CLK(clknet_leaf_1_clk),
    .D(_0079_),
    .RESET_B(net27),
    .Q(\outputs.div.m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2762_ (.CLK(clknet_leaf_31_clk),
    .D(_0080_),
    .RESET_B(net28),
    .Q(\outputs.div.m[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2763_ (.CLK(clknet_leaf_32_clk),
    .D(_0081_),
    .RESET_B(net27),
    .Q(\outputs.div.m[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2764_ (.CLK(clknet_leaf_31_clk),
    .D(_0082_),
    .RESET_B(net33),
    .Q(\outputs.div.m[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2765_ (.CLK(clknet_leaf_30_clk),
    .D(_0083_),
    .RESET_B(net33),
    .Q(\outputs.div.m[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2766_ (.CLK(clknet_leaf_0_clk),
    .D(_0084_),
    .RESET_B(net27),
    .Q(\outputs.div.m[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2767_ (.CLK(clknet_leaf_31_clk),
    .D(_0085_),
    .RESET_B(net37),
    .Q(\outputs.div.m[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2768_ (.CLK(clknet_leaf_0_clk),
    .D(_0086_),
    .RESET_B(net26),
    .Q(\outputs.div.m[9] ));
 sky130_fd_sc_hd__dfrtp_4 _2769_ (.CLK(clknet_leaf_0_clk),
    .D(_0087_),
    .RESET_B(net25),
    .Q(\outputs.div.m[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2770_ (.CLK(clknet_leaf_0_clk),
    .D(_0088_),
    .RESET_B(net26),
    .Q(\outputs.div.m[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2771_ (.CLK(clknet_leaf_1_clk),
    .D(_0089_),
    .RESET_B(net28),
    .Q(\outputs.div.m[12] ));
 sky130_fd_sc_hd__dfrtp_4 _2772_ (.CLK(clknet_leaf_1_clk),
    .D(_0090_),
    .RESET_B(net28),
    .Q(\outputs.div.m[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2773_ (.CLK(clknet_leaf_11_clk),
    .D(_0091_),
    .RESET_B(net41),
    .Q(\outputs.div.m[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2774_ (.CLK(clknet_leaf_11_clk),
    .D(_0092_),
    .RESET_B(net51),
    .Q(\outputs.div.m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2775_ (.CLK(clknet_leaf_11_clk),
    .D(_0093_),
    .RESET_B(net51),
    .Q(\outputs.div.m[16] ));
 sky130_fd_sc_hd__dfrtp_4 _2776_ (.CLK(clknet_leaf_11_clk),
    .D(_0094_),
    .RESET_B(net51),
    .Q(\outputs.div.m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2777_ (.CLK(clknet_leaf_1_clk),
    .D(_0095_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2778_ (.CLK(clknet_leaf_31_clk),
    .D(_0096_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2779_ (.CLK(clknet_leaf_32_clk),
    .D(_0097_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2780_ (.CLK(clknet_leaf_32_clk),
    .D(_0098_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2781_ (.CLK(clknet_leaf_32_clk),
    .D(_0099_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2782_ (.CLK(clknet_leaf_31_clk),
    .D(_0100_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2783_ (.CLK(clknet_leaf_30_clk),
    .D(_0101_),
    .RESET_B(net33),
    .Q(\outputs.div.divisor[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2784_ (.CLK(clknet_leaf_0_clk),
    .D(_0102_),
    .RESET_B(net27),
    .Q(\outputs.div.divisor[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2785_ (.CLK(clknet_leaf_31_clk),
    .D(_0103_),
    .RESET_B(net29),
    .Q(\outputs.div.divisor[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2786_ (.CLK(clknet_leaf_0_clk),
    .D(_0104_),
    .RESET_B(net25),
    .Q(\outputs.div.divisor[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2787_ (.CLK(clknet_leaf_0_clk),
    .D(_0105_),
    .RESET_B(net25),
    .Q(\outputs.div.divisor[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2788_ (.CLK(clknet_leaf_36_clk),
    .D(_0106_),
    .RESET_B(net26),
    .Q(\outputs.div.divisor[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2789_ (.CLK(clknet_leaf_0_clk),
    .D(_0107_),
    .RESET_B(net26),
    .Q(\outputs.div.divisor[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2790_ (.CLK(clknet_leaf_1_clk),
    .D(_0108_),
    .RESET_B(net28),
    .Q(\outputs.div.divisor[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2791_ (.CLK(clknet_leaf_1_clk),
    .D(_0109_),
    .RESET_B(net28),
    .Q(\outputs.div.divisor[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2792_ (.CLK(clknet_leaf_31_clk),
    .D(_0110_),
    .RESET_B(net37),
    .Q(\outputs.div.divisor[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2793_ (.CLK(clknet_leaf_31_clk),
    .D(_0111_),
    .RESET_B(net37),
    .Q(\outputs.div.divisor[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2794_ (.CLK(clknet_leaf_11_clk),
    .D(_0112_),
    .RESET_B(net41),
    .Q(\outputs.div.divisor[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2795_ (.CLK(clknet_leaf_1_clk),
    .D(_0113_),
    .RESET_B(net28),
    .Q(\outputs.divider_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2796_ (.CLK(clknet_leaf_1_clk),
    .D(_0114_),
    .RESET_B(net29),
    .Q(\outputs.divider_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2797_ (.CLK(clknet_leaf_1_clk),
    .D(_0115_),
    .RESET_B(net28),
    .Q(\outputs.divider_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2798_ (.CLK(clknet_leaf_1_clk),
    .D(_0116_),
    .RESET_B(net29),
    .Q(\outputs.divider_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2799_ (.CLK(clknet_leaf_1_clk),
    .D(_0117_),
    .RESET_B(net29),
    .Q(\outputs.divider_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2800_ (.CLK(clknet_leaf_1_clk),
    .D(_0118_),
    .RESET_B(net28),
    .Q(\outputs.divider_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2801_ (.CLK(clknet_leaf_2_clk),
    .D(_0119_),
    .RESET_B(net41),
    .Q(\outputs.divider_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2802_ (.CLK(clknet_leaf_0_clk),
    .D(_0120_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2803_ (.CLK(clknet_leaf_1_clk),
    .D(_0121_),
    .RESET_B(net29),
    .Q(\outputs.divider_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2804_ (.CLK(clknet_leaf_0_clk),
    .D(_0122_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2805_ (.CLK(clknet_leaf_3_clk),
    .D(_0123_),
    .RESET_B(net39),
    .Q(\outputs.divider_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2806_ (.CLK(clknet_leaf_37_clk),
    .D(_0124_),
    .RESET_B(net26),
    .Q(\outputs.divider_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2807_ (.CLK(clknet_leaf_3_clk),
    .D(_0125_),
    .RESET_B(net39),
    .Q(\outputs.divider_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2808_ (.CLK(clknet_leaf_2_clk),
    .D(_0126_),
    .RESET_B(net41),
    .Q(\outputs.divider_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2809_ (.CLK(clknet_leaf_2_clk),
    .D(_0127_),
    .RESET_B(net41),
    .Q(\outputs.divider_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2810_ (.CLK(clknet_leaf_11_clk),
    .D(_0128_),
    .RESET_B(net42),
    .Q(\outputs.divider_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_2 _2811_ (.CLK(clknet_leaf_11_clk),
    .D(_0129_),
    .RESET_B(net52),
    .Q(\outputs.divider_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2812_ (.CLK(clknet_leaf_11_clk),
    .D(_0130_),
    .RESET_B(net42),
    .Q(\outputs.divider_buffer[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2813_ (.CLK(clknet_leaf_2_clk),
    .D(_0131_),
    .RESET_B(net41),
    .Q(\outputs.signal_buffer2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2814_ (.CLK(clknet_leaf_2_clk),
    .D(_0132_),
    .RESET_B(net41),
    .Q(\outputs.signal_buffer2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2815_ (.CLK(clknet_leaf_11_clk),
    .D(_0133_),
    .RESET_B(net42),
    .Q(\outputs.signal_buffer2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2816_ (.CLK(clknet_leaf_12_clk),
    .D(net109),
    .RESET_B(net42),
    .Q(\outputs.signal_buffer2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2817_ (.CLK(clknet_leaf_2_clk),
    .D(_0135_),
    .RESET_B(net42),
    .Q(\outputs.signal_buffer2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2818_ (.CLK(clknet_leaf_13_clk),
    .D(net124),
    .RESET_B(net46),
    .Q(\outputs.signal_buffer2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2819_ (.CLK(clknet_leaf_9_clk),
    .D(net102),
    .RESET_B(net46),
    .Q(\outputs.signal_buffer2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2820_ (.CLK(clknet_leaf_9_clk),
    .D(net121),
    .RESET_B(net46),
    .Q(\outputs.signal_buffer2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2821_ (.CLK(clknet_leaf_7_clk),
    .D(net130),
    .RESET_B(net44),
    .Q(\outputs.signal_buffer2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2822_ (.CLK(clknet_leaf_6_clk),
    .D(net117),
    .RESET_B(net45),
    .Q(\outputs.signal_buffer2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2823_ (.CLK(clknet_leaf_6_clk),
    .D(net132),
    .RESET_B(net45),
    .Q(\outputs.signal_buffer2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2824_ (.CLK(clknet_leaf_6_clk),
    .D(net113),
    .RESET_B(net45),
    .Q(\outputs.signal_buffer2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2825_ (.CLK(clknet_leaf_7_clk),
    .D(net104),
    .RESET_B(net48),
    .Q(\outputs.signal_buffer2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2826_ (.CLK(clknet_leaf_8_clk),
    .D(net115),
    .RESET_B(net48),
    .Q(\outputs.signal_buffer2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2827_ (.CLK(clknet_leaf_8_clk),
    .D(net107),
    .RESET_B(net49),
    .Q(\outputs.signal_buffer2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2828_ (.CLK(clknet_leaf_8_clk),
    .D(net136),
    .RESET_B(net49),
    .Q(\outputs.signal_buffer2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2829_ (.CLK(clknet_leaf_13_clk),
    .D(net127),
    .RESET_B(net49),
    .Q(\outputs.signal_buffer2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2830_ (.CLK(clknet_leaf_9_clk),
    .D(_0148_),
    .RESET_B(net46),
    .Q(\outputs.signal_buffer2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2831_ (.CLK(clknet_leaf_3_clk),
    .D(_0149_),
    .RESET_B(net39),
    .Q(\outputs.div.oscillator_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2832_ (.CLK(clknet_leaf_2_clk),
    .D(_0150_),
    .RESET_B(net41),
    .Q(\outputs.div.oscillator_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2833_ (.CLK(clknet_leaf_2_clk),
    .D(_0151_),
    .RESET_B(net41),
    .Q(\outputs.div.oscillator_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2834_ (.CLK(clknet_leaf_10_clk),
    .D(_0152_),
    .RESET_B(net42),
    .Q(\outputs.div.oscillator_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2835_ (.CLK(clknet_leaf_3_clk),
    .D(_0153_),
    .RESET_B(net39),
    .Q(\outputs.div.oscillator_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2836_ (.CLK(clknet_leaf_10_clk),
    .D(_0154_),
    .RESET_B(net46),
    .Q(\outputs.div.oscillator_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2837_ (.CLK(clknet_leaf_10_clk),
    .D(_0155_),
    .RESET_B(net42),
    .Q(\outputs.div.oscillator_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2838_ (.CLK(clknet_leaf_7_clk),
    .D(_0156_),
    .RESET_B(net46),
    .Q(\outputs.div.oscillator_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2839_ (.CLK(clknet_leaf_5_clk),
    .D(_0157_),
    .RESET_B(net44),
    .Q(\outputs.div.oscillator_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2840_ (.CLK(clknet_leaf_5_clk),
    .D(_0158_),
    .RESET_B(net44),
    .Q(\outputs.div.oscillator_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2841_ (.CLK(clknet_leaf_6_clk),
    .D(_0159_),
    .RESET_B(net45),
    .Q(\outputs.div.oscillator_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2842_ (.CLK(clknet_leaf_6_clk),
    .D(_0160_),
    .RESET_B(net50),
    .Q(\outputs.div.oscillator_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2843_ (.CLK(clknet_leaf_6_clk),
    .D(_0161_),
    .RESET_B(net50),
    .Q(\outputs.div.oscillator_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2844_ (.CLK(clknet_leaf_6_clk),
    .D(_0162_),
    .RESET_B(net50),
    .Q(\outputs.div.oscillator_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2845_ (.CLK(clknet_leaf_7_clk),
    .D(_0163_),
    .RESET_B(net48),
    .Q(\outputs.div.oscillator_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2846_ (.CLK(clknet_leaf_7_clk),
    .D(_0164_),
    .RESET_B(net48),
    .Q(\outputs.div.oscillator_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2847_ (.CLK(clknet_leaf_7_clk),
    .D(_0165_),
    .RESET_B(net48),
    .Q(\outputs.div.oscillator_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2848_ (.CLK(clknet_leaf_9_clk),
    .D(_0166_),
    .RESET_B(net46),
    .Q(\outputs.div.oscillator_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2849_ (.CLK(clknet_leaf_11_clk),
    .D(_0167_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2850_ (.CLK(clknet_leaf_2_clk),
    .D(_0168_),
    .RESET_B(net41),
    .Q(\outputs.shaper.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2851_ (.CLK(clknet_leaf_11_clk),
    .D(_0169_),
    .RESET_B(net42),
    .Q(\outputs.shaper.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2852_ (.CLK(clknet_leaf_11_clk),
    .D(_0170_),
    .RESET_B(net43),
    .Q(\outputs.shaper.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2853_ (.CLK(clknet_leaf_2_clk),
    .D(_0171_),
    .RESET_B(net43),
    .Q(\outputs.shaper.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2854_ (.CLK(clknet_leaf_13_clk),
    .D(_0172_),
    .RESET_B(net47),
    .Q(\outputs.shaper.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2855_ (.CLK(clknet_leaf_9_clk),
    .D(_0173_),
    .RESET_B(net47),
    .Q(\outputs.shaper.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2856_ (.CLK(clknet_leaf_9_clk),
    .D(_0174_),
    .RESET_B(net47),
    .Q(\outputs.shaper.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2857_ (.CLK(clknet_leaf_7_clk),
    .D(_0175_),
    .RESET_B(net45),
    .Q(\outputs.shaper.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2858_ (.CLK(clknet_leaf_5_clk),
    .D(_0176_),
    .RESET_B(net45),
    .Q(\outputs.shaper.count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2859_ (.CLK(clknet_leaf_6_clk),
    .D(_0177_),
    .RESET_B(net45),
    .Q(\outputs.shaper.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2860_ (.CLK(clknet_leaf_6_clk),
    .D(_0178_),
    .RESET_B(net50),
    .Q(\outputs.shaper.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2861_ (.CLK(clknet_leaf_7_clk),
    .D(_0179_),
    .RESET_B(net48),
    .Q(\outputs.shaper.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2862_ (.CLK(clknet_leaf_8_clk),
    .D(_0180_),
    .RESET_B(net48),
    .Q(\outputs.shaper.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2863_ (.CLK(clknet_leaf_8_clk),
    .D(_0181_),
    .RESET_B(net49),
    .Q(\outputs.shaper.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2864_ (.CLK(clknet_leaf_8_clk),
    .D(_0182_),
    .RESET_B(net47),
    .Q(\outputs.shaper.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2865_ (.CLK(clknet_leaf_8_clk),
    .D(_0183_),
    .RESET_B(net49),
    .Q(\outputs.shaper.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2866_ (.CLK(clknet_leaf_9_clk),
    .D(_0184_),
    .RESET_B(net47),
    .Q(\outputs.shaper.count[17] ));
 sky130_fd_sc_hd__dfstp_1 _2867_ (.CLK(clknet_leaf_34_clk),
    .D(_0185_),
    .SET_B(net22),
    .Q(\inputs.frequency_lut.rng[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2868_ (.CLK(clknet_leaf_34_clk),
    .D(_0186_),
    .RESET_B(net22),
    .Q(\inputs.frequency_lut.rng[1] ));
 sky130_fd_sc_hd__dfstp_2 _2869_ (.CLK(clknet_leaf_34_clk),
    .D(_0187_),
    .SET_B(net22),
    .Q(\inputs.frequency_lut.rng[2] ));
 sky130_fd_sc_hd__dfstp_1 _2870_ (.CLK(clknet_leaf_34_clk),
    .D(_0188_),
    .SET_B(net22),
    .Q(\inputs.frequency_lut.rng[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2871_ (.CLK(clknet_leaf_35_clk),
    .D(_0189_),
    .RESET_B(net23),
    .Q(\inputs.frequency_lut.rng[4] ));
 sky130_fd_sc_hd__dfstp_1 _2872_ (.CLK(clknet_leaf_35_clk),
    .D(_0190_),
    .SET_B(net23),
    .Q(\inputs.frequency_lut.rng[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2873_ (.CLK(clknet_leaf_24_clk),
    .D(net75),
    .RESET_B(net35),
    .Q(\outputs.pwm_output ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net38),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net38),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net29),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net38),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net38),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net37),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net36),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net19),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net43),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net43),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net19),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net50),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net50),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net50),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net19),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net62),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net62),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net56),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net62),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net62),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net62),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net61),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net19),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\inputs.keypad_synchronizer.half_sync[12] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\inputs.keypad_synchronizer.half_sync[2] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\outputs.div.q_out[5] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0074_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\outputs.div.q_out[0] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0069_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\outputs.div.a[14] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\outputs.div.q[13] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0043_),
    .X(net168));
 sky130_fd_sc_hd__buf_1 hold107 (.A(\inputs.random_update_clock.count[0] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\outputs.div.q_out[3] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0072_),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\inputs.keypad_synchronizer.half_sync[11] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\outputs.div.a[16] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\outputs.div.a[0] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\outputs.div.q_out[4] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0073_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\outputs.div.count[2] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\outputs.output_gen.count[7] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\outputs.div.q[21] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0051_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\outputs.div.a[10] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\outputs.div.a[12] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\inputs.random_note_generator.out[14] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\outputs.div.a[4] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\outputs.div.q[10] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0040_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\inputs.random_update_clock.count[14] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0971_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\outputs.div.q[19] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\outputs.div.a[23] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\outputs.div.q[9] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\outputs.div.a[6] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\outputs.div.a[5] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\outputs.output_gen.pwm_ff ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\outputs.div.a[8] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\outputs.div.q[18] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0048_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\outputs.div.q[8] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\outputs.div.q[14] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0044_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\outputs.div.q_out[6] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0075_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\inputs.random_update_clock.count[4] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\outputs.div.q[22] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\inputs.keypad_synchronizer.half_sync[8] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\inputs.random_update_clock.count[2] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0937_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\outputs.div.q[24] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0054_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\inputs.random_update_clock.count[16] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\outputs.sig_gen.count[17] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\outputs.div.q[12] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0042_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\outputs.div.a[1] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\outputs.div.a[7] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\inputs.random_note_generator.out[11] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\inputs.random_update_clock.count[3] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\inputs.random_update_clock.count[9] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\inputs.random_update_clock.count[1] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\outputs.div.a[24] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\outputs.div.q[26] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0055_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\inputs.random_update_clock.count[19] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\outputs.div.q_out[7] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0076_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\inputs.random_update_clock.count[11] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\inputs.keypad_synchronizer.half_sync[4] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\outputs.div.divisor[2] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\outputs.sample_rate.count[6] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\outputs.div.a[13] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\outputs.div.a[11] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\inputs.random_update_clock.count[20] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\inputs.random_update_clock.count[15] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\outputs.div.a[15] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\outputs.div.a[17] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\outputs.div.divisor[14] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\outputs.div.a[2] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\inputs.random_note_generator.out[3] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\outputs.div.divisor[16] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\outputs.div.q[2] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0032_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\outputs.div.count[4] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\outputs.div.a[20] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\inputs.random_update_clock.count[6] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\outputs.div.a[21] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\outputs.div.divisor[15] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\outputs.div.divisor[3] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\outputs.output_gen.count[2] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\inputs.random_note_generator.out[9] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0985_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\outputs.div.a[22] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\outputs.div.q[1] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\outputs.output_gen.count[4] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\outputs.div.count[1] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\inputs.random_update_clock.count[7] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\outputs.sig_gen.count[0] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\outputs.output_gen.count[5] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0989_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\outputs.div.a[19] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\inputs.random_note_generator.out[1] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\outputs.div.q[3] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0033_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\inputs.mode_edge.det_edge ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\inputs.wavetype_fsm.next_state[1] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\outputs.div.divisor[12] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\outputs.div.q[0] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\outputs.div.q[5] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0035_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\outputs.div.q[4] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\outputs.output_gen.count[3] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\inputs.keypad_synchronizer.half_sync[7] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\inputs.keypad_synchronizer.half_sync[1] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\outputs.div.q[6] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0036_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\outputs.div.oscillator_out[6] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\outputs.div.oscillator_out[0] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\outputs.div.a[18] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\outputs.div.oscillator_out[3] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\outputs.div.a[9] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\outputs.div.oscillator_out[8] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\outputs.div.oscillator_out[5] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\outputs.div.q[7] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\inputs.random_note_generator.out[6] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\outputs.div.oscillator_out[9] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\outputs.div.divisor[4] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\outputs.div.oscillator_out[4] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\outputs.div.oscillator_out[11] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\outputs.div.oscillator_out[10] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\outputs.div.oscillator_out[7] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\outputs.div.a[3] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\outputs.div.oscillator_out[2] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\outputs.div.divisor[1] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\outputs.div.oscillator_out[1] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\inputs.random_note_generator.out[4] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\outputs.div.divisor[7] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\outputs.div.divisor[0] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\outputs.div.oscillator_out[14] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\outputs.div.divisor[10] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\outputs.div.divisor[13] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\outputs.div.oscillator_out[15] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\outputs.div.divisor[11] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\outputs.div.oscillator_out[12] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\outputs.div.oscillator_out[17] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\outputs.div.oscillator_out[16] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\inputs.random_note_generator.out[2] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\outputs.div.divisor[8] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\inputs.random_update_clock.count[17] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\outputs.div.divisor[5] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\outputs.div.divisor[9] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\inputs.random_update_clock.count[5] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\outputs.div.m[6] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\outputs.shaper.count[11] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\outputs.shaper.count[12] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\outputs.shaper.count[1] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\outputs.shaper.count[8] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\inputs.keypad_synchronizer.half_sync[13] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\outputs.div.a[25] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\outputs.sample_rate.count[7] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\outputs.shaper.count[7] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\outputs.shaper.count[17] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\outputs.div.oscillator_out[13] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\outputs.sig_gen.count[5] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\outputs.scaled_buffer[7] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\outputs.divider_buffer[6] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\outputs.divider_buffer[14] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\outputs.divider_buffer[0] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\inputs.random_note_generator.out[0] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\outputs.divider_buffer[17] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\outputs.div.oscillator_out[15] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\outputs.div.oscillator_out[12] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\outputs.div.oscillator_out[2] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\inputs.random_note_generator.out[12] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\inputs.keypad_synchronizer.half_sync[16] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\inputs.keypad_synchronizer.half_sync[6] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\inputs.random_note_generator.out[13] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\inputs.keypad_synchronizer.half_sync[5] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\inputs.key_encoder.octave_key_up ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\inputs.random_note_generator.out[10] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\inputs.keypad_synchronizer.half_sync[0] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\inputs.keypad_synchronizer.half_sync[10] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\outputs.div.q[23] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0053_),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\outputs.div.q[11] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0041_),
    .X(net99));
 sky130_fd_sc_hd__buf_1 hold38 (.A(\outputs.output_gen.count[0] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\outputs.signal_buffer2[6] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\inputs.keypad_synchronizer.half_sync[3] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0137_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\outputs.signal_buffer2[12] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0143_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\outputs.signal_buffer2[4] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\outputs.signal_buffer2[14] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0145_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\outputs.signal_buffer2[3] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0134_),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\outputs.signal_buffer2[2] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\outputs.signal_buffer2[17] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\inputs.keypad_synchronizer.half_sync[14] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\outputs.signal_buffer2[11] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0142_),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\outputs.signal_buffer2[13] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0144_),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\outputs.signal_buffer2[9] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0140_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\inputs.random_update_clock.count[22] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\inputs.random_update_clock.next_count[22] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\outputs.signal_buffer2[7] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0138_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\inputs.random_note_generator.out[7] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\outputs.div.divisor[17] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\outputs.signal_buffer2[5] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0136_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\outputs.signal_buffer2[1] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\outputs.signal_buffer2[16] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0147_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\outputs.signal_buffer2[0] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\outputs.signal_buffer2[8] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0139_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\outputs.signal_buffer2[10] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\inputs.random_note_generator.out[5] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0141_),
    .X(net132));
 sky130_fd_sc_hd__buf_1 hold71 (.A(\outputs.sample_rate.count[0] ),
    .X(net133));
 sky130_fd_sc_hd__buf_1 hold72 (.A(\inputs.keypad_synchronizer.half_sync[15] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\outputs.signal_buffer2[15] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0146_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\outputs.div.q[16] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0046_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\outputs.sample_rate.count[5] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0999_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\outputs.div.q[20] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\inputs.random_note_generator.out[8] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0050_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\outputs.div.q[17] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0047_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\outputs.sample_rate.count[4] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\inputs.key_encoder.sync_keys[15] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\inputs.key_encoder.mode_key ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\outputs.sample_rate.count[1] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\inputs.mode_edge.ff_out ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\outputs.div.q[15] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0045_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\inputs.keypad_synchronizer.half_sync[9] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\outputs.sample_rate.count[3] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\outputs.output_gen.count[1] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\outputs.div.q_out[1] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0070_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\outputs.sample_rate.count[2] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0997_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\outputs.sample_rate.next_count[2] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\outputs.div.divisor[6] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\outputs.div.q_out[2] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0071_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(cs),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(gpio[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(gpio[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(gpio[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(gpio[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(gpio[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(gpio[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(gpio[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(gpio[8]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(gpio[9]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(nrst),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(gpio[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(gpio[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(gpio[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(gpio[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(gpio[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(gpio[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(gpio[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(gpio[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(pwm));
 sky130_fd_sc_hd__buf_4 wire21 (.A(_1155_),
    .X(net21));
endmodule

