VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pushing_pixels
  CLASS BLOCK ;
  FOREIGN pushing_pixels ;
  ORIGIN 0.000 0.000 ;
  SIZE 740.850 BY 751.570 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 737.470 747.570 737.750 751.570 ;
    END
  END clk
  PIN color[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END color[0]
  PIN color[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END color[10]
  PIN color[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END color[11]
  PIN color[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.290 747.570 193.570 751.570 ;
    END
  END color[12]
  PIN color[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 466.990 747.570 467.270 751.570 ;
    END
  END color[13]
  PIN color[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END color[14]
  PIN color[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 367.240 740.850 367.840 ;
    END
  END color[15]
  PIN color[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END color[16]
  PIN color[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 462.440 740.850 463.040 ;
    END
  END color[17]
  PIN color[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END color[18]
  PIN color[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END color[19]
  PIN color[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 557.150 747.570 557.430 751.570 ;
    END
  END color[1]
  PIN color[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 647.310 747.570 647.590 751.570 ;
    END
  END color[20]
  PIN color[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END color[21]
  PIN color[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 78.240 740.850 78.840 ;
    END
  END color[22]
  PIN color[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END color[23]
  PIN color[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END color[2]
  PIN color[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END color[3]
  PIN color[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END color[4]
  PIN color[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END color[5]
  PIN color[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 747.570 103.410 751.570 ;
    END
  END color[6]
  PIN color[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 173.440 740.850 174.040 ;
    END
  END color[7]
  PIN color[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END color[8]
  PIN color[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 557.640 740.850 558.240 ;
    END
  END color[9]
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 736.850 652.840 740.850 653.440 ;
    END
  END cs
  PIN is_mandelbrot
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 286.670 747.570 286.950 751.570 ;
    END
  END is_mandelbrot
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 376.830 747.570 377.110 751.570 ;
    END
  END nrst
  PIN spi_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END spi_clk
  PIN spi_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END spi_data
  PIN spi_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 747.570 13.250 751.570 ;
    END
  END spi_en
  PIN valid_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 736.850 272.040 740.850 272.640 ;
    END
  END valid_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 740.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 740.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 740.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 735.080 739.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 735.380 740.080 ;
      LAYER met2 ;
        RECT 0.100 747.290 12.690 747.570 ;
        RECT 13.530 747.290 102.850 747.570 ;
        RECT 103.690 747.290 193.010 747.570 ;
        RECT 193.850 747.290 286.390 747.570 ;
        RECT 287.230 747.290 376.550 747.570 ;
        RECT 377.390 747.290 466.710 747.570 ;
        RECT 467.550 747.290 556.870 747.570 ;
        RECT 557.710 747.290 647.030 747.570 ;
        RECT 647.870 747.290 737.190 747.570 ;
        RECT 0.100 4.280 737.750 747.290 ;
        RECT 0.650 4.000 89.970 4.280 ;
        RECT 90.810 4.000 180.130 4.280 ;
        RECT 180.970 4.000 270.290 4.280 ;
        RECT 271.130 4.000 360.450 4.280 ;
        RECT 361.290 4.000 450.610 4.280 ;
        RECT 451.450 4.000 543.990 4.280 ;
        RECT 544.830 4.000 634.150 4.280 ;
        RECT 634.990 4.000 724.310 4.280 ;
        RECT 725.150 4.000 737.750 4.280 ;
      LAYER met3 ;
        RECT 4.000 670.840 737.775 740.005 ;
        RECT 4.400 669.440 737.775 670.840 ;
        RECT 4.000 653.840 737.775 669.440 ;
        RECT 4.000 652.440 736.450 653.840 ;
        RECT 4.000 575.640 737.775 652.440 ;
        RECT 4.400 574.240 737.775 575.640 ;
        RECT 4.000 558.640 737.775 574.240 ;
        RECT 4.000 557.240 736.450 558.640 ;
        RECT 4.000 477.040 737.775 557.240 ;
        RECT 4.400 475.640 737.775 477.040 ;
        RECT 4.000 463.440 737.775 475.640 ;
        RECT 4.000 462.040 736.450 463.440 ;
        RECT 4.000 381.840 737.775 462.040 ;
        RECT 4.400 380.440 737.775 381.840 ;
        RECT 4.000 368.240 737.775 380.440 ;
        RECT 4.000 366.840 736.450 368.240 ;
        RECT 4.000 286.640 737.775 366.840 ;
        RECT 4.400 285.240 737.775 286.640 ;
        RECT 4.000 273.040 737.775 285.240 ;
        RECT 4.000 271.640 736.450 273.040 ;
        RECT 4.000 191.440 737.775 271.640 ;
        RECT 4.400 190.040 737.775 191.440 ;
        RECT 4.000 174.440 737.775 190.040 ;
        RECT 4.000 173.040 736.450 174.440 ;
        RECT 4.000 96.240 737.775 173.040 ;
        RECT 4.400 94.840 737.775 96.240 ;
        RECT 4.000 79.240 737.775 94.840 ;
        RECT 4.000 77.840 736.450 79.240 ;
        RECT 4.000 10.715 737.775 77.840 ;
      LAYER met4 ;
        RECT 19.190 13.095 20.640 738.985 ;
        RECT 23.040 13.095 97.440 738.985 ;
        RECT 99.840 13.095 174.240 738.985 ;
        RECT 176.640 13.095 251.040 738.985 ;
        RECT 253.440 13.095 327.840 738.985 ;
        RECT 330.240 13.095 404.640 738.985 ;
        RECT 407.040 13.095 481.440 738.985 ;
        RECT 483.840 13.095 558.240 738.985 ;
        RECT 560.640 13.095 635.040 738.985 ;
        RECT 637.440 13.095 711.840 738.985 ;
        RECT 714.240 13.095 732.450 738.985 ;
      LAYER met5 ;
        RECT 18.980 106.300 732.660 692.700 ;
  END
END pushing_pixels
END LIBRARY

