* NGSPICE file created from Eighty_Twos.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

.subckt Eighty_Twos clk cs gpi[0] gpi[10] gpi[11] gpi[12] gpi[13] gpi[14] gpi[15]
+ gpi[16] gpi[17] gpi[18] gpi[19] gpi[1] gpi[20] gpi[21] gpi[22] gpi[23] gpi[24] gpi[25]
+ gpi[26] gpi[27] gpi[28] gpi[29] gpi[2] gpi[30] gpi[31] gpi[32] gpi[33] gpi[3] gpi[4]
+ gpi[5] gpi[6] gpi[7] gpi[8] gpi[9] gpo[0] gpo[10] gpo[11] gpo[12] gpo[13] gpo[14]
+ gpo[15] gpo[16] gpo[17] gpo[18] gpo[19] gpo[1] gpo[20] gpo[21] gpo[22] gpo[23] gpo[24]
+ gpo[25] gpo[26] gpo[27] gpo[28] gpo[29] gpo[2] gpo[30] gpo[31] gpo[32] gpo[33] gpo[3]
+ gpo[4] gpo[5] gpo[6] gpo[7] gpo[8] gpo[9] nrst store_en vccd1 vssd1
X_2106_ _0630_ _0265_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o21ai_4
X_2037_ ByteBuffer.instr\[19\] net1 net4 _0261_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__and4_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2655_ net109 _0132_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.D\[6\] sky130_fd_sc_hd__dfrtp_2
X_1606_ ALU.flags_to_alu\[7\] _0788_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1399_ RegFile.H\[1\] _0707_ _0709_ RegFile.D\[1\] vssd1 vssd1 vccd1 vccd1 _0742_
+ sky130_fd_sc_hd__a22o_1
X_1537_ _0654_ _0876_ _0879_ _0828_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__a211o_2
X_1468_ RegFile.E\[2\] _0761_ _0771_ RegFile.B\[2\] vssd1 vssd1 vccd1 vccd1 _0811_
+ sky130_fd_sc_hd__a22o_1
X_2586_ ALU.immediate\[15\] _0585_ _0615_ _0540_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1322_ _0622_ _0618_ _0647_ _0619_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__o211a_1
X_2371_ ByteBuffer.counter\[0\] ByteBuffer.counter\[1\] _0659_ vssd1 vssd1 vccd1 vccd1
+ _0496_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2638_ net92 _0115_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[5\] sky130_fd_sc_hd__dfrtp_2
X_2569_ PC.i_mem_addr\[12\] _0597_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1940_ _1061_ _1172_ _1256_ _1056_ _0177_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ _1092_ _1160_ _1151_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2285_ RegFile.A\[5\] net1 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__and2_1
X_2354_ _0426_ ALU.immediate\[8\] _0407_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__mux2_1
X_1305_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0648_
+ sky130_fd_sc_hd__and2_4
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _0655_ _0267_ _0269_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1854_ _0645_ _0700_ _0661_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__a21o_1
X_1923_ _1093_ _1136_ _1213_ _1252_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1785_ _0806_ _1127_ _1074_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2406_ clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__buf_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2337_ _0479_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
X_2268_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__buf_6
X_2199_ _1221_ _1265_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2469__4 clknet_1_0__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__inv_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _0855_ _0844_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2122_ _0316_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
X_2053_ _1265_ _0262_ _0263_ net7 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a22o_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2424__25 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__inv_2
XFILLER_0_44_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1906_ _0655_ _1239_ _1246_ _0631_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a22o_1
X_1837_ _1158_ _1161_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1768_ _0868_ _0881_ _1108_ _1110_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a2bb2o_1
X_1699_ ByteBuffer.instr\[20\] _0645_ _0672_ _1041_ _0648_ vssd1 vssd1 vccd1 vccd1
+ _1042_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpo[6] sky130_fd_sc_hd__buf_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpo[27] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 gpo[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2671_ net125 _0148_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.B\[6\] sky130_fd_sc_hd__dfrtp_4
X_1622_ RegFile.A\[6\] vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1484_ ALU.flags_to_alu\[2\] _0704_ _0826_ _0629_ vssd1 vssd1 vccd1 vccd1 _0827_
+ sky130_fd_sc_hd__o211a_1
X_1553_ _0629_ _0892_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o21ai_4
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2105_ _0630_ _0286_ _1202_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a21oi_4
X_2036_ ByteBuffer.instr\[19\] _0261_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__nand2_4
XFILLER_0_27_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654_ net108 _0131_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.D\[5\] sky130_fd_sc_hd__dfrtp_2
X_1536_ ALU.flags_to_alu\[1\] _0711_ _0878_ _0654_ vssd1 vssd1 vccd1 vccd1 _0879_
+ sky130_fd_sc_hd__a211oi_1
X_1605_ RegFile.A\[7\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or3_1
X_2585_ PC.i_mem_addr\[15\] _0611_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1398_ RegFile.A\[1\] _0704_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__nor2_1
X_1467_ ALU.flags_to_alu\[2\] _0765_ _0763_ RegFile.H\[2\] vssd1 vssd1 vccd1 vccd1
+ _0810_ sky130_fd_sc_hd__a22o_1
X_2019_ _1184_ RegFile.B\[7\] _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2370_ _0495_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
X_1321_ _0626_ _0657_ _0635_ _0659_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o311a_4
XFILLER_0_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1519_ _0859_ _0860_ _0861_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__nor3_1
X_2637_ net91 _0114_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[4\] sky130_fd_sc_hd__dfrtp_2
X_2568_ _0601_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_2499_ _0543_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1870_ _1156_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__or2_1
X_2353_ _0486_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1304_ _0624_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__inv_2
X_2284_ _0450_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1999_ _1109_ _1123_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2445__45 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__inv_2
X_2460__59 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _0937_ _1210_ _1259_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o211a_1
X_1853_ _1194_ _1195_ _0626_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__a21oi_1
X_1784_ _0937_ _1056_ _1063_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__or3_2
X_2405_ clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__buf_1
X_2336_ _0732_ _0476_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and2_1
X_2267_ _0440_ _0655_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or2_1
X_2198_ _0377_ _0375_ _0376_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _0275_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
X_2121_ _0249_ RegFile.H\[0\] _0308_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1905_ _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ _0622_ _0624_ _0621_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1767_ _0908_ _0885_ _0896_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__a31o_1
X_1836_ _0960_ _1162_ _1170_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__a211o_1
X_2319_ PC.i_mem_addr\[11\] net46 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or2_1
X_2471__6 clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__inv_2
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpo[7] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 gpo[18] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpo[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1621_ RegFile.L\[6\] _0770_ _0763_ RegFile.H\[6\] net51 vssd1 vssd1 vccd1 vccd1
+ _0964_ sky130_fd_sc_hd__a221oi_1
X_2670_ net124 _0147_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.B\[5\] sky130_fd_sc_hd__dfrtp_2
X_1552_ _0893_ _0894_ _0693_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1483_ RegFile.C\[2\] _0705_ _0707_ RegFile.L\[2\] _0825_ vssd1 vssd1 vccd1 vccd1
+ _0826_ sky130_fd_sc_hd__a221o_1
X_2104_ _0306_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2035_ _0621_ _0628_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1819_ _1043_ _1160_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1535_ RegFile.C\[1\] _0705_ _0707_ RegFile.L\[1\] _0877_ vssd1 vssd1 vccd1 vccd1
+ _0878_ sky130_fd_sc_hd__a221o_1
X_2653_ net107 _0130_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.D\[4\] sky130_fd_sc_hd__dfrtp_2
X_2584_ _0614_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
X_1604_ _0780_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nand2_4
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1397_ RegFile.A\[1\] _0652_ _0676_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o211ai_4
X_1466_ RegFile.D\[2\] _0767_ _0807_ _0808_ net51 vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2018_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ _0645_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2636_ net90 _0113_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1518_ ALU.flags_to_alu\[1\] _0765_ _0761_ RegFile.E\[1\] vssd1 vssd1 vccd1 vccd1
+ _0861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1449_ _0648_ _0783_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__nor2_2
X_2567_ PC.i_mem_addr\[11\] _0600_ _0542_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__mux2_1
X_2498_ PC.i_mem_addr\[0\] _0541_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2283_ RegFile.A\[4\] net1 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__and2_1
X_1303_ _0619_ _0640_ _0644_ _0632_ _0645_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2352_ net128 _0438_ _0431_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2619_ net73 _0096_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1998_ _0885_ _0896_ _1172_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a21oi_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1852_ _0647_ _0656_ _0660_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__or3b_1
X_1921_ _1072_ _1172_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__o21ba_1
X_1783_ _1121_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2266_ ByteBuffer.instr\[19\] _0621_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or2_1
X_2335_ _0478_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_2404_ _0513_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2197_ _0375_ _0376_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 ALU.flags_to_alu\[4\] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2120_ _0315_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ RegFile.C\[5\] _0274_ _0270_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__mux2_1
X_1904_ _1011_ _1241_ _1243_ _1049_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1835_ _0908_ _1043_ _1165_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a31o_1
X_1697_ _0619_ _0620_ _0647_ ByteBuffer.instr\[19\] _1039_ vssd1 vssd1 vccd1 vccd1
+ _1040_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1766_ ALU.flags_to_alu\[0\] vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__inv_2
X_2318_ PC.i_mem_addr\[10\] net46 _0468_ _0445_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__o211a_1
X_2249_ _0420_ _0423_ net2 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a21o_1
X_2415__16 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__inv_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpo[19] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpo[29] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpo[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1620_ ALU.flags_to_alu\[6\] _0765_ _0767_ RegFile.D\[6\] _0962_ vssd1 vssd1 vccd1
+ vccd1 _0963_ sky130_fd_sc_hd__a221oi_1
X_1482_ RegFile.E\[2\] _0703_ _0699_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21a_1
X_1551_ ALU.flags_to_alu\[0\] _0711_ _0707_ RegFile.L\[0\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0894_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2103_ RegFile.E\[0\] _0284_ net48 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__mux2_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2034_ _0260_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1818_ _1092_ _1160_ _1151_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__o21a_1
X_1749_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2652_ net106 _0129_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.D\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1603_ _0629_ _0943_ _0944_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__o22a_2
X_1534_ RegFile.E\[1\] _0699_ _0706_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__and3_1
X_1465_ RegFile.L\[2\] _0638_ _0681_ _0762_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__and4_1
X_2583_ PC.i_mem_addr\[14\] _0613_ _0542_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1396_ RegFile.H\[1\] net54 _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a21o_1
X_2017_ _1188_ _1191_ _1201_ _1193_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2635_ net89 _0112_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1517_ RegFile.B\[1\] _0771_ _0763_ RegFile.H\[1\] vssd1 vssd1 vccd1 vccd1 _0860_
+ sky130_fd_sc_hd__a22o_1
X_1448_ ALU.flags_to_alu\[5\] _0788_ _0790_ _0711_ vssd1 vssd1 vccd1 vccd1 _0791_
+ sky130_fd_sc_hd__a22o_1
X_2566_ _0540_ _0598_ _0599_ _0585_ ALU.immediate\[11\] vssd1 vssd1 vccd1 vccd1 _0600_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2497_ _0659_ _0412_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__nor2_8
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1379_ RegFile.H\[3\] _0707_ _0709_ RegFile.D\[3\] vssd1 vssd1 vccd1 vccd1 _0722_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2282_ _0449_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
X_2351_ net130 _0416_ _0439_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__a21o_1
X_1302_ ByteBuffer.instr\[23\] vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__buf_8
XFILLER_0_51_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1997_ _1059_ _1140_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__and2_1
X_2618_ net72 _0095_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2549_ net47 _0583_ _0584_ _0585_ ALU.immediate\[8\] vssd1 vssd1 vccd1 vccd1 _0586_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2436__36 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__inv_2
X_1851_ _0622_ ByteBuffer.instr\[19\] _0624_ _0619_ vssd1 vssd1 vccd1 vccd1 _1194_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1920_ _0934_ _1255_ _1164_ _0855_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__a22o_1
X_2403_ _0418_ ALU.immediate\[7\] _0409_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__mux2_1
X_1782_ _1101_ _1120_ _1098_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o21ai_1
X_2334_ _0744_ _0476_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__and2_1
X_2265_ net141 _0413_ _0416_ _0627_ _0439_ vssd1 vssd1 vccd1 vccd1 FSM.next_state\[1\]
+ sky130_fd_sc_hd__a221o_1
X_2196_ _0855_ _1092_ _0347_ _0175_ _0182_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_47_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold11 ALU.flags_to_alu\[3\] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _1239_ _0262_ _0263_ net8 vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a22o_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1903_ _1241_ _1243_ _1011_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1765_ _0885_ _0896_ _0908_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a21o_1
X_1834_ _1172_ _1067_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__o21ai_1
X_1696_ ByteBuffer.instr\[20\] _0622_ _0624_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2317_ _0208_ net46 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2248_ net3 net5 vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__or2b_1
X_2179_ _0355_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 gpo[0] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpo[2] sky130_fd_sc_hd__clkbuf_4
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpo[1] sky130_fd_sc_hd__clkbuf_4
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpo[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1481_ RegFile.A\[2\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__or3_1
X_1550_ RegFile.C\[0\] _0705_ _0709_ RegFile.E\[0\] vssd1 vssd1 vccd1 vccd1 _0893_
+ sky130_fd_sc_hd__a22o_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2102_ _0305_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_2033_ _0249_ RegFile.B\[0\] _0252_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__mux2_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1748_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1817_ _1122_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__and2_2
X_1679_ _1020_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1602_ RegFile.L\[7\] net54 net53 RegFile.C\[7\] vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2651_ net105 _0128_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.D\[2\] sky130_fd_sc_hd__dfrtp_4
X_2582_ _0540_ _0611_ _0612_ _0585_ ALU.immediate\[14\] vssd1 vssd1 vccd1 vccd1 _0613_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1533_ _0870_ _0871_ net50 _0741_ _0789_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__a32o_1
X_1395_ RegFile.D\[1\] _0683_ net53 RegFile.B\[1\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0738_ sky130_fd_sc_hd__a221o_1
X_1464_ RegFile.C\[2\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2016_ _0250_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2634_ net88 _0111_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[1\] sky130_fd_sc_hd__dfrtp_2
X_1516_ RegFile.D\[1\] _0767_ _0857_ _0858_ net51 vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2565_ PC.i_mem_addr\[9\] PC.i_mem_addr\[10\] _0582_ PC.i_mem_addr\[11\] vssd1 vssd1
+ vccd1 vccd1 _0599_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1447_ RegFile.E\[5\] _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__or2_1
X_1378_ RegFile.A\[3\] _0652_ _0676_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o211a_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2496_ _0522_ _0455_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__mux2_1
X_2457__56 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__inv_2
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2281_ RegFile.A\[3\] net1 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__and2_1
X_1301_ _0618_ _0641_ _0635_ _0642_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__o221ai_4
X_2350_ net131 _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ _0231_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ net71 _0094_ net61 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[0\] sky130_fd_sc_hd__dfrtp_4
X_2548_ _0534_ _0537_ _0520_ _0539_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__o211a_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ ByteBuffer.instr\[19\] _0639_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ _0700_ _1185_ _1187_ ByteBuffer.instr\[21\] _0645_ vssd1 vssd1 vccd1 vccd1
+ _1193_ sky130_fd_sc_hd__a221o_2
X_1781_ _1043_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2333_ _0477_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_2402_ _0512_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2195_ _0373_ _0374_ _0361_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2264_ _0432_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ _1139_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__xor2_1
Xhold12 ALU.flags_to_alu\[5\] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1902_ _1000_ _1020_ _1242_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1764_ _0868_ _0881_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nand2_1
X_1833_ _1174_ _1175_ _0947_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__mux2_1
X_1695_ _0715_ _1026_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__o21a_1
X_2316_ _0467_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2247_ net7 _0417_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and2_1
X_2178_ _0357_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__xnor2_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpo[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 store_en sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 gpo[10] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 gpo[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1480_ _0819_ _0821_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__or3_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2101_ RegFile.E\[1\] _0282_ net48 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__mux2_1
X_2032_ _0259_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2420__21 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__inv_2
X_1678_ _1014_ _1018_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__nand2_1
X_1747_ _1037_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1816_ ByteBuffer.instr\[21\] _0645_ _1045_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ net104 _0127_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.D\[1\] sky130_fd_sc_hd__dfrtp_2
X_1532_ RegFile.L\[1\] _0817_ _0872_ _0873_ _0874_ vssd1 vssd1 vccd1 vccd1 _0875_
+ sky130_fd_sc_hd__a2111oi_1
X_1601_ ALU.flags_to_alu\[7\] _0687_ _0683_ RegFile.E\[7\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0944_ sky130_fd_sc_hd__a221o_1
X_2581_ PC.i_mem_addr\[14\] _0606_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1394_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__inv_2
X_1463_ _0804_ _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2015_ RegFile.A\[0\] _0249_ _1203_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2702_ clknet_2_0__leaf_clk ByteBuffer.next_counter\[1\] net57 vssd1 vssd1 vccd1
+ vccd1 ByteBuffer.counter\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1515_ RegFile.C\[1\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2633_ net87 _0110_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.H\[0\] sky130_fd_sc_hd__dfrtp_2
X_2564_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__inv_2
X_2495_ _0534_ _0537_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1377_ RegFile.H\[3\] net54 _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a21o_1
X_1446_ _0678_ _0785_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nand2_4
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1300_ ByteBuffer.instr\[21\] _0624_ ByteBuffer.instr\[17\] ByteBuffer.instr\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or4bb_1
X_2280_ _0448_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ RegFile.A\[1\] _0230_ _1203_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2616_ clknet_2_3__leaf_clk _0093_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1429_ _0638_ _0646_ _0650_ _0760_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__nor4_1
X_2478_ _0678_ _0636_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nor2_1
X_2547_ PC.i_mem_addr\[6\] PC.i_mem_addr\[7\] _0567_ PC.i_mem_addr\[8\] vssd1 vssd1
+ vccd1 vccd1 _0584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _1047_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_2
XFILLER_0_21_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2332_ _0752_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2401_ _0429_ ALU.immediate\[6\] _0409_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2194_ _0361_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ net9 _0418_ _0433_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2427__27 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__inv_2
XFILLER_0_30_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1978_ _1108_ _1110_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__nand2_1
Xhold13 ALU.flags_to_alu\[6\] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlygate4sd3_1
X_2441__41 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__inv_2
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1901_ _1151_ _1021_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1832_ _1043_ _1173_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_2
X_1694_ _1034_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__nand2_1
X_1763_ _0816_ _0831_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2315_ _0445_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__and2_1
X_2246_ net8 _0417_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2177_ _0908_ _0232_ _1092_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpo[21] sky130_fd_sc_hd__buf_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 gpo[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 gpo[11] sky130_fd_sc_hd__clkbuf_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2100_ _0304_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2031_ _0230_ RegFile.B\[1\] _0252_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1815_ _0960_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1677_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1746_ _0718_ _1088_ _0716_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2229_ net132 _0659_ vssd1 vssd1 vccd1 vccd1 ByteBuffer.next_counter\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1600_ _0939_ _0941_ _0942_ _0774_ RegFile.A\[7\] vssd1 vssd1 vccd1 vccd1 _0943_
+ sky130_fd_sc_hd__o32a_1
X_1531_ RegFile.E\[1\] _0789_ _0699_ _0703_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2580_ PC.i_mem_addr\[14\] _0606_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1462_ _0781_ _0803_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1393_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__and2_1
X_2014_ _0655_ _0243_ _0248_ _0631_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1729_ _0780_ _0921_ _0929_ _0933_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand4_2
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2632_ net86 _0109_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.L\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ clknet_2_1__leaf_clk ByteBuffer.next_counter\[0\] net61 vssd1 vssd1 vccd1
+ vccd1 ByteBuffer.counter\[0\] sky130_fd_sc_hd__dfrtp_1
X_1514_ RegFile.L\[1\] _0638_ _0681_ _0762_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1445_ _0783_ _0708_ _0703_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__and3_2
X_2563_ PC.i_mem_addr\[10\] PC.i_mem_addr\[11\] _0588_ vssd1 vssd1 vccd1 vccd1 _0597_
+ sky130_fd_sc_hd__and3_1
X_2494_ _0525_ _0527_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or3_2
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1376_ RegFile.D\[3\] _0683_ net53 RegFile.B\[3\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2448__47 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__inv_2
Xfanout60 net61 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2462__61 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XFILLER_0_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1994_ _0655_ _0224_ _0229_ _0631_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2615_ clknet_2_0__leaf_clk _0092_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1428_ net56 _0650_ _0766_ _0638_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o211a_4
X_2546_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__inv_2
X_2477_ ALU.immediate\[0\] _0520_ _0521_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__a21o_1
X_1359_ ByteBuffer.instr\[21\] _0667_ _0668_ _0696_ vssd1 vssd1 vccd1 vccd1 _0702_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2400_ _0511_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2331_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2262_ net2 _0434_ _0435_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2193_ _0365_ _0366_ _0372_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1977_ _1141_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2529_ _0567_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nor2_1
Xhold14 ByteDecoder.state\[1\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1900_ _1022_ _1085_ _1240_ _1151_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__a211o_1
X_1831_ _1151_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__nand2_1
X_1693_ _1035_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__inv_2
X_1762_ _0937_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__or2_1
X_2314_ PC.i_mem_addr\[9\] _0229_ net46 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__mux2_1
X_2245_ net5 net3 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or2b_1
X_2176_ _0781_ _1049_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a21oi_1
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 gpo[32] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpo[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 gpo[12] sky130_fd_sc_hd__clkbuf_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2030_ _0258_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ _1011_ _1022_ _1085_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a31o_1
X_1814_ _1069_ _1153_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a21o_1
X_1676_ _1014_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2228_ _0406_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
X_2159_ _1201_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2411__12 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__inv_2
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1530_ RegFile.D\[1\] _0785_ _0708_ _0703_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1392_ _0729_ _0733_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__or2_1
X_1461_ _0781_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2013_ _0246_ _0247_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__nor2_2
X_1728_ _0782_ _0802_ _0781_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__a21o_1
X_1659_ RegFile.H\[5\] net54 _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__a21o_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2631_ net85 _0108_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.L\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2562_ _0596_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_2700_ clknet_2_1__leaf_clk FSM.next_state\[1\] net61 vssd1 vssd1 vccd1 vccd1 ByteDecoder.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1444_ RegFile.H\[5\] _0784_ _0786_ RegFile.D\[5\] vssd1 vssd1 vccd1 vccd1 _0787_
+ sky130_fd_sc_hd__a22o_1
X_1375_ _0716_ _0717_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nor2_2
X_2493_ ByteBuffer.instr\[21\] _0621_ _0648_ _0647_ vssd1 vssd1 vccd1 vccd1 _0538_
+ sky130_fd_sc_hd__o211a_1
X_1513_ _0844_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout61 net11 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2545_ PC.i_mem_addr\[7\] PC.i_mem_addr\[8\] _0573_ vssd1 vssd1 vccd1 vccd1 _0582_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2614_ clknet_2_1__leaf_clk _0091_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1427_ _0638_ _0681_ _0762_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__and3_2
X_1358_ _0645_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__nand2_1
X_2476_ _0903_ _0906_ _0519_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__and3_1
X_1289_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0632_
+ sky130_fd_sc_hd__nand2b_4
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2330_ net1 net4 net46 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__nand3_1
X_2192_ _0365_ _0366_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2261_ net3 _0417_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1976_ _1139_ _1059_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2528_ PC.i_mem_addr\[4\] _0556_ PC.i_mem_addr\[5\] vssd1 vssd1 vccd1 vccd1 _0568_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2432__32 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__inv_2
X_1761_ _0855_ _0844_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__and2b_1
X_1830_ ByteBuffer.instr\[21\] _0670_ _1044_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__and3_1
X_1692_ _1029_ _1033_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__nor2_1
X_2313_ _0465_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2244_ net9 _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__nand2_1
X_2175_ _1043_ _1229_ _1235_ _1092_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1959_ _1062_ _1172_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__nor2_1
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 gpo[33] sky130_fd_sc_hd__buf_2
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 gpo[13] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpo[23] sky130_fd_sc_hd__clkbuf_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1008_ _1086_ _1010_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a21oi_1
X_1813_ _0983_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ ALU.immediate\[12\] _0675_ _0693_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a22o_1
X_2089_ RegFile.E\[7\] _0264_ _0298_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__mux2_1
X_2227_ ALU.flags_to_alu\[0\] _0405_ _0335_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__mux2_1
X_2158_ _1182_ _0339_ _0340_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__or4_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1391_ _0729_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand2_1
X_1460_ _0782_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2012_ _0756_ _0244_ _0245_ _1049_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1658_ RegFile.D\[5\] _0683_ net53 RegFile.B\[5\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _1001_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1727_ _1069_ _0982_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ RegFile.E\[4\] _0699_ _0706_ _0654_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__a31o_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ net84 _0107_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.L\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2561_ PC.i_mem_addr\[10\] _0595_ _0542_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__mux2_1
X_2492_ _0535_ _0536_ _0388_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__mux2_1
X_1512_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__clkbuf_4
X_1443_ _0785_ _0708_ _0703_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__and3_2
X_1374_ _0690_ _0714_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_8
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1992_ _1054_ _0226_ _0227_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2544_ _0581_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2613_ clknet_2_0__leaf_clk _0090_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2475_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__inv_2
X_1426_ ALU.flags_to_alu\[5\] _0765_ _0767_ RegFile.D\[5\] _0768_ vssd1 vssd1 vccd1
+ vccd1 _0769_ sky130_fd_sc_hd__a221o_1
X_1288_ _0618_ _0621_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__o21a_2
X_1357_ ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2453__52 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__inv_2
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2191_ _0208_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__xnor2_1
X_2260_ net5 _0417_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1975_ _0211_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1409_ RegFile.A\[0\] _0704_ _0751_ _0630_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2527_ PC.i_mem_addr\[4\] PC.i_mem_addr\[5\] _0556_ vssd1 vssd1 vccd1 vccd1 _0567_
+ sky130_fd_sc_hd__and3_1
X_2418__19 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__inv_2
X_2389_ _0426_ ALU.immediate\[0\] _0409_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1691_ _1029_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nand2_1
X_1760_ _1101_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__nor2_1
X_2312_ _0445_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2243_ net10 _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__and2_2
X_2174_ _0349_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__xnor2_1
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 gpo[14] sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpo[24] sky130_fd_sc_hd__buf_2
XFILLER_0_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ _0912_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 gpo[3] sky130_fd_sc_hd__clkbuf_4
X_1889_ _1069_ _1165_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1674_ RegFile.A\[4\] _0704_ _1016_ _0630_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__o211a_1
X_1743_ _1014_ _1018_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1812_ _1132_ _1154_ _0804_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o21ba_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _0284_ _0404_ _1201_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__mux2_1
X_2088_ _1192_ _0655_ _0288_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__a21oi_4
X_2157_ _1221_ _1239_ _1265_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1390_ ALU.immediate\[10\] _0675_ _0693_ _0732_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2011_ _0244_ _0245_ _0756_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1588_ RegFile.C\[4\] _0705_ _0707_ RegFile.L\[4\] vssd1 vssd1 vccd1 vccd1 _0931_
+ sky130_fd_sc_hd__a22o_1
X_1657_ _0726_ _0997_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__a21oi_1
X_1726_ _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ ALU.flags_to_alu\[2\] _0389_ _0335_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__mux2_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2560_ _0540_ _0593_ _0594_ _0585_ ALU.immediate\[10\] vssd1 vssd1 vccd1 vccd1 _0595_
+ sky130_fd_sc_hd__a32o_1
X_1442_ _0645_ _0647_ _0642_ _0672_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__a22o_2
X_2491_ _0636_ _0525_ _0697_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and3b_1
X_1511_ _0780_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1373_ _0690_ _0714_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1709_ _0726_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__inv_2
X_2689_ clknet_2_2__leaf_clk _0166_ net58 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout63 net11 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_6
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2439__39 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__inv_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1991_ _1054_ _0226_ _1049_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a21oi_1
X_2612_ clknet_2_1__leaf_clk _0089_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1425_ RegFile.C\[5\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__and4_1
X_2543_ PC.i_mem_addr\[7\] _0580_ _0542_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__mux2_1
X_2474_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1356_ _0694_ _0698_ _0648_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__a21o_4
X_1287_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__buf_8
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2190_ _0367_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1974_ RegFile.A\[2\] _0210_ _1203_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1408_ RegFile.B\[0\] _0705_ _0750_ _0711_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2526_ ALU.immediate\[5\] _0565_ _0519_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__mux2_1
X_2388_ _0505_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
X_1339_ _0638_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1690_ ALU.immediate\[15\] _0675_ _0693_ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2242_ net4 net1 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__and2b_2
XFILLER_0_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2311_ PC.i_mem_addr\[8\] _0248_ net46 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__mux2_1
X_2173_ _0351_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__xnor2_1
X_1957_ _0911_ _0882_ _0910_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 gpo[15] sky130_fd_sc_hd__clkbuf_4
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpo[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2509_ _0550_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__nor2_1
X_1888_ _1132_ _1154_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1811_ _0935_ _0938_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nor2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1673_ RegFile.B\[4\] _0705_ _1015_ _0711_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__a211o_1
X_1742_ _1052_ _0736_ _1082_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _0393_ _0399_ _0403_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2087_ _0297_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_2156_ _0183_ _0204_ _0224_ _0243_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ net49 _0990_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1725_ _0780_ _0969_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__and2_1
X_1587_ ALU.flags_to_alu\[4\] _0699_ _0703_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__and3_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ _0998_ _0725_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0325_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_2208_ _0280_ _0388_ _1201_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2467__2 clknet_1_0__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1510_ _0629_ _0850_ _0851_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1441_ _0783_ _0708_ _0706_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__and3_4
X_2490_ _0678_ _0526_ _0531_ _0523_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1372_ _0691_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1708_ _1037_ _0715_ _1026_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2688_ clknet_2_2__leaf_clk _0165_ net58 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ _0693_ _0978_ _0981_ _0675_ ALU.immediate\[6\] vssd1 vssd1 vccd1 vccd1 _0982_
+ sky130_fd_sc_hd__a32o_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1990_ _0225_ _1080_ net49 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2542_ _0578_ _0579_ net47 vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2611_ clknet_2_1__leaf_clk _0088_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1424_ net56 _0650_ _0766_ _0684_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o211a_2
X_1355_ _0695_ _0696_ _0672_ _0642_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__o2111ai_4
X_2473_ _0659_ _0669_ _0648_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__and3_1
X_2407__8 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_2
X_1286_ _0623_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__nor2_8
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1973_ _0655_ _0204_ _0209_ _0631_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a22o_1
X_2525_ _0630_ _0775_ _0778_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1407_ RegFile.H\[0\] _0707_ _0709_ RegFile.D\[0\] vssd1 vssd1 vccd1 vccd1 _0750_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1338_ _0619_ _0640_ _0644_ _0632_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__a22o_4
X_2387_ _0418_ _0645_ _0497_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2310_ _1182_ _0442_ _0463_ _0445_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__o211a_1
X_2241_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] vssd1 vssd1 vccd1 vccd1 _0416_
+ sky130_fd_sc_hd__or2_1
X_2172_ _0197_ _1092_ _1093_ _0212_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__o221a_1
X_2423__24 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__inv_2
X_1956_ _1057_ _1107_ _1111_ _1236_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1887_ _1134_ _1227_ _1207_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 gpo[16] sky130_fd_sc_hd__clkbuf_4
X_2508_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] PC.i_mem_addr\[2\] vssd1 vssd1 vccd1
+ vccd1 _0551_ sky130_fd_sc_hd__and3_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1741_ _0721_ _0725_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1810_ _0982_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__inv_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1672_ RegFile.H\[4\] _0707_ _0709_ RegFile.D\[4\] vssd1 vssd1 vccd1 vccd1 _1015_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2224_ _0347_ _1038_ _0401_ _0402_ _0630_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__o311a_1
X_2155_ _0229_ _0248_ _0630_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2086_ RegFile.D\[0\] _0249_ _0289_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1939_ _0922_ _1253_ _0176_ _1093_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1724_ _1066_ _0959_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _0923_ _0928_ _0629_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a21o_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _0721_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _0284_ RegFile.L\[0\] _0317_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__mux2_1
X_2069_ _0655_ _0286_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__and2_2
X_2207_ _0655_ _0378_ _0379_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1371_ ALU.immediate\[14\] _0675_ _0693_ _0713_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a22o_1
X_1440_ _0672_ _0642_ _0624_ _0670_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1707_ net49 _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__nor2_2
X_1638_ _0655_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__or2_1
X_2687_ clknet_2_2__leaf_clk _0164_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1569_ _0882_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__a21oi_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2541_ PC.i_mem_addr\[7\] _0573_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2610_ clknet_2_1__leaf_clk _0087_ net58 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1423_ _0670_ _0757_ _0759_ _0650_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__a31o_1
X_1354_ ByteBuffer.instr\[20\] vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__inv_2
X_1285_ _0624_ _0626_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__or3_4
XFILLER_0_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2444__44 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__inv_2
XFILLER_0_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2524_ _0564_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
X_1406_ RegFile.A\[0\] _0652_ _0676_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__o211a_1
X_1337_ _0677_ _0679_ _0638_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a21oi_4
X_2386_ _0504_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2240_ ByteDecoder.state\[1\] _0413_ _0414_ net128 _0415_ vssd1 vssd1 vccd1 vccd1
+ FSM.next_state\[0\] sky130_fd_sc_hd__a221o_1
X_2171_ _1050_ _0218_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _1107_ _1111_ _1057_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1886_ _1136_ _1146_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2507_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] PC.i_mem_addr\[2\] vssd1 vssd1 vccd1
+ vccd1 _0550_ sky130_fd_sc_hd__a21oi_1
X_2369_ _0418_ ALU.immediate\[15\] _0407_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__mux2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1671_ RegFile.A\[4\] _0652_ _0676_ _1013_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1740_ _0721_ _0725_ _0729_ _0733_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2085_ _0296_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
X_2154_ _1094_ _0187_ _0338_ _0630_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__o31a_1
X_2223_ _1034_ _1089_ _1035_ _1093_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1938_ _0855_ _1175_ _1214_ _0816_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1869_ _0983_ _1155_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1654_ _0737_ _0746_ _0994_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a31o_1
X_1723_ _0780_ _0946_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ RegFile.L\[4\] _0817_ _0924_ _0925_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_
+ sky130_fd_sc_hd__a2111o_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _0655_ _0386_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2137_ _0324_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
X_2068_ _0266_ _1191_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1370_ RegFile.A\[6\] _0704_ _0712_ _0630_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465__64 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
X_1637_ ALU.flags_to_alu\[6\] _0711_ _0709_ RegFile.E\[6\] _0979_ vssd1 vssd1 vccd1
+ vccd1 _0980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2686_ clknet_2_2__leaf_clk _0163_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1706_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nand2_8
X_1499_ ALU.flags_to_alu\[3\] _0704_ _0841_ _0629_ vssd1 vssd1 vccd1 vccd1 _0842_
+ sky130_fd_sc_hd__o211a_1
X_1568_ _0816_ _0831_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__xnor2_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0517_ clknet_0__0517_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0517_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1422_ net56 _0650_ _0762_ _0684_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o211a_2
X_2540_ ALU.immediate\[7\] _0946_ _0519_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__mux2_1
X_1353_ _0619_ _0624_ _0622_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__or3b_4
X_1284_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] vssd1 vssd1 vccd1 vccd1 _0627_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2669_ net123 _0146_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.B\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1971_ _0736_ _0206_ _0207_ _1049_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a211o_2
X_1405_ RegFile.B\[0\] net53 _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2385_ _0429_ ByteBuffer.instr\[22\] _0497_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__mux2_1
X_2523_ PC.i_mem_addr\[4\] _0563_ _0542_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__mux2_1
X_1336_ _0622_ _0624_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__or3_4
Xinput1 cs vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2170_ _1050_ _0195_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a21oi_1
X_1954_ _1143_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__nor2_1
X_1885_ _1226_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2506_ ALU.immediate\[2\] _0815_ _0519_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__mux2_1
X_2368_ _0494_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__clkbuf_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ ByteBuffer.instr\[22\] _0618_ _0660_ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2299_ PC.i_mem_addr\[2\] net46 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or2_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2414__15 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__inv_2
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap52 _0772_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1670_ RegFile.H\[4\] net54 _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__a21o_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _0400_ _1033_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__nor2_1
X_2084_ RegFile.D\[1\] _0230_ _0289_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_1
X_2153_ _1224_ _1246_ _1268_ _0209_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1937_ _1113_ _0174_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1799_ _1139_ _1141_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__nand2_1
X_1868_ _1043_ _1160_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1584_ ALU.flags_to_alu\[4\] _0788_ _0926_ _0711_ vssd1 vssd1 vccd1 vccd1 _0927_
+ sky130_fd_sc_hd__a22o_1
X_1653_ _0995_ _0733_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _0806_ _0937_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nor2_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0183_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2136_ _0282_ RegFile.L\[1\] _0317_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_1
X_2067_ _0285_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1705_ _0645_ _1044_ _1045_ ByteBuffer.instr\[19\] vssd1 vssd1 vccd1 vccd1 _1048_
+ sky130_fd_sc_hd__o211ai_4
X_1636_ RegFile.C\[6\] _0705_ _0707_ RegFile.L\[6\] vssd1 vssd1 vccd1 vccd1 _0979_
+ sky130_fd_sc_hd__a22o_1
X_1567_ _0883_ _0884_ _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a21o_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2685_ clknet_2_0__leaf_clk _0162_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2119_ _0230_ RegFile.H\[1\] _0308_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1498_ RegFile.C\[3\] _0705_ _0707_ RegFile.L\[3\] _0840_ vssd1 vssd1 vccd1 vccd1
+ _0841_ sky130_fd_sc_hd__a221o_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__0516_ clknet_0__0516_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0516_
+ sky130_fd_sc_hd__clkbuf_16
X_1421_ RegFile.E\[5\] _0761_ _0763_ RegFile.H\[5\] vssd1 vssd1 vccd1 vccd1 _0764_
+ sky130_fd_sc_hd__a22o_1
X_1352_ ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__inv_2
X_1283_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2668_ net122 _0145_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.B\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1619_ RegFile.C\[6\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2599_ clknet_2_3__leaf_clk _0076_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2435__35 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__inv_2
X_1970_ _0736_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2450__49 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__inv_2
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2522_ _0561_ _0562_ net47 vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__mux2_1
X_1404_ RegFile.H\[0\] _0680_ _0683_ RegFile.D\[0\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0747_ sky130_fd_sc_hd__a221o_1
X_1335_ _0645_ ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_8
X_2384_ _0503_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 gpi[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1884_ RegFile.A\[6\] _1225_ _1203_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1953_ _1137_ _1142_ _1207_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__a21bo_1
X_2505_ _0548_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ _0619_ _0622_ _0624_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2298_ _0224_ _0442_ _0457_ _0445_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__o211a_1
X_2367_ _0429_ ALU.immediate\[14\] _0407_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap53 _0685_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_4
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _0335_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_2221_ _1029_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
X_2083_ _0295_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1936_ _0832_ _0912_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1867_ _1148_ _1207_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1798_ ALU.flags_to_alu\[0\] _1059_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1721_ _1056_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1583_ RegFile.E\[4\] _0789_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or2_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _0729_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__inv_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0323_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _0383_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2066_ RegFile.C\[0\] _0284_ _0270_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1919_ _0781_ _1253_ _1256_ _0922_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2684_ clknet_2_0__leaf_clk _0161_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1704_ _0670_ _1044_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__a21oi_4
X_1635_ _0971_ _0977_ _0629_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__a21o_1
X_1497_ RegFile.E\[3\] _0703_ _0699_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1566_ _0885_ _0896_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__a21oi_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2456__55 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__inv_2
X_2049_ _0273_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2118_ _0314_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout57 net58 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_6
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__0515_ clknet_0__0515_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0515_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1420_ net56 _0650_ _0762_ _0638_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o211a_2
X_1351_ _0670_ _0619_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__or2_2
X_1282_ ByteBuffer.instr\[23\] ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0625_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1618_ RegFile.E\[6\] _0761_ _0771_ RegFile.B\[6\] vssd1 vssd1 vccd1 vccd1 _0961_
+ sky130_fd_sc_hd__a22oi_1
X_2667_ net121 _0144_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.B\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1549_ _0886_ _0888_ _0890_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__o31a_1
X_2598_ clknet_2_3__leaf_clk _0075_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2521_ PC.i_mem_addr\[4\] _0556_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__xor2_1
X_1334_ _0619_ _0640_ _0644_ _0632_ _0645_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__a221o_2
X_1403_ _0740_ _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__nand2_1
X_2383_ _0421_ ByteBuffer.instr\[21\] _0497_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__mux2_1
Xinput3 gpi[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0517_ _0517_ vssd1 vssd1 vccd1 vccd1 clknet_0__0517_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1952_ _0189_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1883_ _0655_ _1221_ _1224_ _0631_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2504_ PC.i_mem_addr\[1\] _0547_ _0542_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__mux2_1
X_2366_ _0493_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__clkbuf_1
X_1317_ ByteBuffer.instr\[20\] ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _0660_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2297_ PC.i_mem_addr\[1\] net46 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap54 _0680_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2082_ RegFile.D\[2\] _0210_ _0289_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__mux2_1
X_2151_ _0336_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
X_2220_ _1049_ _0244_ _0398_ _0655_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1935_ _1143_ _1145_ _1207_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__o21a_1
X_1797_ _0908_ _0885_ _0896_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nand3b_1
X_1866_ _1131_ _1147_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__or2_1
X_2349_ _0485_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2472__7 clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__inv_2
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1651_ _0756_ _0990_ _0991_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__a211o_1
X_1720_ _1057_ _1060_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__o211a_1
X_1582_ RegFile.C\[4\] _0793_ _0794_ RegFile.B\[4\] vssd1 vssd1 vccd1 vccd1 _0925_
+ sky130_fd_sc_hd__a22o_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _0280_ RegFile.L\[2\] _0317_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_1
X_2065_ _0243_ _0262_ _0263_ net2 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a22o_1
X_2203_ _1239_ _0224_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1849_ _1188_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__nand2_4
X_1918_ _1257_ _1175_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1634_ _0972_ _0973_ _0975_ _0976_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2683_ clknet_2_0__leaf_clk _0160_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1703_ _0645_ _1044_ _1045_ ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _1046_
+ sky130_fd_sc_hd__o211a_1
X_1496_ RegFile.A\[3\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__or3_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__buf_2
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ RegFile.C\[6\] _0272_ _0270_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__mux2_1
X_2117_ _0210_ RegFile.H\[2\] _0308_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__mux2_1
Xfanout58 net61 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_8
XFILLER_0_67_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__0514_ clknet_0__0514_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0514_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1350_ _0664_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__nor2_8
X_1281_ ByteBuffer.instr\[18\] vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2666_ net120 _0143_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.B\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2597_ clknet_2_3__leaf_clk _0074_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1617_ _0947_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1479_ RegFile.C\[2\] _0793_ _0786_ RegFile.D\[2\] vssd1 vssd1 vccd1 vccd1 _0822_
+ sky130_fd_sc_hd__a22o_1
X_1548_ RegFile.A\[0\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1402_ ALU.immediate\[9\] _0675_ _0693_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2520_ ALU.immediate\[4\] _0921_ _0519_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__mux2_1
Xinput4 gpi[23] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
X_1333_ _0655_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nor2_4
X_2382_ _0502_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0516_ _0516_ vssd1 vssd1 vccd1 vccd1 clknet_0__0516_ sky130_fd_sc_hd__clkbuf_16
X_2649_ net103 _0126_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.D\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2440__40 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__inv_2
X_1951_ RegFile.A\[3\] _0188_ _1203_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__mux2_1
X_1882_ _1092_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2365_ _0421_ ALU.immediate\[13\] _0407_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__mux2_1
X_2503_ _0545_ _0546_ net47 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1316_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__buf_4
X_2296_ _0243_ _0442_ _0456_ _0445_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__o211a_1
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap55 _0706_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2081_ _0294_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_2150_ ALU.flags_to_alu\[7\] _0328_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1934_ _1114_ _1272_ _1236_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1796_ _1138_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__clkbuf_2
X_1865_ _1151_ _1123_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ MemControl.state\[2\] MemControl.state\[1\] _0411_ vssd1 vssd1 vccd1 vccd1
+ _0485_ sky130_fd_sc_hd__mux2_1
X_2279_ RegFile.A\[2\] net1 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1581_ RegFile.H\[4\] _0784_ _0786_ RegFile.D\[4\] vssd1 vssd1 vccd1 vccd1 _0924_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1650_ _0992_ _0753_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _0381_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2064_ _0283_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
X_2133_ _0322_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1917_ _0780_ _0921_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1848_ ByteBuffer.instr\[20\] _1187_ _1190_ _0700_ _0645_ vssd1 vssd1 vccd1 vccd1
+ _1191_ sky130_fd_sc_hd__a221o_2
X_1779_ _0645_ _1044_ _1045_ ByteBuffer.instr\[19\] vssd1 vssd1 vccd1 vccd1 _1122_
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1633_ RegFile.H\[6\] _0784_ _0817_ RegFile.L\[6\] vssd1 vssd1 vccd1 vccd1 _0976_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ _0622_ _0624_ _0678_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a21o_1
X_2682_ clknet_2_0__leaf_clk _0159_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1564_ _0780_ _0903_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__and3_1
X_1495_ _0834_ _0836_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__or3_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2116_ _0313_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
X_2047_ _1221_ _0262_ _0263_ net9 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a22o_1
Xfanout59 net61 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_8
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2447__46 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__inv_2
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1280_ _0619_ _0622_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2461__60 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
XFILLER_0_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2665_ net119 _0142_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.B\[0\] sky130_fd_sc_hd__dfrtp_2
X_1547_ RegFile.L\[0\] _0817_ _0889_ _0711_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2596_ clknet_2_3__leaf_clk _0073_ net59 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1616_ _0955_ _0693_ _0958_ _0675_ ALU.immediate\[7\] vssd1 vssd1 vccd1 vccd1 _0959_
+ sky130_fd_sc_hd__a32o_2
X_1478_ RegFile.H\[2\] _0784_ _0820_ _0711_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ _0741_ _0743_ _0630_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__and3b_1
X_2381_ _0422_ ByteBuffer.instr\[20\] _0497_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__mux2_1
Xinput5 gpi[2] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
X_1332_ _0664_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__nor2_8
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__0515_ _0515_ vssd1 vssd1 vccd1 vccd1 clknet_0__0515_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2648_ net102 _0125_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.E\[7\] sky130_fd_sc_hd__dfrtp_1
X_2579_ _0610_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ _0655_ _0183_ _0187_ _0631_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1881_ _0718_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__xor2_2
X_2502_ PC.i_mem_addr\[1\] PC.i_mem_addr\[0\] vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__xor2_1
X_2364_ _0492_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
X_1315_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] vssd1 vssd1 vccd1 vccd1 _0658_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2295_ _0455_ _0442_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nand2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap56 _0646_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ RegFile.D\[3\] _0188_ _0289_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1933_ _1113_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1795_ _0883_ _0884_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and2_1
X_1864_ _1120_ _1205_ _1131_ _1166_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__a2bb2o_1
X_2347_ _0484_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
X_2278_ _0447_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2410__11 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__inv_2
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1580_ RegFile.A\[4\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2132_ _0278_ RegFile.L\[3\] _0317_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _1182_ _0204_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ RegFile.C\[1\] _0282_ _0270_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1847_ _1189_ _0666_ _0665_ ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _1190_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1916_ _1254_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__nor2_1
X_1778_ _1098_ _1101_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2681_ clknet_2_0__leaf_clk _0158_ net57 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1701_ _0656_ _0700_ _0624_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__and3b_2
X_1632_ RegFile.B\[6\] _0794_ _0974_ _0711_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a22o_1
X_1494_ RegFile.C\[3\] _0793_ _0786_ RegFile.D\[3\] vssd1 vssd1 vccd1 vccd1 _0837_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1563_ _0904_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__or2_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ _0188_ RegFile.H\[3\] _0308_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ _0271_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2664_ net118 _0141_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.C\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1615_ RegFile.E\[7\] _0709_ _0957_ _0654_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a211o_1
X_1546_ RegFile.E\[0\] _0789_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__or2_1
X_1477_ RegFile.E\[2\] _0789_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__or2_1
X_2595_ clknet_2_2__leaf_clk _0072_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2029_ _0210_ RegFile.B\[2\] _0252_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1400_ RegFile.B\[1\] _0705_ _0742_ _0711_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__a211o_1
X_1331_ _0666_ _0626_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__o21ai_4
X_2380_ _0501_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 gpi[3] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
X_2647_ net101 _0124_ net61 vssd1 vssd1 vccd1 vccd1 RegFile.E\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0514_ _0514_ vssd1 vssd1 vccd1 vccd1 clknet_0__0514_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1529_ RegFile.B\[1\] _0785_ _0708_ _0706_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__and4_1
X_2578_ PC.i_mem_addr\[13\] _0609_ _0542_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1025_ _1088_ net49 vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2431__31 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__inv_2
XFILLER_0_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2501_ _0867_ _0519_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2363_ _0422_ ALU.immediate\[12\] _0407_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
X_2294_ PC.i_mem_addr\[0\] vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
X_1314_ ByteBuffer.instr\[21\] _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1932_ _1106_ _1112_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2_1
X_1863_ _1103_ _1119_ _1124_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ _1057_ _1060_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2346_ _1032_ _0476_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2277_ RegFile.A\[1\] _0445_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _0321_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2062_ _0224_ _0262_ _0263_ net3 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a22o_1
X_2200_ _0243_ _0380_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1846_ _0668_ _0696_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1915_ _1151_ _1048_ _1159_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__and3_1
X_1777_ _1103_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__and2_1
X_2329_ _0474_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ RegFile.E\[6\] _0789_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__or2_1
X_2680_ net70 _0157_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.A\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ _0678_ _1039_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__o21ai_4
X_1493_ RegFile.H\[3\] _0784_ _0835_ _0711_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__a22o_1
X_1562_ RegFile.L\[0\] _0680_ _0687_ ALU.flags_to_alu\[0\] vssd1 vssd1 vccd1 vccd1
+ _0905_ sky130_fd_sc_hd__a22o_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ RegFile.C\[7\] _0264_ _0270_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2114_ _0312_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1829_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2663_ net117 _0140_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.C\[6\] sky130_fd_sc_hd__dfrtp_2
X_1614_ ALU.flags_to_alu\[7\] _0711_ _0707_ RegFile.L\[7\] _0956_ vssd1 vssd1 vccd1
+ vccd1 _0957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2594_ clknet_2_2__leaf_clk _0071_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1476_ ALU.flags_to_alu\[2\] _0788_ _0817_ RegFile.L\[2\] _0818_ vssd1 vssd1 vccd1
+ vccd1 _0819_ sky130_fd_sc_hd__a221o_1
X_1545_ RegFile.H\[0\] _0784_ _0788_ ALU.flags_to_alu\[0\] _0887_ vssd1 vssd1 vccd1
+ vccd1 _0888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2028_ _0257_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2452__51 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__inv_2
XFILLER_0_32_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1330_ _0669_ _0671_ _0672_ _0659_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__o211a_1
Xinput7 gpi[4] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2646_ net100 _0123_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.E\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2577_ _0540_ _0607_ _0608_ _0585_ ALU.immediate\[13\] vssd1 vssd1 vccd1 vccd1 _0609_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1528_ RegFile.H\[1\] _0784_ _0788_ ALU.flags_to_alu\[1\] vssd1 vssd1 vccd1 vccd1
+ _0871_ sky130_fd_sc_hd__a22oi_1
X_1459_ _0630_ _0798_ _0801_ _0693_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__o211ai_4
X_2417__18 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__inv_2
XFILLER_0_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2500_ ALU.immediate\[1\] _0519_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2362_ _0491_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
X_2293_ _0454_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_1313_ _0619_ _0622_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2629_ net83 _0106_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.L\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap47 _0540_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 gpi[7] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dlymetal6s2s_1
X_1862_ _1204_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1931_ _1270_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1793_ _1127_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nand2_2
X_2345_ _0483_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
X_2276_ _0446_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _0276_ RegFile.L\[4\] _0317_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_1
X_2061_ _0281_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1914_ _1151_ _1173_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1845_ _0700_ _1186_ _1187_ ByteBuffer.instr\[19\] _0645_ vssd1 vssd1 vccd1 vccd1
+ _1188_ sky130_fd_sc_hd__a221o_2
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1776_ _0806_ _0936_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2328_ _0445_ _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2259_ _0418_ _0429_ _0419_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ RegFile.C\[6\] _0793_ _0786_ RegFile.D\[6\] vssd1 vssd1 vccd1 vccd1 _0973_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1492_ RegFile.E\[3\] _0789_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__or2_1
X_1561_ RegFile.E\[0\] _0683_ _0685_ RegFile.C\[0\] _0654_ vssd1 vssd1 vccd1 vccd1
+ _0904_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _1269_ RegFile.H\[4\] _0308_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__mux2_1
X_2044_ _0655_ _0265_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__o211a_4
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1828_ _1151_ _1122_ _1159_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__or3b_1
X_1759_ _1100_ _0805_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2438__38 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__inv_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1613_ RegFile.C\[7\] _0708_ net55 vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__and3_1
X_2662_ net116 _0139_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.C\[5\] sky130_fd_sc_hd__dfrtp_2
X_1544_ RegFile.C\[0\] _0792_ _0699_ _0706_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__and4_1
X_2593_ clknet_2_3__leaf_clk _0070_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_1475_ RegFile.B\[2\] _0785_ _0708_ _0706_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__and4_1
X_2027_ _0188_ RegFile.B\[3\] _0252_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 gpi[5] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1527_ RegFile.C\[1\] _0793_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nand2_1
X_2645_ net99 _0122_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.E\[4\] sky130_fd_sc_hd__dfrtp_2
X_2576_ PC.i_mem_addr\[12\] _0597_ PC.i_mem_addr\[13\] vssd1 vssd1 vccd1 vccd1 _0608_
+ sky130_fd_sc_hd__a21o_1
X_1458_ ALU.flags_to_alu\[5\] _0711_ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_
+ sky130_fd_sc_hd__a211o_1
X_1389_ RegFile.A\[2\] _0704_ _0731_ _0630_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2361_ _0490_ ALU.immediate\[11\] _0407_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1312_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__buf_8
X_2292_ _0445_ net46 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2628_ net82 _0105_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.L\[3\] sky130_fd_sc_hd__dfrtp_2
X_2559_ PC.i_mem_addr\[10\] _0588_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap48 _0298_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1930_ RegFile.A\[4\] _1269_ _1203_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput11 nrst vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_2
X_1861_ RegFile.A\[7\] _1184_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1792_ _0935_ _0936_ _1064_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2344_ _0713_ _0476_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ RegFile.A\[0\] _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ RegFile.C\[2\] _0280_ _0270_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _1165_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__inv_2
X_1844_ _0700_ _0641_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nand2_1
X_1775_ _1105_ _1116_ _1117_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2327_ _0440_ _0326_ _0442_ PC.i_mem_addr\[15\] vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__a2bb2o_1
X_2258_ net8 _0420_ _0426_ net7 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__and4bb_1
X_2459__58 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__inv_2
X_2189_ _0248_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ RegFile.A\[0\] net52 _0898_ _0902_ _0629_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2112_ _0311_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
X_1491_ ALU.flags_to_alu\[3\] _0788_ _0817_ RegFile.L\[3\] _0833_ vssd1 vssd1 vccd1
+ vccd1 _0834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ _0655_ _1193_ _1201_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1827_ _1069_ _1164_ _1167_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a211o_1
X_1689_ RegFile.A\[7\] _0704_ _1031_ _0630_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1758_ _1100_ _0805_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2661_ net115 _0138_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.C\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1474_ _0789_ _0699_ net55 vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and3_2
X_1612_ _0948_ _0954_ _0629_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__a21o_1
X_1543_ RegFile.D\[0\] _0786_ _0794_ RegFile.B\[0\] vssd1 vssd1 vccd1 vccd1 _0886_
+ sky130_fd_sc_hd__a22o_1
X_2592_ clknet_2_0__leaf_clk _0069_ net57 vssd1 vssd1 vccd1 vccd1 ByteDecoder.num_bytes\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2026_ _0256_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 gpi[6] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
X_2644_ net98 _0121_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.E\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1457_ RegFile.E\[5\] _0699_ _0706_ _0654_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__a31o_1
X_2575_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__inv_2
X_1526_ ALU.immediate\[1\] _0675_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1388_ RegFile.B\[2\] _0705_ _0730_ _0711_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a211o_1
X_2009_ net49 _1079_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1311_ _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__clkbuf_8
X_2291_ _0262_ _0413_ _0445_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__a21boi_2
X_2360_ net6 _0417_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2422__23 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__inv_2
XFILLER_0_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2627_ net81 _0104_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.L\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1509_ RegFile.L\[3\] net54 _0685_ RegFile.C\[3\] vssd1 vssd1 vccd1 vccd1 _0852_
+ sky130_fd_sc_hd__a22o_1
X_2558_ PC.i_mem_addr\[10\] _0588_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__nand2_1
X_2489_ _0523_ _0529_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__o21ai_2
Xmax_cap49 _1043_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_6
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _1192_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__nor2_4
XFILLER_0_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1791_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__xnor2_1
X_2343_ _0482_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
X_2274_ net1 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__buf_6
X_1989_ _0756_ _0990_ _0993_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__0517_ clknet_0__0517_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0517_
+ sky130_fd_sc_hd__clkbuf_16
X_1843_ ByteBuffer.instr\[20\] _0665_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _0938_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__or2_1
X_1774_ _0806_ _0936_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__xnor2_1
X_2326_ _1224_ _0442_ _0472_ _0445_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__o211a_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2257_ _0419_ _0425_ _0430_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__o211ai_2
X_2188_ _1069_ _1092_ _1093_ _1131_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1490_ RegFile.B\[3\] _0785_ _0708_ _0706_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _1247_ RegFile.H\[5\] _0308_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2042_ _0630_ _0267_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or2_2
Xhold1 ByteDecoder.num_bytes\[1\] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1826_ _1075_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__nor2_1
X_1688_ RegFile.B\[7\] _0705_ _1030_ _0711_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1757_ _1099_ _1095_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2309_ PC.i_mem_addr\[7\] net46 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ _0949_ _0950_ _0952_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or4_1
X_2660_ net114 _0137_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.C\[3\] sky130_fd_sc_hd__dfrtp_1
X_2591_ clknet_2_0__leaf_clk _0068_ net57 vssd1 vssd1 vccd1 vccd1 ByteDecoder.num_bytes\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1473_ _0780_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_4
X_1542_ ALU.immediate\[0\] _0664_ _0692_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__o21ai_2
X_2429__29 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__inv_2
X_2025_ _1269_ RegFile.B\[4\] _0252_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1809_ _1130_ _1148_ _1149_ _1151_ _1123_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a2111oi_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2443__43 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__inv_2
XFILLER_0_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2643_ net97 _0120_ net61 vssd1 vssd1 vccd1 vccd1 RegFile.E\[2\] sky130_fd_sc_hd__dfrtp_1
X_2574_ PC.i_mem_addr\[12\] PC.i_mem_addr\[13\] _0597_ vssd1 vssd1 vccd1 vccd1 _0606_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1456_ RegFile.C\[5\] _0705_ _0707_ RegFile.L\[5\] vssd1 vssd1 vccd1 vccd1 _0799_
+ sky130_fd_sc_hd__a22o_1
X_1387_ RegFile.H\[2\] _0707_ _0709_ RegFile.D\[2\] vssd1 vssd1 vccd1 vccd1 _0730_
+ sky130_fd_sc_hd__a22o_1
X_1525_ _0675_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2008_ _1166_ _0232_ _0236_ _0242_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a211o_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2290_ _0453_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_1310_ _0623_ _0628_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2626_ net80 _0103_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.L\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2557_ _0592_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ ALU.flags_to_alu\[3\] _0687_ _0683_ RegFile.E\[3\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0851_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _0678_ _0636_ _0526_ _0530_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__o41a_1
X_1439_ ALU.immediate\[5\] _0675_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1790_ _1072_ _1127_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nand2_1
X_2342_ _1006_ _0476_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and2_1
X_2273_ MemControl.state\[0\] _0443_ _0444_ net134 vssd1 vssd1 vccd1 vccd1 _0000_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1988_ _1142_ _1207_ _0213_ _0223_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a31o_4
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2609_ clknet_2_0__leaf_clk _0086_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__0516_ clknet_0__0516_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0516_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1842_ _0642_ _0666_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nor2_1
X_1911_ _0937_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__nor2_1
X_1773_ _1114_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
X_2325_ PC.i_mem_addr\[14\] net46 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__or2_1
X_2187_ _1050_ _1212_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nand2_1
X_2256_ ByteDecoder.state\[1\] ByteDecoder.state\[0\] vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _0310_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2041_ _0266_ _1191_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nor2_1
Xhold2 FSM.next_state\[0\] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dlygate4sd3_1
X_2464__63 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1756_ _0970_ _0982_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1825_ _1043_ _1122_ _1159_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__or3b_4
X_1687_ RegFile.H\[7\] _0707_ _0709_ RegFile.D\[7\] vssd1 vssd1 vccd1 vccd1 _1030_
+ sky130_fd_sc_hd__a22o_1
X_2308_ _1221_ _0442_ _0462_ _0445_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__o211a_1
X_2239_ ByteDecoder.state\[0\] vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1610_ RegFile.H\[7\] _0784_ _0817_ RegFile.L\[7\] vssd1 vssd1 vccd1 vccd1 _0953_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2590_ clknet_2_0__leaf_clk _0067_ net57 vssd1 vssd1 vccd1 vccd1 ByteDecoder.num_bytes\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1472_ _0629_ _0812_ _0813_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1541_ _0675_ _0867_ _0869_ _0880_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__o211ai_1
X_2024_ _0255_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1739_ _1054_ _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__a21o_1
X_1808_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__buf_6
XFILLER_0_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2642_ net96 _0119_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.E\[1\] sky130_fd_sc_hd__dfrtp_2
X_1524_ _0629_ _0862_ _0863_ _0865_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__o32a_4
X_2573_ _0605_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1455_ _0787_ _0791_ _0796_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o31a_1
X_1386_ RegFile.A\[2\] _0652_ _0676_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2007_ _0237_ _0238_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1507_ _0847_ _0848_ _0849_ _0774_ RegFile.A\[3\] vssd1 vssd1 vccd1 vccd1 _0850_
+ sky130_fd_sc_hd__o32a_1
X_2625_ net79 _0102_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.L\[0\] sky130_fd_sc_hd__dfrtp_2
X_2556_ PC.i_mem_addr\[9\] _0591_ _0542_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__mux2_1
X_2487_ ByteBuffer.instr\[20\] _0343_ _0531_ _0636_ vssd1 vssd1 vccd1 vccd1 _0532_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1369_ RegFile.B\[6\] _0705_ _0710_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1438_ _0629_ _0775_ _0778_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2413__14 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__inv_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2341_ _0481_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2272_ _0411_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _1166_ _0212_ _0215_ _1124_ _0222_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2608_ clknet_2_1__leaf_clk _0085_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_2539_ _0577_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1910_ _0832_ _0856_ _0912_ _0913_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o31a_1
Xclkbuf_1_0__f__0515_ clknet_0__0515_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0515_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1841_ _0631_ _1094_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a21bo_1
X_1772_ _0937_ _0913_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2324_ _1246_ _0442_ _0471_ _0445_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__o211a_1
X_2186_ _1066_ _1092_ _1158_ _0347_ _1181_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o221a_1
X_2255_ _0427_ _0428_ _0418_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2040_ _1188_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
Xhold3 ByteDecoder.num_bytes\[2\] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1686_ RegFile.A\[7\] _0652_ _1028_ _0676_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1755_ _1096_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__and2_1
X_1824_ ALU.flags_to_alu\[0\] _1151_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_
+ sky130_fd_sc_hd__a31o_1
X_2307_ PC.i_mem_addr\[6\] net46 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__or2_1
X_2238_ ByteDecoder.state\[1\] ByteDecoder.num_bytes\[2\] ByteDecoder.num_bytes\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nor3_1
X_2169_ _0816_ _1049_ _1166_ _1137_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2468__3 clknet_1_0__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ _0675_ _0867_ _0880_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__or3_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1471_ RegFile.L\[2\] _0680_ _0685_ RegFile.C\[2\] vssd1 vssd1 vccd1 vccd1 _0814_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2023_ _1247_ RegFile.B\[5\] _0252_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1807_ _0678_ _1039_ _1042_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1669_ RegFile.D\[4\] _0683_ net53 RegFile.B\[4\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _1012_ sky130_fd_sc_hd__a221o_1
X_1738_ _0740_ _0745_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__and2b_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2419__20 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__inv_2
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2434__34 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__inv_2
X_1523_ ALU.flags_to_alu\[1\] _0652_ _0629_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__o21ai_1
X_1454_ RegFile.A\[5\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__or3_1
X_2641_ net95 _0118_ net59 vssd1 vssd1 vccd1 vccd1 RegFile.E\[0\] sky130_fd_sc_hd__dfrtp_2
X_2572_ PC.i_mem_addr\[12\] _0604_ _0542_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1385_ RegFile.H\[2\] _0680_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a21o_1
X_2408__9 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_2
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _1140_ _0239_ _0240_ _1043_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2624_ net78 _0101_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1506_ ALU.flags_to_alu\[3\] _0765_ _0763_ RegFile.H\[3\] vssd1 vssd1 vccd1 vccd1
+ _0849_ sky130_fd_sc_hd__a22o_1
X_2555_ _0540_ _0589_ _0590_ _0585_ ALU.immediate\[9\] vssd1 vssd1 vccd1 vccd1 _0591_
+ sky130_fd_sc_hd__a32o_1
X_2486_ _0678_ _0524_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1437_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__buf_4
X_1368_ _0708_ net55 vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__nor2_8
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1299_ ByteBuffer.instr\[17\] _0624_ ByteBuffer.instr\[19\] _0619_ vssd1 vssd1 vccd1
+ vccd1 _0642_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _1017_ _0476_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__and2_1
X_2271_ _0261_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1986_ _0816_ _1253_ _0216_ _0221_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2607_ clknet_2_1__leaf_clk _0084_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2538_ PC.i_mem_addr\[6\] _0576_ _0542_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__mux2_1
Xwire50 _0875_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1840_ _0655_ _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0514_ clknet_0__0514_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0514_
+ sky130_fd_sc_hd__clkbuf_16
X_1771_ _1106_ _1112_ _1113_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2323_ PC.i_mem_addr\[13\] net46 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2254_ net9 _0417_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__and2_1
X_2185_ _0363_ _0364_ _0362_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _0205_ _1082_ net49 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 ByteDecoder.num_bytes\[3\] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1823_ _1151_ _1049_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nor2_4
X_1685_ RegFile.H\[7\] net54 _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1754_ _0960_ _1095_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__or2_1
X_2237_ _0410_ _0411_ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__or3_2
X_2306_ _1239_ _0442_ _0461_ _0445_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__o211a_1
X_2455__54 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__inv_2
X_2099_ RegFile.E\[2\] _0280_ net48 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _1093_ _1136_ _0347_ _1252_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ ALU.flags_to_alu\[2\] _0687_ _0683_ RegFile.E\[2\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2022_ _0254_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _1130_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__nor2_1
X_1599_ RegFile.L\[7\] _0770_ _0763_ RegFile.H\[7\] net52 vssd1 vssd1 vccd1 vccd1
+ _0942_ sky130_fd_sc_hd__a221o_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _1009_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1737_ _1055_ _1079_ _0754_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a21bo_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470__5 clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__inv_2
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ net94 _0117_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1522_ RegFile.L\[1\] net54 _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__a21oi_1
X_1453_ RegFile.C\[5\] _0793_ _0794_ RegFile.B\[5\] _0795_ vssd1 vssd1 vccd1 vccd1
+ _0796_ sky130_fd_sc_hd__a221o_1
X_2571_ _0540_ _0602_ _0603_ _0585_ ALU.immediate\[12\] vssd1 vssd1 vccd1 vccd1 _0604_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1384_ RegFile.D\[2\] _0683_ net53 RegFile.B\[2\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0727_ sky130_fd_sc_hd__a221o_1
X_2005_ _0947_ _1214_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ net77 _0100_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[6\] sky130_fd_sc_hd__dfrtp_2
X_2554_ PC.i_mem_addr\[9\] _0582_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1367_ RegFile.H\[6\] _0707_ _0709_ RegFile.D\[6\] vssd1 vssd1 vccd1 vccd1 _0710_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1505_ RegFile.D\[3\] _0767_ _0771_ RegFile.B\[3\] vssd1 vssd1 vccd1 vccd1 _0848_
+ sky130_fd_sc_hd__a22o_1
X_2485_ _0327_ _0525_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1436_ _0664_ _0674_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__or2_1
X_1298_ _0619_ _0622_ _0624_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2270_ net133 _0411_ _0410_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _1213_ _0218_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__o21ba_1
X_2537_ _0572_ _0575_ net47 vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2606_ clknet_2_1__leaf_clk _0083_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1419_ _0670_ _0757_ _0759_ _0650_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__a31oi_4
X_2399_ _0421_ ALU.immediate\[5\] _0409_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire51 _0772_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ _1104_ _0856_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2322_ _1268_ _0442_ _0470_ _0445_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__o211a_1
X_2184_ _0362_ _0363_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__or3_1
X_2253_ net2 _0420_ _0421_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1899_ _1086_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__inv_2
X_1968_ _0746_ _0994_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 ByteBuffer.counter\[0\] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1753_ _0960_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__nand2_1
X_1822_ _1048_ _1163_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nor2_2
X_1684_ RegFile.D\[7\] _0683_ net53 RegFile.B\[7\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _1027_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2236_ MemControl.state\[2\] MemControl.state\[1\] MemControl.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _0412_ sky130_fd_sc_hd__o21ba_2
X_2167_ _1257_ _1049_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand2_1
X_2305_ PC.i_mem_addr\[5\] net46 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or2_1
X_2098_ _0303_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2021_ _1225_ RegFile.B\[6\] _0252_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1736_ _0960_ _0983_ _1064_ _1065_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__a41o_1
X_1805_ _1131_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__nand2_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1598_ ALU.flags_to_alu\[7\] _0765_ _0767_ RegFile.D\[7\] _0940_ vssd1 vssd1 vccd1
+ vccd1 _0941_ sky130_fd_sc_hd__a221o_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1003_ _1007_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nor2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2219_ _1213_ _0990_ _0394_ _0396_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2570_ PC.i_mem_addr\[12\] _0597_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1521_ RegFile.E\[1\] _0683_ _0685_ RegFile.C\[1\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0864_ sky130_fd_sc_hd__a221o_1
X_1452_ RegFile.L\[5\] _0789_ _0699_ net55 vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__and4_1
X_1383_ _0721_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2004_ _1059_ _1161_ _1255_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1719_ _0816_ _0831_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__or2b_1
X_2699_ clknet_2_1__leaf_clk net129 net61 vssd1 vssd1 vccd1 vccd1 ByteDecoder.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2622_ net76 _0099_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[5\] sky130_fd_sc_hd__dfrtp_4
X_1504_ RegFile.E\[3\] _0761_ _0845_ _0846_ net51 vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2553_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1435_ _0776_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__or2_2
X_1366_ _0708_ _0703_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__nor2_4
X_2484_ _0524_ _0525_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__mux2_1
X_1297_ ByteBuffer.instr\[20\] _0639_ _0632_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1984_ _0197_ _1254_ _1164_ _0908_ _0219_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2536_ _0573_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__nor2_1
X_2605_ clknet_2_0__leaf_clk _0082_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1418_ _0684_ _0677_ _0679_ _0760_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__and4_4
X_1349_ _0666_ _0626_ _0673_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o21a_2
XFILLER_0_3_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _0510_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2321_ PC.i_mem_addr\[12\] net46 vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or2_1
X_2183_ _1092_ _1223_ _0228_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2252_ net3 net5 net6 _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__or4b_1
XFILLER_0_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _1166_ _1137_ _0191_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1898_ _1147_ _1228_ _1234_ _1238_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__o211ai_4
X_2519_ _0560_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6 MemControl.state\[2\] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1683_ _0718_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nor2_1
X_1752_ _0970_ _0982_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1821_ _1122_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__nor2_2
X_2304_ _1265_ _0442_ _0460_ _0445_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__o211a_1
X_2097_ RegFile.E\[3\] _0278_ net48 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__mux2_1
X_2166_ _1151_ _1092_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__nand2_2
X_2235_ _0670_ _0659_ _0662_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__and3_2
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2020_ _0253_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1666_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1804_ _1134_ _1136_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nor3_2
X_1735_ _1067_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ RegFile.C\[7\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__and4_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2149_ _0659_ _1201_ _0333_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a31o_2
X_2218_ _0908_ _1165_ _0240_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1520_ RegFile.A\[1\] _0774_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__nor2_1
X_1451_ _0785_ _0708_ _0706_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__and3_2
X_1382_ ALU.immediate\[11\] _0675_ _0693_ _0724_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a22o_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2003_ _0908_ _1175_ _1165_ _0197_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2425__26 clknet_1_1__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__inv_2
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1649_ _0749_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__inv_2
X_2698_ clknet_2_1__leaf_clk _0001_ net61 vssd1 vssd1 vccd1 vccd1 MemControl.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1718_ _0855_ _0844_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1503_ RegFile.L\[3\] _0638_ _0681_ _0762_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__and4_1
X_2621_ net75 _0098_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2552_ PC.i_mem_addr\[9\] _0582_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__and2_1
X_2483_ _0404_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1434_ RegFile.L\[5\] net54 _0687_ ALU.flags_to_alu\[5\] vssd1 vssd1 vccd1 vccd1
+ _0777_ sky130_fd_sc_hd__a22o_1
X_1365_ _0694_ _0698_ _0648_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1296_ _0624_ ByteBuffer.instr\[17\] vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1983_ _0197_ _1175_ _1162_ _1139_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a2bb2o_1
X_2604_ clknet_2_1__leaf_clk _0081_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1417_ _0670_ _0757_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and3_4
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2535_ PC.i_mem_addr\[6\] _0567_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1348_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__inv_2
X_1279_ ByteBuffer.instr\[17\] vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__buf_6
X_2397_ _0422_ ALU.immediate\[4\] _0409_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2320_ _0187_ _0442_ _0469_ _0445_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__o211a_1
X_2251_ net2 _0417_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__and2_1
X_2182_ _1092_ _1223_ _0228_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1966_ _0192_ _0193_ _0202_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1897_ _1049_ _1235_ _1237_ _1118_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__o22a_1
X_2518_ PC.i_mem_addr\[3\] _0559_ _0542_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 MemControl.state\[1\] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1820_ ByteBuffer.instr\[21\] _0645_ _1044_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__or3b_2
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1682_ _1000_ _1011_ _1022_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o31a_1
X_1751_ _1038_ _1051_ _1090_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o22ai_4
X_2234_ MemControl.state\[0\] _0261_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__and2_1
X_2303_ PC.i_mem_addr\[4\] net46 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or2_1
X_2096_ _0302_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2165_ _1094_ _0187_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__xor2_1
X_1949_ _0726_ _0185_ _0186_ _1092_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1803_ _1143_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__nand2_1
X_1596_ RegFile.E\[7\] _0761_ _0771_ RegFile.B\[7\] vssd1 vssd1 vccd1 vccd1 _0939_
+ sky130_fd_sc_hd__a22o_1
X_1665_ _1003_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1734_ _1070_ _1074_ _1075_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__a211o_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ ALU.flags_to_alu\[0\] _1151_ _1122_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_
+ sky130_fd_sc_hd__a31o_1
X_2079_ _0293_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
X_2148_ _1192_ _0630_ _1202_ _0287_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1450_ _0792_ _0699_ _0706_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__and3_2
X_1381_ RegFile.A\[3\] _0704_ _0723_ _0630_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2002_ ALU.flags_to_alu\[0\] _1151_ _1164_ _1254_ _0908_ vssd1 vssd1 vccd1 vccd1
+ _0237_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1648_ _0740_ _0745_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__nor2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2697_ clknet_2_1__leaf_clk net135 net61 vssd1 vssd1 vccd1 vccd1 MemControl.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1717_ _1058_ _1059_ _0883_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o21a_1
X_1579_ _0780_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__nand2_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2430__30 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__inv_2
X_2620_ net74 _0097_ net59 vssd1 vssd1 vccd1 vccd1 ALU.flags_to_alu\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1433_ RegFile.E\[5\] _0683_ _0685_ RegFile.C\[5\] _0654_ vssd1 vssd1 vccd1 vccd1
+ _0776_ sky130_fd_sc_hd__a221o_1
X_1502_ RegFile.C\[3\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2482_ _0678_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nor2_1
X_2551_ _0587_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
X_1364_ _0699_ net55 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nor2_8
XFILLER_0_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1295_ _0622_ _0632_ _0634_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1982_ _0910_ _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__nand2_1
X_2534_ PC.i_mem_addr\[6\] _0567_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2603_ clknet_2_1__leaf_clk _0080_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1347_ RegFile.A\[6\] _0652_ _0676_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o211a_1
X_1416_ _0700_ _0758_ _0647_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2396_ _0509_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1278_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or2_2
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _0420_ _0421_ _0422_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o31a_1
X_2181_ _1246_ _1268_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1965_ _1213_ _0195_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1896_ _1117_ _1105_ _1116_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2517_ _0555_ _0558_ net47 vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2379_ _0490_ ByteBuffer.instr\[19\] _0497_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 _0000_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ net49 _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nand2_4
XFILLER_0_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1681_ _1023_ _1007_ _1011_ _1020_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o22a_1
X_2164_ _0278_ _0334_ _0337_ net138 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__a22o_1
X_2233_ _0407_ _0409_ vssd1 vssd1 vccd1 vccd1 ByteBuffer.next_counter\[1\] sky130_fd_sc_hd__nand2_1
X_2302_ _0183_ _0442_ _0459_ _0445_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__o211a_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2095_ RegFile.E\[4\] _0276_ net48 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1948_ _0726_ _0185_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__nand2_1
X_1879_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1802_ _1144_ _1113_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1733_ _1069_ _0982_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__nor2_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ ALU.immediate\[13\] _0675_ _0693_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1595_ _0832_ _0856_ _0912_ _0913_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o311a_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ _0332_ _0626_ _0645_ _1197_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2216_ ALU.flags_to_alu\[0\] _1151_ _1173_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2078_ RegFile.D\[4\] _1269_ _0289_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_1
X_2451__50 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__inv_2
XFILLER_0_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ RegFile.B\[3\] _0705_ _0722_ _0711_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2001_ _0232_ _0233_ _0234_ _1162_ _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__o32a_1
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2696_ clknet_2_2__leaf_clk _0173_ net58 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1716_ _0885_ _0896_ _0908_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a21bo_1
X_1578_ _0629_ _0918_ _0919_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__o22a_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1647_ _0806_ _0938_ _0984_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a31o_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2416__17 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__inv_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ PC.i_mem_addr\[8\] _0586_ _0542_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1432_ _0764_ _0769_ _0773_ _0774_ RegFile.A\[5\] vssd1 vssd1 vccd1 vccd1 _0775_
+ sky130_fd_sc_hd__o32a_2
X_1363_ _0622_ _0701_ _0702_ _0626_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__o22ai_4
X_2481_ ByteBuffer.instr\[20\] _0639_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__nand2_1
X_1501_ ALU.immediate\[3\] _0674_ _0843_ _0830_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1294_ _0626_ _0635_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__and3b_1
X_2679_ net69 _0156_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.A\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1981_ _1139_ _0909_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__nand2_1
X_2602_ clknet_2_1__leaf_clk _0079_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_2533_ ALU.immediate\[6\] _0969_ _0519_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1346_ RegFile.H\[6\] net54 _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1415_ _0619_ _0622_ ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__a21bo_1
X_2395_ _0490_ ALU.immediate\[3\] _0409_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__mux2_1
X_1277_ ByteBuffer.instr\[17\] vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2180_ _0346_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1964_ _0196_ _0198_ _0199_ _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__or4b_1
X_1895_ _1043_ _1123_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2516_ _0556_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _0645_ ByteBuffer.instr\[22\] vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__xnor2_4
X_2378_ _0500_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold9 ALU.flags_to_alu\[1\] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _1003_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__inv_2
X_2301_ PC.i_mem_addr\[3\] net46 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
X_2163_ _0276_ _0334_ _0337_ net137 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a22o_1
X_2232_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__clkbuf_4
X_2094_ _0301_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1947_ _0997_ _0184_ net49 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _1206_ _1209_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2437__37 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__inv_2
XFILLER_0_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1663_ RegFile.A\[5\] _0704_ _1005_ _0630_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1732_ _1066_ _0959_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nor2_1
X_1801_ _1057_ _1060_ _1062_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1594_ _0935_ _0936_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _0292_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
X_2146_ _0647_ _0329_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__o21a_1
X_2215_ _1149_ _1079_ _1207_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2000_ _1059_ _1123_ _1141_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2695_ clknet_2_2__leaf_clk _0172_ net59 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1715_ _0675_ _0867_ _0869_ _0880_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1646_ _0984_ _0985_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a21bo_1
X_1577_ RegFile.L\[4\] net54 net53 RegFile.C\[4\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a22o_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2129_ _0320_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1500_ _0655_ _0838_ _0839_ _0842_ _0828_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__a311o_1
X_2480_ _0678_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1362_ _0699_ _0703_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__nor2_8
X_1431_ _0760_ _0652_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__or2_2
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1293_ _0624_ _0622_ ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1629_ ALU.flags_to_alu\[6\] _0788_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__and2_1
X_2678_ net68 _0155_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.A\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1980_ _0883_ _1172_ _1168_ _1058_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2532_ _0571_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
X_2601_ clknet_2_1__leaf_clk _0078_ net58 vssd1 vssd1 vccd1 vccd1 ByteBuffer.instr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1345_ RegFile.D\[6\] _0683_ net53 RegFile.B\[6\] _0687_ vssd1 vssd1 vccd1 vccd1
+ _0688_ sky130_fd_sc_hd__a221o_1
X_1414_ ByteBuffer.instr\[22\] _0642_ _0635_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__or3_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2394_ _0508_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
X_1276_ ByteBuffer.instr\[16\] vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1963_ _1256_ _1175_ _0816_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__mux2_1
X_1894_ _1151_ _1134_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2_1
X_2446_ clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__buf_1
X_2515_ PC.i_mem_addr\[3\] _0551_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
X_2458__57 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__inv_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1328_ _0670_ _0661_ _0639_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__or3_1
X_2377_ _0435_ _0624_ _0497_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2231_ ByteBuffer.counter\[1\] _0659_ ByteBuffer.counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0408_ sky130_fd_sc_hd__or3b_1
X_2300_ _0204_ _0442_ _0458_ _0445_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__o211a_1
X_2093_ RegFile.E\[5\] _0274_ net48 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__mux2_1
X_2162_ _0274_ _0334_ _0337_ net139 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1946_ _0736_ _1082_ _0734_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1877_ _1100_ _1210_ _1212_ _1213_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1800_ _1137_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1662_ RegFile.B\[5\] _0705_ _1004_ _0711_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1731_ _1071_ _1072_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__a21o_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _1124_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1593_ _0922_ _0934_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2076_ RegFile.D\[5\] _1247_ _0289_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__mux2_1
X_2145_ _0330_ _0696_ _0618_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__a21o_1
X_1929_ _0655_ _1265_ _1268_ _0631_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1576_ ALU.flags_to_alu\[4\] _0687_ _0683_ RegFile.E\[4\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0919_ sky130_fd_sc_hd__a221o_1
X_2694_ clknet_2_2__leaf_clk _0171_ net59 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1645_ _0986_ _0970_ _0982_ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__o31a_1
X_1714_ _0816_ _0831_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__xor2_4
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2128_ _0274_ RegFile.L\[5\] _0317_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__mux2_1
X_2059_ _0204_ _0262_ _0263_ net5 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a22o_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1430_ RegFile.L\[5\] _0770_ _0771_ RegFile.B\[5\] net52 vssd1 vssd1 vccd1 vccd1
+ _0773_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1361_ _0699_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__nand2_8
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1292_ ByteBuffer.instr\[17\] _0624_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__xor2_4
X_2421__22 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__inv_2
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1628_ RegFile.A\[6\] _0792_ _0704_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__or3_1
X_2677_ net67 _0154_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.A\[4\] sky130_fd_sc_hd__dfrtp_4
X_1559_ RegFile.E\[0\] _0761_ _0899_ _0900_ _0901_ vssd1 vssd1 vccd1 vccd1 _0902_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2600_ clknet_2_3__leaf_clk _0077_ net57 vssd1 vssd1 vccd1 vccd1 ALU.immediate\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1413_ _0754_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nand2_2
XFILLER_0_23_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2393_ _0435_ ALU.immediate\[2\] _0409_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
X_2531_ PC.i_mem_addr\[5\] _0570_ _0542_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1344_ _0686_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__clkbuf_8
X_1275_ ByteBuffer.instr\[19\] vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _1210_ _1168_ _1057_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1893_ _0806_ _1210_ _1229_ _1213_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__o221a_1
X_2376_ _0499_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
X_2514_ PC.i_mem_addr\[3\] _0551_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__and2_1
X_1327_ _0645_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2230_ ByteBuffer.counter\[1\] ByteBuffer.next_counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0407_ sky130_fd_sc_hd__nand2_4
X_2092_ _0300_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2161_ net140 _0337_ _0344_ _0345_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1945_ _1273_ _0180_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__o21a_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1876_ _1070_ _1172_ _1216_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2359_ _0489_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1661_ RegFile.H\[5\] _0707_ _0709_ RegFile.D\[5\] vssd1 vssd1 vccd1 vccd1 _1004_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ _0922_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nor2_2
X_1730_ _0781_ _0782_ _0802_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__nand2_1
X_2213_ _1096_ _1125_ _0986_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
X_2075_ _0291_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
X_2428__28 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__inv_2
XFILLER_0_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1859_ _0630_ _1193_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__o21bai_4
X_1928_ _1022_ _1266_ _1267_ _1092_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2442__42 clknet_1_1__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__inv_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1713_ _0855_ _0844_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__nor2_1
X_1575_ _0914_ _0916_ _0917_ _0774_ RegFile.A\[4\] vssd1 vssd1 vccd1 vccd1 _0918_
+ sky130_fd_sc_hd__o32a_1
X_2693_ clknet_2_2__leaf_clk _0170_ net59 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1644_ _0947_ _0959_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__or2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _0319_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2058_ _0279_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _0622_ _0701_ _0702_ _0626_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o22a_4
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1291_ ByteBuffer.instr\[20\] _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2676_ net66 _0153_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.A\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1558_ net56 _0650_ _0762_ _0684_ ALU.flags_to_alu\[0\] vssd1 vssd1 vccd1 vccd1 _0901_
+ sky130_fd_sc_hd__o2111a_1
X_1627_ _0780_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nand2_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _0816_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__nor2_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2530_ _0566_ _0569_ net47 vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__mux2_1
X_1343_ _0684_ _0677_ _0679_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__and3_1
X_1412_ _0749_ _0753_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__or2_1
X_2392_ _0507_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2659_ net113 _0136_ net61 vssd1 vssd1 vccd1 vccd1 RegFile.C\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1961_ _0855_ _1165_ _1164_ _0197_ _1166_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__a221o_1
X_1892_ _1073_ _1168_ _1231_ _1232_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2513_ ALU.immediate\[3\] _0853_ _0519_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__mux2_1
X_1326_ _0667_ _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nor2_1
X_2375_ _0436_ _0622_ _0497_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2449__48 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__inv_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2160_ _1201_ _0272_ _0335_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2091_ RegFile.E\[6\] _0272_ _0298_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_1
X_2463__62 clknet_1_1__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
XFILLER_0_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1944_ _0181_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_1875_ _1175_ _1174_ _1069_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2289_ RegFile.A\[7\] net1 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__and2_1
X_1309_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__buf_4
X_2358_ _0435_ ALU.immediate\[10\] _0407_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ RegFile.A\[5\] _0652_ _0676_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__o211a_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ ALU.immediate\[4\] _0675_ _0929_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _0282_ _0391_ _0335_ net136 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__o22a_1
X_2143_ _0619_ _0668_ _0620_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a21oi_1
X_2074_ RegFile.D\[6\] _1225_ _0289_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1927_ _1022_ _1266_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nand2_1
X_1858_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__clkbuf_4
X_1789_ _0806_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2692_ clknet_2_2__leaf_clk _0169_ net59 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1712_ _0756_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__inv_2
X_1643_ _0947_ _0959_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1574_ RegFile.L\[4\] _0770_ _0771_ RegFile.B\[4\] net52 vssd1 vssd1 vccd1 vccd1
+ _0917_ sky130_fd_sc_hd__a221o_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _0272_ RegFile.L\[6\] _0317_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__mux2_1
X_2057_ RegFile.C\[3\] _0278_ _0270_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__mux2_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1290_ _0619_ _0622_ _0624_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_58_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1626_ _0654_ _0966_ _0967_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o2bb2a_2
X_2675_ net65 _0152_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.A\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1557_ net56 _0650_ _0766_ _0684_ RegFile.D\[0\] vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__o2111a_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ ALU.immediate\[2\] _0674_ _0829_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__o211a_4
X_2109_ _1225_ RegFile.H\[6\] _0308_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2412__13 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__inv_2
X_2466__1 clknet_1_1__leaf__0514_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1342_ _0677_ _0679_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__a21oi_4
X_1411_ _0749_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__nand2_1
X_2391_ _0436_ ALU.immediate\[1\] _0409_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1609_ RegFile.B\[7\] _0794_ _0951_ _0711_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__a22o_1
X_2658_ net112 _0135_ net60 vssd1 vssd1 vccd1 vccd1 RegFile.C\[1\] sky130_fd_sc_hd__dfrtp_2
X_2589_ clknet_2_1__leaf_clk _0066_ net58 vssd1 vssd1 vccd1 vccd1 MemControl.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1960_ _0675_ _0867_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__nor2_1
X_1891_ _1174_ _1175_ _0781_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2512_ _0554_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1325_ ByteBuffer.instr\[20\] ByteBuffer.instr\[21\] vssd1 vssd1 vccd1 vccd1 _0668_
+ sky130_fd_sc_hd__nand2b_1
X_2374_ _0498_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ _0299_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1943_ _1093_ _1145_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__nor2_1
X_1874_ _0781_ _1214_ _1076_ _1168_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__o221a_1
X_2426_ clknet_1_0__leaf__0514_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1308_ _0638_ net56 _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or3_1
X_2288_ _0452_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2357_ _0488_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _0930_ _0931_ _0932_ _0693_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2073_ _0290_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _0334_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2142_ _0264_ _0327_ _1201_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1926_ _1000_ _1085_ net49 vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__mux2_1
X_1857_ _1196_ _0627_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1788_ _0983_ _1128_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433__33 clknet_1_0__leaf__0516_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__inv_2
XFILLER_0_45_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2691_ clknet_2_2__leaf_clk _0168_ net59 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_1711_ _0746_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1642_ _0804_ _0935_ _0805_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1573_ ALU.flags_to_alu\[4\] _0765_ _0767_ RegFile.D\[4\] _0915_ vssd1 vssd1 vccd1
+ vccd1 _0916_ sky130_fd_sc_hd__a221o_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _0318_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
X_2056_ _0183_ _0262_ _0263_ net6 vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a22o_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1909_ _1136_ _1146_ _1207_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1625_ RegFile.L\[6\] net54 _0685_ RegFile.C\[6\] vssd1 vssd1 vccd1 vccd1 _0968_
+ sky130_fd_sc_hd__a22o_1
X_2674_ net64 _0151_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.A\[1\] sky130_fd_sc_hd__dfrtp_4
X_1556_ net56 _0650_ _0762_ _0638_ RegFile.H\[0\] vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _0664_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__inv_2
X_2108_ _0309_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
X_2039_ _1188_ _1191_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1410_ ALU.immediate\[8\] _0675_ _0693_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1341_ _0637_ _0634_ _0632_ _0622_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2390_ _0506_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1608_ RegFile.E\[7\] _0789_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__or2_1
X_2657_ net111 _0134_ net61 vssd1 vssd1 vccd1 vccd1 RegFile.C\[0\] sky130_fd_sc_hd__dfrtp_1
X_2588_ _0617_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_1539_ _0868_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ _1071_ _1172_ _1214_ _0922_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__o221a_1
X_2511_ PC.i_mem_addr\[2\] _0553_ _0542_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2373_ _0426_ _0619_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__mux2_1
X_1324_ _0622_ _0624_ ByteBuffer.instr\[19\] _0619_ vssd1 vssd1 vccd1 vccd1 _0667_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1942_ _1146_ _1274_ _0175_ _1161_ _0179_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1873_ _1066_ _1165_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2356_ _0436_ ALU.immediate\[9\] _0407_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__mux2_1
X_2287_ RegFile.A\[6\] net1 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__and2_1
X_1307_ _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2454__53 clknet_1_0__leaf__0517_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__inv_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _0390_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2072_ RegFile.D\[7\] _1184_ _0289_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2141_ _1183_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1925_ _1227_ _1249_ _1263_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__a211o_4
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1856_ _0632_ _1197_ _1198_ _0663_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1787_ _0960_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__xnor2_1
X_2339_ _0480_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1572_ RegFile.C\[4\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__and4_1
X_1710_ _0991_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__inv_2
X_2690_ clknet_2_2__leaf_clk _0167_ net58 vssd1 vssd1 vccd1 vccd1 PC.i_mem_addr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1641_ _0960_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__nor2_1
X_2124_ _0264_ RegFile.L\[7\] _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__mux2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _0277_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1908_ _1248_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1839_ _1126_ _1152_ _1180_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__o31a_2
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 gpo[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1624_ ALU.flags_to_alu\[6\] _0687_ _0683_ RegFile.E\[6\] _0654_ vssd1 vssd1 vccd1
+ vccd1 _0967_ sky130_fd_sc_hd__a221o_1
X_1555_ RegFile.L\[0\] _0770_ _0771_ RegFile.B\[0\] _0897_ vssd1 vssd1 vccd1 vccd1
+ _0898_ sky130_fd_sc_hd__a221o_1
X_2673_ net127 _0150_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.A\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2107_ _1184_ RegFile.H\[7\] _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__mux2_1
X_1486_ _0654_ _0823_ _0824_ _0827_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__a311o_2
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2038_ _1182_ _0262_ _0263_ net10 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1340_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2656_ net110 _0133_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.D\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1607_ RegFile.C\[7\] _0793_ _0786_ RegFile.D\[7\] vssd1 vssd1 vccd1 vccd1 _0950_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1469_ _0809_ _0810_ _0811_ _0774_ RegFile.A\[2\] vssd1 vssd1 vccd1 vccd1 _0812_
+ sky130_fd_sc_hd__o32a_1
X_2587_ PC.i_mem_addr\[15\] _0616_ _0542_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__mux2_1
X_1538_ _0869_ _0880_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ _0549_ _0552_ net47 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1323_ _0633_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__or2_2
X_2372_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2639_ net93 _0116_ net62 vssd1 vssd1 vccd1 vccd1 RegFile.H\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1941_ _1113_ _1210_ _0178_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1872_ _1122_ _1163_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__or2_2
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1306_ _0620_ _0647_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__and3_1
X_2355_ _0487_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
X_2286_ _0451_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _0630_ _1094_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2071_ _0287_ _0288_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nor2_4
X_1855_ ByteBuffer.instr\[19\] _0660_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nand2_1
X_1924_ _0937_ _1114_ _1116_ _1124_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1786_ _1100_ _1128_ _1070_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2338_ _0724_ _0476_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__and2_1
X_2269_ _0442_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__inv_6
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1571_ RegFile.E\[4\] _0761_ _0763_ RegFile.H\[4\] vssd1 vssd1 vccd1 vccd1 _0914_
+ sky130_fd_sc_hd__a22o_1
X_1640_ _0970_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__xnor2_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0268_ _0307_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__nand2_8
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ RegFile.C\[4\] _0276_ _0270_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__mux2_1
X_2409__10 clknet_1_0__leaf__0515_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__inv_2
X_1907_ RegFile.A\[5\] _1247_ _1203_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1838_ _1130_ _1166_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand2_1
X_1769_ _1107_ _1111_ _0832_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpo[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpo[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2672_ net126 _0149_ net63 vssd1 vssd1 vccd1 vccd1 RegFile.B\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1623_ _0961_ _0963_ _0964_ net51 _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a32o_1
X_1554_ RegFile.C\[0\] _0638_ _0681_ _0760_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__and4_1
X_1485_ _0664_ _0692_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__or2_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

