// This is the unpowered netlist.
module top8227 (M10ClkOut,
    clk,
    dataBusEnable,
    dataBusSelect,
    functionalClockOut,
    interruptRequest,
    nonMaskableInterrupt,
    nrst,
    readNotWrite,
    ready,
    setOverflow,
    sync,
    addressBusHigh,
    addressBusLow,
    dataBusInput,
    dataBusOutput);
 output M10ClkOut;
 input clk;
 input dataBusEnable;
 output dataBusSelect;
 output functionalClockOut;
 input interruptRequest;
 input nonMaskableInterrupt;
 input nrst;
 output readNotWrite;
 input ready;
 input setOverflow;
 output sync;
 output [7:0] addressBusHigh;
 output [7:0] addressBusLow;
 input [7:0] dataBusInput;
 output [7:0] dataBusOutput;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire \branch_ff.branchBackward ;
 wire \branch_ff.branchForward ;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \demux.PSR_C ;
 wire \demux.PSR_N ;
 wire \demux.PSR_V ;
 wire \demux.PSR_Z ;
 wire \demux.isAddressing ;
 wire \demux.nmi ;
 wire \demux.reset ;
 wire \demux.setInterruptFlag ;
 wire \demux.state_machine.currentAddress[0] ;
 wire \demux.state_machine.currentAddress[10] ;
 wire \demux.state_machine.currentAddress[11] ;
 wire \demux.state_machine.currentAddress[12] ;
 wire \demux.state_machine.currentAddress[1] ;
 wire \demux.state_machine.currentAddress[2] ;
 wire \demux.state_machine.currentAddress[3] ;
 wire \demux.state_machine.currentAddress[4] ;
 wire \demux.state_machine.currentAddress[5] ;
 wire \demux.state_machine.currentAddress[6] ;
 wire \demux.state_machine.currentAddress[7] ;
 wire \demux.state_machine.currentAddress[8] ;
 wire \demux.state_machine.currentAddress[9] ;
 wire \demux.state_machine.currentInstruction[0] ;
 wire \demux.state_machine.currentInstruction[1] ;
 wire \demux.state_machine.currentInstruction[2] ;
 wire \demux.state_machine.currentInstruction[3] ;
 wire \demux.state_machine.currentInstruction[4] ;
 wire \demux.state_machine.currentInstruction[5] ;
 wire \demux.state_machine.timeState[0] ;
 wire \demux.state_machine.timeState[1] ;
 wire \demux.state_machine.timeState[2] ;
 wire \demux.state_machine.timeState[3] ;
 wire \demux.state_machine.timeState[4] ;
 wire \demux.state_machine.timeState[5] ;
 wire \demux.state_machine.timeState[6] ;
 wire \free_carry_ff.freeCarry ;
 wire \instructionLoader.interruptInjector.interruptRequest ;
 wire \instructionLoader.interruptInjector.irqGenerated ;
 wire \instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ;
 wire \instructionLoader.interruptInjector.irqSync.nextQ2 ;
 wire \instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ;
 wire \instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ;
 wire \instructionLoader.interruptInjector.nmiSync.in ;
 wire \instructionLoader.interruptInjector.nmiSync.nextQ2 ;
 wire \instructionLoader.interruptInjector.processStatusRegIFlag ;
 wire \instructionLoader.interruptInjector.resetDetected ;
 wire \internalDataflow.accRegToDB[0] ;
 wire \internalDataflow.accRegToDB[1] ;
 wire \internalDataflow.accRegToDB[2] ;
 wire \internalDataflow.accRegToDB[3] ;
 wire \internalDataflow.accRegToDB[4] ;
 wire \internalDataflow.accRegToDB[5] ;
 wire \internalDataflow.accRegToDB[6] ;
 wire \internalDataflow.accRegToDB[7] ;
 wire \internalDataflow.addressHighBusModule.busInputs[16] ;
 wire \internalDataflow.addressHighBusModule.busInputs[17] ;
 wire \internalDataflow.addressHighBusModule.busInputs[18] ;
 wire \internalDataflow.addressHighBusModule.busInputs[19] ;
 wire \internalDataflow.addressHighBusModule.busInputs[20] ;
 wire \internalDataflow.addressHighBusModule.busInputs[21] ;
 wire \internalDataflow.addressHighBusModule.busInputs[22] ;
 wire \internalDataflow.addressHighBusModule.busInputs[23] ;
 wire \internalDataflow.addressLowBusModule.busInputs[16] ;
 wire \internalDataflow.addressLowBusModule.busInputs[17] ;
 wire \internalDataflow.addressLowBusModule.busInputs[18] ;
 wire \internalDataflow.addressLowBusModule.busInputs[19] ;
 wire \internalDataflow.addressLowBusModule.busInputs[20] ;
 wire \internalDataflow.addressLowBusModule.busInputs[21] ;
 wire \internalDataflow.addressLowBusModule.busInputs[22] ;
 wire \internalDataflow.addressLowBusModule.busInputs[23] ;
 wire \internalDataflow.addressLowBusModule.busInputs[24] ;
 wire \internalDataflow.addressLowBusModule.busInputs[25] ;
 wire \internalDataflow.addressLowBusModule.busInputs[26] ;
 wire \internalDataflow.addressLowBusModule.busInputs[27] ;
 wire \internalDataflow.addressLowBusModule.busInputs[28] ;
 wire \internalDataflow.addressLowBusModule.busInputs[29] ;
 wire \internalDataflow.addressLowBusModule.busInputs[30] ;
 wire \internalDataflow.addressLowBusModule.busInputs[31] ;
 wire \internalDataflow.addressLowBusModule.busInputs[32] ;
 wire \internalDataflow.addressLowBusModule.busInputs[33] ;
 wire \internalDataflow.addressLowBusModule.busInputs[34] ;
 wire \internalDataflow.addressLowBusModule.busInputs[35] ;
 wire \internalDataflow.addressLowBusModule.busInputs[36] ;
 wire \internalDataflow.addressLowBusModule.busInputs[37] ;
 wire \internalDataflow.addressLowBusModule.busInputs[38] ;
 wire \internalDataflow.addressLowBusModule.busInputs[39] ;
 wire \internalDataflow.dataBusModule.busInputs[43] ;
 wire \internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ;
 wire \internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ;
 wire \internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ;
 wire \internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ;
 wire \internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ;
 wire \internalDataflow.stackBusModule.busInputs[32] ;
 wire \internalDataflow.stackBusModule.busInputs[33] ;
 wire \internalDataflow.stackBusModule.busInputs[34] ;
 wire \internalDataflow.stackBusModule.busInputs[35] ;
 wire \internalDataflow.stackBusModule.busInputs[36] ;
 wire \internalDataflow.stackBusModule.busInputs[37] ;
 wire \internalDataflow.stackBusModule.busInputs[38] ;
 wire \internalDataflow.stackBusModule.busInputs[39] ;
 wire \internalDataflow.stackBusModule.busInputs[40] ;
 wire \internalDataflow.stackBusModule.busInputs[41] ;
 wire \internalDataflow.stackBusModule.busInputs[42] ;
 wire \internalDataflow.stackBusModule.busInputs[43] ;
 wire \internalDataflow.stackBusModule.busInputs[44] ;
 wire \internalDataflow.stackBusModule.busInputs[45] ;
 wire \internalDataflow.stackBusModule.busInputs[46] ;
 wire \internalDataflow.stackBusModule.busInputs[47] ;
 wire \negEdgeDetector.q1 ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \pulse_slower.currentEnableState[0] ;
 wire \pulse_slower.currentEnableState[1] ;
 wire \pulse_slower.nextEnableState[0] ;
 wire \pulse_slower.nextEnableState[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0968_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__clkbuf_2 _1503_ (.A(\demux.state_machine.currentInstruction[2] ),
    .X(_0810_));
 sky130_fd_sc_hd__buf_2 _1504_ (.A(\demux.state_machine.currentInstruction[3] ),
    .X(_0811_));
 sky130_fd_sc_hd__buf_2 _1505_ (.A(\demux.state_machine.currentInstruction[1] ),
    .X(_0812_));
 sky130_fd_sc_hd__clkbuf_2 _1506_ (.A(\demux.state_machine.currentInstruction[0] ),
    .X(_0813_));
 sky130_fd_sc_hd__or4bb_1 _1507_ (.A(_0810_),
    .B(_0811_),
    .C_N(_0812_),
    .D_N(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__buf_4 _1508_ (.A(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__or4_2 _1509_ (.A(_0812_),
    .B(_0813_),
    .C(_0810_),
    .D(_0811_),
    .X(_0816_));
 sky130_fd_sc_hd__or4b_1 _1510_ (.A(\demux.state_machine.currentInstruction[0] ),
    .B(\demux.state_machine.currentInstruction[2] ),
    .C(\demux.state_machine.currentInstruction[3] ),
    .D_N(\demux.state_machine.currentInstruction[1] ),
    .X(_0817_));
 sky130_fd_sc_hd__buf_4 _1511_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__buf_4 _1512_ (.A(\demux.state_machine.currentInstruction[5] ),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _1513_ (.A(\demux.state_machine.currentInstruction[4] ),
    .X(_0820_));
 sky130_fd_sc_hd__nand2_4 _1514_ (.A(_0819_),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__a31o_2 _1515_ (.A1(_0815_),
    .A2(_0816_),
    .A3(_0818_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__inv_2 _1516_ (.A(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__or4b_1 _1517_ (.A(_0812_),
    .B(_0813_),
    .C(_0811_),
    .D_N(_0810_),
    .X(_0824_));
 sky130_fd_sc_hd__buf_4 _1518_ (.A(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nand2b_4 _1519_ (.A_N(\demux.state_machine.currentInstruction[5] ),
    .B(_0820_),
    .Y(_0826_));
 sky130_fd_sc_hd__buf_4 _1520_ (.A(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__a21oi_1 _1521_ (.A1(_0815_),
    .A2(_0825_),
    .B1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2b_4 _1522_ (.A_N(\demux.state_machine.currentInstruction[4] ),
    .B(_0819_),
    .Y(_0829_));
 sky130_fd_sc_hd__clkbuf_8 _1523_ (.A(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_2 _1524_ (.A(_0830_),
    .B(_0816_),
    .Y(_0831_));
 sky130_fd_sc_hd__clkbuf_4 _1525_ (.A(_0812_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_4 _1526_ (.A(_0813_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_4 _1527_ (.A(_0810_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_4 _1528_ (.A(_0811_),
    .X(_0835_));
 sky130_fd_sc_hd__nand4_4 _1529_ (.A(_0832_),
    .B(_0833_),
    .C(_0834_),
    .D(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__nor2_1 _1530_ (.A(_0827_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand4b_2 _1531_ (.A_N(_0833_),
    .B(_0834_),
    .C(_0835_),
    .D(_0832_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_2 _1532_ (.A(_0827_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__or3_2 _1533_ (.A(_0831_),
    .B(_0837_),
    .C(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__or2_2 _1534_ (.A(\demux.state_machine.currentInstruction[5] ),
    .B(\demux.state_machine.currentInstruction[4] ),
    .X(_0841_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(_0841_),
    .B(_0836_),
    .Y(_0842_));
 sky130_fd_sc_hd__or4b_1 _1536_ (.A(\demux.state_machine.currentInstruction[1] ),
    .B(\demux.state_machine.currentInstruction[2] ),
    .C(\demux.state_machine.currentInstruction[3] ),
    .D_N(\demux.state_machine.currentInstruction[0] ),
    .X(_0843_));
 sky130_fd_sc_hd__clkbuf_4 _1537_ (.A(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__nor2_1 _1538_ (.A(_0826_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nor2_1 _1539_ (.A(_0826_),
    .B(_0816_),
    .Y(_0846_));
 sky130_fd_sc_hd__nor2_4 _1540_ (.A(_0826_),
    .B(_0818_),
    .Y(_0847_));
 sky130_fd_sc_hd__or4_2 _1541_ (.A(_0842_),
    .B(_0845_),
    .C(_0846_),
    .D(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__or4_1 _1542_ (.A(_0823_),
    .B(_0828_),
    .C(_0840_),
    .D(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_0830_),
    .B(_0836_),
    .Y(_0850_));
 sky130_fd_sc_hd__or4bb_1 _1544_ (.A(_0812_),
    .B(_0813_),
    .C_N(_0810_),
    .D_N(_0811_),
    .X(_0851_));
 sky130_fd_sc_hd__buf_4 _1545_ (.A(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _1546_ (.A(_0821_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__or4bb_1 _1547_ (.A(\demux.state_machine.currentInstruction[1] ),
    .B(_0811_),
    .C_N(_0810_),
    .D_N(_0813_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_4 _1548_ (.A(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__a21oi_1 _1549_ (.A1(_0855_),
    .A2(_0825_),
    .B1(_0821_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand4b_4 _1550_ (.A_N(_0812_),
    .B(_0833_),
    .C(_0834_),
    .D(_0835_),
    .Y(_0857_));
 sky130_fd_sc_hd__or2b_1 _1551_ (.A(_0834_),
    .B_N(_0835_),
    .X(_0858_));
 sky130_fd_sc_hd__or4bb_1 _1552_ (.A(_0813_),
    .B(_0811_),
    .C_N(_0810_),
    .D_N(_0812_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_4 _1553_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nand4b_4 _1554_ (.A_N(_0835_),
    .B(_0834_),
    .C(_0833_),
    .D(_0832_),
    .Y(_0861_));
 sky130_fd_sc_hd__a41o_1 _1555_ (.A1(_0857_),
    .A2(_0858_),
    .A3(_0860_),
    .A4(_0861_),
    .B1(_0821_),
    .X(_0862_));
 sky130_fd_sc_hd__or4b_1 _1556_ (.A(_0850_),
    .B(_0853_),
    .C(_0856_),
    .D_N(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__or4bb_1 _1557_ (.A(_0813_),
    .B(_0810_),
    .C_N(_0811_),
    .D_N(_0812_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_8 _1558_ (.A(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__buf_4 _1559_ (.A(_0827_),
    .X(_0866_));
 sky130_fd_sc_hd__a21oi_2 _1560_ (.A1(_0865_),
    .A2(_0860_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nor2_4 _1561_ (.A(_0829_),
    .B(_0852_),
    .Y(_0868_));
 sky130_fd_sc_hd__clkbuf_4 _1562_ (.A(_0841_),
    .X(_0869_));
 sky130_fd_sc_hd__a21oi_2 _1563_ (.A1(_0844_),
    .A2(_0818_),
    .B1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__buf_4 _1564_ (.A(_0830_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(_0871_),
    .B(_0818_),
    .Y(_0872_));
 sky130_fd_sc_hd__nor2_4 _1566_ (.A(_0869_),
    .B(_0861_),
    .Y(_0873_));
 sky130_fd_sc_hd__or4_1 _1567_ (.A(_0868_),
    .B(_0870_),
    .C(_0872_),
    .D(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_4 _1568_ (.A(\demux.state_machine.timeState[4] ),
    .X(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _1569_ (.A(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _1570_ (.A(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__o41a_1 _1571_ (.A1(_0849_),
    .A2(_0863_),
    .A3(_0867_),
    .A4(_0874_),
    .B1(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_4 _1572_ (.A(\demux.state_machine.timeState[6] ),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _1573_ (.A(_0869_),
    .B(_0865_),
    .X(_0880_));
 sky130_fd_sc_hd__or4b_1 _1574_ (.A(\demux.state_machine.currentInstruction[1] ),
    .B(_0813_),
    .C(\demux.state_machine.currentInstruction[2] ),
    .D_N(\demux.state_machine.currentInstruction[3] ),
    .X(_0881_));
 sky130_fd_sc_hd__buf_4 _1575_ (.A(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__or4b_1 _1576_ (.A(_0819_),
    .B(_0882_),
    .C(_0820_),
    .D_N(\demux.PSR_N ),
    .X(_0883_));
 sky130_fd_sc_hd__or4bb_1 _1577_ (.A(_0812_),
    .B(_0810_),
    .C_N(_0811_),
    .D_N(_0813_),
    .X(_0884_));
 sky130_fd_sc_hd__clkbuf_4 _1578_ (.A(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__or3_1 _1579_ (.A(\demux.PSR_Z ),
    .B(_0869_),
    .C(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or4b_1 _1580_ (.A(_0819_),
    .B(_0855_),
    .C(_0820_),
    .D_N(\demux.PSR_C ),
    .X(_0887_));
 sky130_fd_sc_hd__o2111a_2 _1581_ (.A1(\demux.PSR_N ),
    .A2(_0880_),
    .B1(_0883_),
    .C1(_0886_),
    .D1(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_1 _1582_ (.A(_0869_),
    .B(_0860_),
    .Y(_0889_));
 sky130_fd_sc_hd__and4b_1 _1583_ (.A_N(_0832_),
    .B(_0833_),
    .C(_0834_),
    .D(_0835_),
    .X(_0890_));
 sky130_fd_sc_hd__nor2_4 _1584_ (.A(_0819_),
    .B(_0820_),
    .Y(_0891_));
 sky130_fd_sc_hd__and3_1 _1585_ (.A(\demux.PSR_V ),
    .B(_0890_),
    .C(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__nor3_1 _1586_ (.A(\demux.PSR_C ),
    .B(_0869_),
    .C(_0825_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor3_1 _1587_ (.A(\demux.PSR_V ),
    .B(_0869_),
    .C(_0852_),
    .Y(_0894_));
 sky130_fd_sc_hd__a2111oi_1 _1588_ (.A1(\demux.PSR_Z ),
    .A2(_0889_),
    .B1(_0892_),
    .C1(_0893_),
    .D1(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__buf_2 _1589_ (.A(\demux.state_machine.timeState[2] ),
    .X(_0896_));
 sky130_fd_sc_hd__buf_4 _1590_ (.A(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_1 _1591_ (.A(\branch_ff.branchForward ),
    .B(\branch_ff.branchBackward ),
    .Y(_0898_));
 sky130_fd_sc_hd__and2_1 _1592_ (.A(_0897_),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__a31o_1 _1593_ (.A1(_0877_),
    .A2(_0888_),
    .A3(net53),
    .B1(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__buf_4 _1594_ (.A(_0869_),
    .X(_0901_));
 sky130_fd_sc_hd__a41o_1 _1595_ (.A1(_0857_),
    .A2(_0882_),
    .A3(_0825_),
    .A4(_0865_),
    .B1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a41o_1 _1596_ (.A1(_0885_),
    .A2(_0855_),
    .A3(_0860_),
    .A4(_0852_),
    .B1(_0901_),
    .X(_0903_));
 sky130_fd_sc_hd__nand2_2 _1597_ (.A(_0902_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__clkbuf_4 _1598_ (.A(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__o21a_1 _1599_ (.A1(_0879_),
    .A2(_0900_),
    .B1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nor2_1 _1600_ (.A(_0857_),
    .B(_0829_),
    .Y(_0907_));
 sky130_fd_sc_hd__nor2_1 _1601_ (.A(_0829_),
    .B(_0838_),
    .Y(_0908_));
 sky130_fd_sc_hd__nand4b_4 _1602_ (.A_N(_0810_),
    .B(_0811_),
    .C(_0812_),
    .D(_0833_),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_4 _1603_ (.A(_0826_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__or3_2 _1604_ (.A(_0907_),
    .B(_0908_),
    .C(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__nor2_4 _1605_ (.A(_0826_),
    .B(_0857_),
    .Y(_0912_));
 sky130_fd_sc_hd__a21oi_4 _1606_ (.A1(_0909_),
    .A2(_0865_),
    .B1(_0871_),
    .Y(_0913_));
 sky130_fd_sc_hd__o21a_1 _1607_ (.A1(_0912_),
    .A2(_0913_),
    .B1(\demux.state_machine.timeState[5] ),
    .X(_0914_));
 sky130_fd_sc_hd__a21oi_2 _1608_ (.A1(_0882_),
    .A2(_0861_),
    .B1(_0866_),
    .Y(_0915_));
 sky130_fd_sc_hd__and4bb_1 _1609_ (.A_N(_0820_),
    .B_N(_0825_),
    .C(_0896_),
    .D(_0819_),
    .X(_0916_));
 sky130_fd_sc_hd__inv_2 _1610_ (.A(\demux.state_machine.timeState[4] ),
    .Y(_0917_));
 sky130_fd_sc_hd__nor3_1 _1611_ (.A(_0917_),
    .B(_0871_),
    .C(_0815_),
    .Y(_0918_));
 sky130_fd_sc_hd__a211o_1 _1612_ (.A1(_0876_),
    .A2(_0915_),
    .B1(_0916_),
    .C1(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__nor2_2 _1613_ (.A(_0869_),
    .B(_0909_),
    .Y(_0920_));
 sky130_fd_sc_hd__nor2_2 _1614_ (.A(_0869_),
    .B(_0838_),
    .Y(_0921_));
 sky130_fd_sc_hd__a22o_1 _1615_ (.A1(\demux.state_machine.timeState[3] ),
    .A2(_0920_),
    .B1(_0921_),
    .B2(_0875_),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_1 _1616_ (.A(_0871_),
    .B(_0855_),
    .Y(_0923_));
 sky130_fd_sc_hd__and2_1 _1617_ (.A(_0897_),
    .B(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__or4_1 _1618_ (.A(_0914_),
    .B(_0919_),
    .C(_0922_),
    .D(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a31oi_2 _1619_ (.A1(_0885_),
    .A2(_0844_),
    .A3(_0882_),
    .B1(_0830_),
    .Y(_0926_));
 sky130_fd_sc_hd__nor2_4 _1620_ (.A(_0841_),
    .B(_0815_),
    .Y(_0927_));
 sky130_fd_sc_hd__a21o_1 _1621_ (.A1(_0885_),
    .A2(_0855_),
    .B1(_0866_),
    .X(_0928_));
 sky130_fd_sc_hd__or3b_1 _1622_ (.A(_0926_),
    .B(_0927_),
    .C_N(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__a21oi_4 _1623_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0830_),
    .Y(_0930_));
 sky130_fd_sc_hd__o21a_1 _1624_ (.A1(_0929_),
    .A2(_0930_),
    .B1(_0879_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_4 _1625_ (.A(\demux.state_machine.timeState[0] ),
    .X(_0932_));
 sky130_fd_sc_hd__nor2_2 _1626_ (.A(_0827_),
    .B(_0852_),
    .Y(_0933_));
 sky130_fd_sc_hd__and2_1 _1627_ (.A(_0932_),
    .B(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__a2111o_1 _1628_ (.A1(_0877_),
    .A2(_0911_),
    .B1(_0925_),
    .C1(_0931_),
    .D1(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__or2_4 _1629_ (.A(_0896_),
    .B(\demux.state_machine.timeState[6] ),
    .X(_0936_));
 sky130_fd_sc_hd__nor2_1 _1630_ (.A(\demux.state_machine.timeState[2] ),
    .B(\demux.state_machine.timeState[6] ),
    .Y(_0937_));
 sky130_fd_sc_hd__a21oi_1 _1631_ (.A1(_0917_),
    .A2(_0937_),
    .B1(\demux.reset ),
    .Y(_0938_));
 sky130_fd_sc_hd__and2b_2 _1632_ (.A_N(_0820_),
    .B(_0819_),
    .X(_0939_));
 sky130_fd_sc_hd__and2b_1 _1633_ (.A_N(_0835_),
    .B(_0834_),
    .X(_0940_));
 sky130_fd_sc_hd__and4b_2 _1634_ (.A_N(_0832_),
    .B(_0939_),
    .C(_0940_),
    .D(\demux.state_machine.timeState[4] ),
    .X(_0941_));
 sky130_fd_sc_hd__a221oi_2 _1635_ (.A1(_0912_),
    .A2(_0936_),
    .B1(_0920_),
    .B2(_0938_),
    .C1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(_0827_),
    .B(_0885_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2_2 _1637_ (.A(_0827_),
    .B(_0855_),
    .Y(_0944_));
 sky130_fd_sc_hd__or2_2 _1638_ (.A(_0896_),
    .B(\demux.state_machine.timeState[4] ),
    .X(_0945_));
 sky130_fd_sc_hd__o41ai_2 _1639_ (.A1(_0926_),
    .A2(_0943_),
    .A3(_0944_),
    .A4(_0927_),
    .B1(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__nor4_2 _1640_ (.A(\demux.state_machine.currentAddress[8] ),
    .B(\demux.state_machine.currentAddress[0] ),
    .C(\demux.state_machine.currentAddress[2] ),
    .D(\demux.state_machine.currentAddress[9] ),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_4 _1641_ (.A(\demux.isAddressing ),
    .B(net56),
    .Y(_0948_));
 sky130_fd_sc_hd__o21ai_2 _1642_ (.A1(_0932_),
    .A2(_0822_),
    .B1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__a31oi_4 _1643_ (.A1(_0942_),
    .A2(_0946_),
    .A3(_0822_),
    .B1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__or2_2 _1644_ (.A(\pulse_slower.currentEnableState[1] ),
    .B(\pulse_slower.currentEnableState[0] ),
    .X(_0951_));
 sky130_fd_sc_hd__inv_2 _1645_ (.A(_0951_),
    .Y(\pulse_slower.nextEnableState[0] ));
 sky130_fd_sc_hd__o211a_1 _1646_ (.A1(net13),
    .A2(_0950_),
    .B1(\pulse_slower.nextEnableState[0] ),
    .C1(_0948_),
    .X(_0952_));
 sky130_fd_sc_hd__o31a_1 _1647_ (.A1(_0878_),
    .A2(_0906_),
    .A3(_0935_),
    .B1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_2 _1648_ (.A(_0953_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 _1649_ (.A(net6),
    .X(_0954_));
 sky130_fd_sc_hd__nor3_1 _1650_ (.A(\demux.nmi ),
    .B(\instructionLoader.interruptInjector.resetDetected ),
    .C(\instructionLoader.interruptInjector.irqGenerated ),
    .Y(_0955_));
 sky130_fd_sc_hd__clkbuf_4 _1651_ (.A(net55),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_4 _1652_ (.A(net5),
    .X(_0957_));
 sky130_fd_sc_hd__and4b_2 _1653_ (.A_N(_0954_),
    .B(_0956_),
    .C(net4),
    .D(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__inv_2 _1654_ (.A(net13),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(_0950_),
    .Y(net42));
 sky130_fd_sc_hd__a21o_2 _1656_ (.A1(_0959_),
    .A2(net42),
    .B1(_0951_),
    .X(_0960_));
 sky130_fd_sc_hd__buf_4 _1657_ (.A(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__nor2_2 _1658_ (.A(\instructionLoader.interruptInjector.resetDetected ),
    .B(net43),
    .Y(_0962_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(_0961_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__o21ai_4 _1660_ (.A1(net2),
    .A2(net3),
    .B1(_0956_),
    .Y(_0964_));
 sky130_fd_sc_hd__and2_1 _1661_ (.A(_0963_),
    .B(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__clkbuf_4 _1662_ (.A(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_4 _1663_ (.A(net7),
    .X(_0967_));
 sky130_fd_sc_hd__inv_2 _1664_ (.A(net9),
    .Y(_0968_));
 sky130_fd_sc_hd__buf_2 _1665_ (.A(net8),
    .X(_0969_));
 sky130_fd_sc_hd__and3_1 _1666_ (.A(_0968_),
    .B(_0969_),
    .C(_0956_),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _1667_ (.A(_0967_),
    .B(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__buf_2 _1668_ (.A(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_1 _1669_ (.A(_0961_),
    .B(_0962_),
    .X(_0973_));
 sky130_fd_sc_hd__buf_2 _1670_ (.A(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__buf_2 _1671_ (.A(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__buf_2 _1672_ (.A(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__clkbuf_4 _1673_ (.A(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a32o_1 _1674_ (.A1(_0958_),
    .A2(_0966_),
    .A3(_0972_),
    .B1(_0977_),
    .B2(\demux.state_machine.currentAddress[6] ),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _1675_ (.A(_0963_),
    .X(_0978_));
 sky130_fd_sc_hd__clkbuf_4 _1676_ (.A(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\demux.state_machine.currentAddress[7] ),
    .A1(_0958_),
    .S(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__a21boi_1 _1678_ (.A1(_0966_),
    .A2(_0972_),
    .B1_N(_0980_),
    .Y(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _1679_ (.A(_0961_),
    .X(_0981_));
 sky130_fd_sc_hd__buf_4 _1680_ (.A(_0948_),
    .X(_0982_));
 sky130_fd_sc_hd__clkbuf_4 _1681_ (.A(_0897_),
    .X(_0983_));
 sky130_fd_sc_hd__or2_1 _1682_ (.A(\demux.state_machine.currentAddress[4] ),
    .B(\demux.state_machine.currentAddress[10] ),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_4 _1683_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__nor2_1 _1684_ (.A(_0932_),
    .B(_0875_),
    .Y(_0986_));
 sky130_fd_sc_hd__clkbuf_4 _1685_ (.A(\demux.state_machine.currentAddress[1] ),
    .X(_0987_));
 sky130_fd_sc_hd__buf_2 _1686_ (.A(\demux.state_machine.currentAddress[12] ),
    .X(_0988_));
 sky130_fd_sc_hd__nor4b_1 _1687_ (.A(_0932_),
    .B(_0896_),
    .C(_0875_),
    .D_N(\demux.state_machine.timeState[6] ),
    .Y(_0989_));
 sky130_fd_sc_hd__o31a_1 _1688_ (.A1(_0987_),
    .A2(_0988_),
    .A3(\demux.state_machine.currentAddress[6] ),
    .B1(net54),
    .X(_0990_));
 sky130_fd_sc_hd__or3_2 _1689_ (.A(\demux.state_machine.currentAddress[11] ),
    .B(\demux.state_machine.currentAddress[3] ),
    .C(\demux.state_machine.currentAddress[7] ),
    .X(_0991_));
 sky130_fd_sc_hd__and2b_1 _1690_ (.A_N(\demux.state_machine.timeState[0] ),
    .B(\demux.state_machine.timeState[4] ),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_4 _1691_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__and2_1 _1692_ (.A(_0932_),
    .B(\demux.state_machine.currentAddress[5] ),
    .X(_0994_));
 sky130_fd_sc_hd__a21o_1 _1693_ (.A1(_0991_),
    .A2(_0993_),
    .B1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a311oi_2 _1694_ (.A1(_0983_),
    .A2(_0985_),
    .A3(_0986_),
    .B1(_0990_),
    .C1(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__a21oi_1 _1695_ (.A1(_0959_),
    .A2(net42),
    .B1(_0951_),
    .Y(_0997_));
 sky130_fd_sc_hd__clkbuf_4 _1696_ (.A(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__buf_4 _1697_ (.A(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__o211a_2 _1698_ (.A1(_0982_),
    .A2(_0996_),
    .B1(_0962_),
    .C1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__a22o_1 _1699_ (.A1(_0879_),
    .A2(_0981_),
    .B1(_1000_),
    .B2(_0983_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _1700_ (.A1(\demux.state_machine.timeState[5] ),
    .A2(_0981_),
    .B1(_1000_),
    .B2(\demux.state_machine.timeState[1] ),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _1701_ (.A(_0877_),
    .X(_1001_));
 sky130_fd_sc_hd__clkbuf_4 _1702_ (.A(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__buf_4 _1703_ (.A(_0932_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_4 _1704_ (.A(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_4 _1705_ (.A(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__buf_2 _1706_ (.A(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_4 _1707_ (.A(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_4 _1708_ (.A(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__a22o_1 _1709_ (.A1(_1002_),
    .A2(_0981_),
    .B1(_1000_),
    .B2(_1008_),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _1710_ (.A1(net84),
    .A2(_0981_),
    .B1(_1000_),
    .B2(\demux.state_machine.timeState[5] ),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _1711_ (.A1(_0983_),
    .A2(_0981_),
    .B1(_1000_),
    .B2(_1002_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _1712_ (.A1(\demux.state_machine.timeState[1] ),
    .A2(_0981_),
    .B1(_1000_),
    .B2(_0879_),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _1713_ (.A(_1000_),
    .Y(_1009_));
 sky130_fd_sc_hd__o22a_1 _1714_ (.A1(_1008_),
    .A2(_0999_),
    .B1(_1009_),
    .B2(net84),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _1715_ (.A(_0956_),
    .X(_1010_));
 sky130_fd_sc_hd__and4b_1 _1716_ (.A_N(_0957_),
    .B(_0954_),
    .C(_1010_),
    .D(net4),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_4 _1717_ (.A(net9),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_2 _1718_ (.A(_1012_),
    .B(net55),
    .Y(_1013_));
 sky130_fd_sc_hd__nor2_1 _1719_ (.A(_0969_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__and3_1 _1720_ (.A(net3),
    .B(_0979_),
    .C(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _1721_ (.A1(net85),
    .A2(_0977_),
    .B1(_1011_),
    .B2(_1015_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_2 _1722_ (.A(net4),
    .B(_0957_),
    .X(_1016_));
 sky130_fd_sc_hd__o21ai_4 _1723_ (.A1(_0954_),
    .A2(_1016_),
    .B1(_0956_),
    .Y(_1017_));
 sky130_fd_sc_hd__and4b_1 _1724_ (.A_N(net3),
    .B(_0978_),
    .C(_1010_),
    .D(net2),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_4 _1725_ (.A(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__a22o_1 _1726_ (.A1(_0988_),
    .A2(_0977_),
    .B1(_1017_),
    .B2(_1019_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _1727_ (.A0(\demux.state_machine.currentAddress[11] ),
    .A1(_1011_),
    .S(_0979_),
    .X(_1020_));
 sky130_fd_sc_hd__and2b_1 _1728_ (.A_N(_1015_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _1729_ (.A(_1021_),
    .X(_0002_));
 sky130_fd_sc_hd__or3_4 _1730_ (.A(\demux.nmi ),
    .B(\instructionLoader.interruptInjector.resetDetected ),
    .C(\instructionLoader.interruptInjector.irqGenerated ),
    .X(_1022_));
 sky130_fd_sc_hd__or4b_2 _1731_ (.A(net4),
    .B(_0954_),
    .C(_1022_),
    .D_N(_0957_),
    .X(_1023_));
 sky130_fd_sc_hd__and4bb_2 _1732_ (.A_N(_0957_),
    .B_N(_0954_),
    .C(_0956_),
    .D(net4),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(_1013_),
    .B(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_2 _1734_ (.A(net3),
    .B(_0956_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21oi_1 _1735_ (.A1(_1023_),
    .A2(_1025_),
    .B1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__mux2_1 _1736_ (.A0(\demux.state_machine.currentAddress[0] ),
    .A1(_1027_),
    .S(_0979_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _1737_ (.A(_1028_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_1 _1738_ (.A(_0954_),
    .B(_0956_),
    .Y(_1029_));
 sky130_fd_sc_hd__nor2_1 _1739_ (.A(_1016_),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__a22o_1 _1740_ (.A1(_0987_),
    .A2(_0977_),
    .B1(_1019_),
    .B2(_1030_),
    .X(_0004_));
 sky130_fd_sc_hd__o211a_1 _1741_ (.A1(_1026_),
    .A2(_1014_),
    .B1(_1024_),
    .C1(_0979_),
    .X(_1031_));
 sky130_fd_sc_hd__a21o_1 _1742_ (.A1(net101),
    .A2(_0977_),
    .B1(_1031_),
    .X(_0008_));
 sky130_fd_sc_hd__and4_1 _1743_ (.A(net3),
    .B(_0963_),
    .C(_1010_),
    .D(_1017_),
    .X(_1032_));
 sky130_fd_sc_hd__inv_2 _1744_ (.A(_1013_),
    .Y(_1033_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(_0961_),
    .B(_1023_),
    .Y(_1034_));
 sky130_fd_sc_hd__a32o_1 _1746_ (.A1(_0966_),
    .A2(_1033_),
    .A3(_1017_),
    .B1(_1019_),
    .B2(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__a211o_1 _1747_ (.A1(net78),
    .A2(_0977_),
    .B1(_1032_),
    .C1(_1035_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _1748_ (.A(net4),
    .B(_0957_),
    .Y(_1036_));
 sky130_fd_sc_hd__o21a_1 _1749_ (.A1(_1026_),
    .A2(_1016_),
    .B1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o21ai_1 _1750_ (.A1(_1029_),
    .A2(_1037_),
    .B1(_0979_),
    .Y(_1038_));
 sky130_fd_sc_hd__o21a_1 _1751_ (.A1(net81),
    .A2(_0979_),
    .B1(_1038_),
    .X(_0007_));
 sky130_fd_sc_hd__inv_2 _1752_ (.A(net4),
    .Y(_1039_));
 sky130_fd_sc_hd__and3_1 _1753_ (.A(_1039_),
    .B(_0957_),
    .C(_0956_),
    .X(_1040_));
 sky130_fd_sc_hd__and2_2 _1754_ (.A(_0954_),
    .B(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(net86),
    .A2(_0977_),
    .B1(_1019_),
    .B2(_1041_),
    .X(_0001_));
 sky130_fd_sc_hd__a41o_1 _1756_ (.A1(_1012_),
    .A2(_0969_),
    .A3(_1010_),
    .A4(_1024_),
    .B1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__a21o_1 _1757_ (.A1(_1013_),
    .A2(_1017_),
    .B1(_1040_),
    .X(_1043_));
 sky130_fd_sc_hd__a32o_1 _1758_ (.A1(net3),
    .A2(_1010_),
    .A3(_1042_),
    .B1(_1043_),
    .B2(_0964_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _1759_ (.A0(net113),
    .A1(_1044_),
    .S(_0979_),
    .X(_1045_));
 sky130_fd_sc_hd__clkbuf_1 _1760_ (.A(_1045_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _1761_ (.A(_0963_),
    .B(_0964_),
    .C(_1030_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_4 _1762_ (.A(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__a21o_1 _1763_ (.A1(net76),
    .A2(_0977_),
    .B1(_1047_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_4 _1764_ (.A(_0978_),
    .B(_0964_),
    .C(_1041_),
    .X(_1048_));
 sky130_fd_sc_hd__nor2_1 _1765_ (.A(_0836_),
    .B(_0978_),
    .Y(_1049_));
 sky130_fd_sc_hd__a22o_1 _1766_ (.A1(_0972_),
    .A2(_1048_),
    .B1(_1049_),
    .B2(_0939_),
    .X(_1050_));
 sky130_fd_sc_hd__and2b_1 _1767_ (.A_N(_0819_),
    .B(_0820_),
    .X(_1051_));
 sky130_fd_sc_hd__nor2_2 _1768_ (.A(_0962_),
    .B(_1026_),
    .Y(_1052_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(_1017_),
    .B(_1040_),
    .Y(_1053_));
 sky130_fd_sc_hd__and3_2 _1770_ (.A(_0998_),
    .B(_1052_),
    .C(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__and2_2 _1771_ (.A(_0967_),
    .B(_1014_),
    .X(_1055_));
 sky130_fd_sc_hd__a221o_1 _1772_ (.A1(_1051_),
    .A2(_1049_),
    .B1(_1054_),
    .B2(_1055_),
    .C1(_1032_),
    .X(_1056_));
 sky130_fd_sc_hd__or2_1 _1773_ (.A(_1050_),
    .B(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__nor2_1 _1774_ (.A(_0821_),
    .B(_0861_),
    .Y(_1058_));
 sky130_fd_sc_hd__and2b_2 _1775_ (.A_N(_0967_),
    .B(_1014_),
    .X(_1059_));
 sky130_fd_sc_hd__and2_1 _1776_ (.A(_1052_),
    .B(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__a22o_1 _1777_ (.A1(_1058_),
    .A2(_0974_),
    .B1(_1034_),
    .B2(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__and4b_1 _1778_ (.A_N(_0967_),
    .B(_0969_),
    .C(net55),
    .D(_1012_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_2 _1779_ (.A(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__a22o_1 _1780_ (.A1(_0842_),
    .A2(_0975_),
    .B1(_1048_),
    .B2(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__or3_1 _1781_ (.A(_1057_),
    .B(_1061_),
    .C(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_4 _1782_ (.A(_0974_),
    .X(_1066_));
 sky130_fd_sc_hd__buf_2 _1783_ (.A(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__inv_2 _1784_ (.A(_0965_),
    .Y(_1068_));
 sky130_fd_sc_hd__nor2_4 _1785_ (.A(_1068_),
    .B(_1023_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22o_1 _1786_ (.A1(_0910_),
    .A2(_1067_),
    .B1(_1063_),
    .B2(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__nor2_4 _1787_ (.A(_0830_),
    .B(_0909_),
    .Y(_1071_));
 sky130_fd_sc_hd__a32o_1 _1788_ (.A1(_0966_),
    .A2(_0972_),
    .A3(_1017_),
    .B1(_1067_),
    .B2(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__or2_1 _1789_ (.A(_1070_),
    .B(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a211o_1 _1790_ (.A1(_0957_),
    .A2(_0954_),
    .B1(_1022_),
    .C1(_1039_),
    .X(_1074_));
 sky130_fd_sc_hd__inv_2 _1791_ (.A(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__clkbuf_4 _1792_ (.A(_0821_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_2 _1793_ (.A(_0815_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__a32o_1 _1794_ (.A1(_0966_),
    .A2(_1059_),
    .A3(_1075_),
    .B1(_1067_),
    .B2(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_4 _1795_ (.A(_0920_),
    .X(_1079_));
 sky130_fd_sc_hd__o21ai_1 _1796_ (.A1(_1012_),
    .A2(_0969_),
    .B1(_1010_),
    .Y(_1080_));
 sky130_fd_sc_hd__a21boi_4 _1797_ (.A1(_0967_),
    .A2(_1010_),
    .B1_N(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__a31o_1 _1798_ (.A1(_0964_),
    .A2(_1017_),
    .A3(_1081_),
    .B1(_1066_),
    .X(_1082_));
 sky130_fd_sc_hd__o21a_1 _1799_ (.A1(_1079_),
    .A2(_0978_),
    .B1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__and4b_4 _1800_ (.A_N(_0834_),
    .B(_0835_),
    .C(_0832_),
    .D(_0833_),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _1801_ (.A(_0819_),
    .B(_0820_),
    .X(_1085_));
 sky130_fd_sc_hd__or3b_1 _1802_ (.A(_1022_),
    .B(_1012_),
    .C_N(_0969_),
    .X(_1086_));
 sky130_fd_sc_hd__nor2_2 _1803_ (.A(_0967_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__and2_2 _1804_ (.A(_1034_),
    .B(_1052_),
    .X(_1088_));
 sky130_fd_sc_hd__a32o_1 _1805_ (.A1(_1084_),
    .A2(_1085_),
    .A3(_0975_),
    .B1(_1087_),
    .B2(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__a21o_1 _1806_ (.A1(_0967_),
    .A2(_0958_),
    .B1(_1024_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_4 _1807_ (.A(_1066_),
    .X(_1091_));
 sky130_fd_sc_hd__a32o_1 _1808_ (.A1(_0966_),
    .A2(_1080_),
    .A3(_1090_),
    .B1(_1091_),
    .B2(_0873_),
    .X(_1092_));
 sky130_fd_sc_hd__or4_1 _1809_ (.A(_1078_),
    .B(_1083_),
    .C(_1089_),
    .D(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__nor2_2 _1810_ (.A(_0871_),
    .B(_0861_),
    .Y(_1094_));
 sky130_fd_sc_hd__and4bb_4 _1811_ (.A_N(_1012_),
    .B_N(_0969_),
    .C(net55),
    .D(_0967_),
    .X(_1095_));
 sky130_fd_sc_hd__a22o_1 _1812_ (.A1(_1094_),
    .A2(_0975_),
    .B1(_1069_),
    .B2(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nor2_2 _1813_ (.A(_0866_),
    .B(_0861_),
    .Y(_1097_));
 sky130_fd_sc_hd__a22o_1 _1814_ (.A1(_1097_),
    .A2(_1067_),
    .B1(_1059_),
    .B2(_1069_),
    .X(_1098_));
 sky130_fd_sc_hd__or2_1 _1815_ (.A(_1096_),
    .B(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__or4_1 _1816_ (.A(_1065_),
    .B(_1073_),
    .C(_1093_),
    .D(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__a22o_1 _1817_ (.A1(_0907_),
    .A2(_0975_),
    .B1(_1048_),
    .B2(_1095_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_4 _1818_ (.A(_0912_),
    .X(_1102_));
 sky130_fd_sc_hd__a31o_1 _1819_ (.A1(_0964_),
    .A2(_1017_),
    .A3(_1095_),
    .B1(_0974_),
    .X(_1103_));
 sky130_fd_sc_hd__o21a_1 _1820_ (.A1(_1102_),
    .A2(_0978_),
    .B1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a31o_1 _1821_ (.A1(_0890_),
    .A2(_0891_),
    .A3(_0976_),
    .B1(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__a211o_1 _1822_ (.A1(_0972_),
    .A2(_1047_),
    .B1(_1101_),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _1823_ (.A1(_0944_),
    .A2(_1067_),
    .B1(_1054_),
    .B2(_1063_),
    .X(_1107_));
 sky130_fd_sc_hd__nor2_1 _1824_ (.A(_0855_),
    .B(_1076_),
    .Y(_1108_));
 sky130_fd_sc_hd__a22o_1 _1825_ (.A1(_1108_),
    .A2(_1067_),
    .B1(_1055_),
    .B2(_1069_),
    .X(_1109_));
 sky130_fd_sc_hd__a221o_1 _1826_ (.A1(_0923_),
    .A2(_0976_),
    .B1(_1069_),
    .B2(_1081_),
    .C1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__or3_1 _1827_ (.A(_1106_),
    .B(_1107_),
    .C(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__nor2_1 _1828_ (.A(_0961_),
    .B(_1074_),
    .Y(_1112_));
 sky130_fd_sc_hd__and4_2 _1829_ (.A(_1012_),
    .B(_0967_),
    .C(_0969_),
    .D(_1010_),
    .X(_1113_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(net2),
    .Y(_1114_));
 sky130_fd_sc_hd__o2111ai_1 _1831_ (.A1(_1114_),
    .A2(net3),
    .B1(_1010_),
    .C1(_1053_),
    .D1(_1012_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_1 _1832_ (.A(_1055_),
    .B(_1063_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_1 _1833_ (.A(_1074_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__or4_1 _1834_ (.A(_0974_),
    .B(_0964_),
    .C(_1115_),
    .D(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__a21bo_1 _1835_ (.A1(_0943_),
    .A2(_1066_),
    .B1_N(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__a31o_1 _1836_ (.A1(_1052_),
    .A2(_1112_),
    .A3(_1113_),
    .B1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_2 _1837_ (.A(_0830_),
    .B(_0885_),
    .Y(_1121_));
 sky130_fd_sc_hd__and4bb_1 _1838_ (.A_N(_0832_),
    .B_N(_0834_),
    .C(_0835_),
    .D(_0833_),
    .X(_1122_));
 sky130_fd_sc_hd__a32o_1 _1839_ (.A1(_1122_),
    .A2(_1085_),
    .A3(_0974_),
    .B1(_1081_),
    .B2(_1088_),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_1 _1840_ (.A1(_1121_),
    .A2(_0975_),
    .B1(_0972_),
    .B2(_1054_),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a32o_1 _1841_ (.A1(_0891_),
    .A2(_1122_),
    .A3(_1091_),
    .B1(_1047_),
    .B2(_1063_),
    .X(_1125_));
 sky130_fd_sc_hd__or3_1 _1842_ (.A(_1120_),
    .B(_1124_),
    .C(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_1 _1843_ (.A(_0901_),
    .B(_0855_),
    .Y(_1127_));
 sky130_fd_sc_hd__nor2_1 _1844_ (.A(_0857_),
    .B(_1076_),
    .Y(_1128_));
 sky130_fd_sc_hd__a22o_1 _1845_ (.A1(_1128_),
    .A2(_1091_),
    .B1(_1048_),
    .B2(_1059_),
    .X(_1129_));
 sky130_fd_sc_hd__a221o_1 _1846_ (.A1(_1127_),
    .A2(_0976_),
    .B1(_1047_),
    .B2(_1055_),
    .C1(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__nor2_4 _1847_ (.A(_0830_),
    .B(_0815_),
    .Y(_1131_));
 sky130_fd_sc_hd__a22o_1 _1848_ (.A1(_1131_),
    .A2(_0974_),
    .B1(_1018_),
    .B2(_1081_),
    .X(_1132_));
 sky130_fd_sc_hd__or3_2 _1849_ (.A(_0967_),
    .B(_0969_),
    .C(_1013_),
    .X(_1133_));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(_1095_),
    .Y(_1134_));
 sky130_fd_sc_hd__o211a_1 _1851_ (.A1(_1012_),
    .A2(_0969_),
    .B1(_0956_),
    .C1(_1024_),
    .X(_1135_));
 sky130_fd_sc_hd__a31o_1 _1852_ (.A1(_0958_),
    .A2(_1086_),
    .A3(_1134_),
    .B1(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__a22o_1 _1853_ (.A1(_1033_),
    .A2(_1017_),
    .B1(_1133_),
    .B2(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__nor2_1 _1854_ (.A(_0866_),
    .B(_0815_),
    .Y(_1138_));
 sky130_fd_sc_hd__a32o_1 _1855_ (.A1(_0966_),
    .A2(_1116_),
    .A3(_1137_),
    .B1(_1066_),
    .B2(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__or2_1 _1856_ (.A(_1132_),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _1857_ (.A1(_0845_),
    .A2(_1067_),
    .B1(_1048_),
    .B2(_1055_),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _1858_ (.A1(_0927_),
    .A2(_1066_),
    .B1(_1054_),
    .B2(_1081_),
    .X(_1142_));
 sky130_fd_sc_hd__nor2_2 _1859_ (.A(_0901_),
    .B(_0844_),
    .Y(_1143_));
 sky130_fd_sc_hd__nor2_2 _1860_ (.A(_0871_),
    .B(_0844_),
    .Y(_1144_));
 sky130_fd_sc_hd__a22o_1 _1861_ (.A1(_1144_),
    .A2(_1066_),
    .B1(_1054_),
    .B2(_1087_),
    .X(_1145_));
 sky130_fd_sc_hd__a221o_1 _1862_ (.A1(_1143_),
    .A2(_1091_),
    .B1(_0972_),
    .B2(_1019_),
    .C1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__or4_1 _1863_ (.A(_1140_),
    .B(_1141_),
    .C(_1142_),
    .D(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__or3_1 _1864_ (.A(_1126_),
    .B(_1130_),
    .C(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__or3_1 _1865_ (.A(_1100_),
    .B(_1111_),
    .C(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_1 _1866_ (.A(_1149_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_4 _1867_ (.A(_0830_),
    .B(_0860_),
    .Y(_1150_));
 sky130_fd_sc_hd__and2_1 _1868_ (.A(_0999_),
    .B(_1041_),
    .X(_1151_));
 sky130_fd_sc_hd__nor2_1 _1869_ (.A(_0821_),
    .B(_0860_),
    .Y(_1152_));
 sky130_fd_sc_hd__a32o_1 _1870_ (.A1(_1052_),
    .A2(_1133_),
    .A3(_1151_),
    .B1(_1066_),
    .B2(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__a221o_1 _1871_ (.A1(_1150_),
    .A2(_0975_),
    .B1(_0972_),
    .B2(_1069_),
    .C1(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__a22o_1 _1872_ (.A1(_0839_),
    .A2(_0975_),
    .B1(_1018_),
    .B2(_1055_),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _1873_ (.A(_0866_),
    .B(_0860_),
    .Y(_1156_));
 sky130_fd_sc_hd__a22o_1 _1874_ (.A1(_1156_),
    .A2(_0974_),
    .B1(_1063_),
    .B2(_1088_),
    .X(_1157_));
 sky130_fd_sc_hd__a22o_1 _1875_ (.A1(_0908_),
    .A2(_1066_),
    .B1(_1048_),
    .B2(_1113_),
    .X(_1158_));
 sky130_fd_sc_hd__a221o_1 _1876_ (.A1(_0921_),
    .A2(_1067_),
    .B1(_1048_),
    .B2(_1081_),
    .C1(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__or4_1 _1877_ (.A(_1154_),
    .B(_1155_),
    .C(_1157_),
    .D(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__nor2_2 _1878_ (.A(_0901_),
    .B(_0818_),
    .Y(_1161_));
 sky130_fd_sc_hd__a221o_1 _1879_ (.A1(_1161_),
    .A2(_1067_),
    .B1(_1019_),
    .B2(_1095_),
    .C1(_1142_),
    .X(_1162_));
 sky130_fd_sc_hd__a32o_1 _1880_ (.A1(_1034_),
    .A2(_1052_),
    .A3(_1113_),
    .B1(_1091_),
    .B2(_0872_),
    .X(_1163_));
 sky130_fd_sc_hd__a22o_1 _1881_ (.A1(_0889_),
    .A2(_1091_),
    .B1(_1047_),
    .B2(_1113_),
    .X(_1164_));
 sky130_fd_sc_hd__or4_1 _1882_ (.A(_1140_),
    .B(_1162_),
    .C(_1163_),
    .D(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(_0866_),
    .B(_0865_),
    .Y(_1166_));
 sky130_fd_sc_hd__a22o_1 _1884_ (.A1(_1166_),
    .A2(_1067_),
    .B1(_1069_),
    .B2(_1113_),
    .X(_1167_));
 sky130_fd_sc_hd__nor2_4 _1885_ (.A(_0829_),
    .B(_0865_),
    .Y(_1168_));
 sky130_fd_sc_hd__a31o_1 _1886_ (.A1(_0964_),
    .A2(_1017_),
    .A3(_1087_),
    .B1(_0975_),
    .X(_1169_));
 sky130_fd_sc_hd__o21a_1 _1887_ (.A1(_1168_),
    .A2(_0978_),
    .B1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__a2bb2o_1 _1888_ (.A1_N(_0880_),
    .A2_N(_0978_),
    .B1(_1047_),
    .B2(_1081_),
    .X(_1171_));
 sky130_fd_sc_hd__or3_1 _1889_ (.A(_1167_),
    .B(_1170_),
    .C(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__nor2_1 _1890_ (.A(_1076_),
    .B(_0818_),
    .Y(_1173_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(_1076_),
    .B(_0865_),
    .Y(_1174_));
 sky130_fd_sc_hd__a22o_1 _1892_ (.A1(_1088_),
    .A2(_1095_),
    .B1(_1174_),
    .B2(_0975_),
    .X(_1175_));
 sky130_fd_sc_hd__a221o_1 _1893_ (.A1(_1173_),
    .A2(_1091_),
    .B1(_1060_),
    .B2(_1112_),
    .C1(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__a221o_1 _1894_ (.A1(_0847_),
    .A2(_0976_),
    .B1(_1019_),
    .B2(_1063_),
    .C1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__or4_1 _1895_ (.A(_1160_),
    .B(_1165_),
    .C(_1172_),
    .D(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__or2_1 _1896_ (.A(_1100_),
    .B(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _1897_ (.A(_1179_),
    .X(_0021_));
 sky130_fd_sc_hd__nor3_1 _1898_ (.A(_0901_),
    .B(_0825_),
    .C(_0978_),
    .Y(_1180_));
 sky130_fd_sc_hd__a21oi_1 _1899_ (.A1(_0954_),
    .A2(_1010_),
    .B1(_1040_),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_1 _1900_ (.A(_0866_),
    .B(_0825_),
    .Y(_1182_));
 sky130_fd_sc_hd__a32o_1 _1901_ (.A1(_0966_),
    .A2(_1063_),
    .A3(_1181_),
    .B1(_0974_),
    .B2(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__a2111o_1 _1902_ (.A1(_1047_),
    .A2(_1059_),
    .B1(_1092_),
    .C1(_1180_),
    .D1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__nand2_1 _1903_ (.A(_1047_),
    .B(_1087_),
    .Y(_1185_));
 sky130_fd_sc_hd__o31a_1 _1904_ (.A1(_0901_),
    .A2(_0852_),
    .A3(_0978_),
    .B1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__inv_2 _1905_ (.A(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__or4_1 _1906_ (.A(_1065_),
    .B(_1164_),
    .C(_1184_),
    .D(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__nor2_1 _1907_ (.A(_0871_),
    .B(_0825_),
    .Y(_1189_));
 sky130_fd_sc_hd__nor2_1 _1908_ (.A(_1076_),
    .B(_0825_),
    .Y(_1190_));
 sky130_fd_sc_hd__a22o_1 _1909_ (.A1(_1190_),
    .A2(_1091_),
    .B1(_1055_),
    .B2(_1088_),
    .X(_1191_));
 sky130_fd_sc_hd__a221o_1 _1910_ (.A1(_1189_),
    .A2(_0976_),
    .B1(_1069_),
    .B2(_1087_),
    .C1(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _1911_ (.A1(_0868_),
    .A2(_0976_),
    .B1(_1019_),
    .B2(_1113_),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _1912_ (.A1(_0853_),
    .A2(_0974_),
    .B1(_0972_),
    .B2(_1088_),
    .X(_1194_));
 sky130_fd_sc_hd__a32o_1 _1913_ (.A1(_0958_),
    .A2(_0966_),
    .A3(_0970_),
    .B1(_1066_),
    .B2(_0933_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _1914_ (.A(_1194_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__or2_1 _1915_ (.A(_1193_),
    .B(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__or4_1 _1916_ (.A(_1099_),
    .B(_1130_),
    .C(_1192_),
    .D(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__or4_1 _1917_ (.A(_1111_),
    .B(_1160_),
    .C(_1188_),
    .D(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _1918_ (.A(_1199_),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(_0871_),
    .B(_0882_),
    .Y(_1200_));
 sky130_fd_sc_hd__a221o_1 _1920_ (.A1(_1200_),
    .A2(_0976_),
    .B1(_1054_),
    .B2(_1095_),
    .C1(_1158_),
    .X(_1201_));
 sky130_fd_sc_hd__nor2_4 _1921_ (.A(_0827_),
    .B(_0882_),
    .Y(_1202_));
 sky130_fd_sc_hd__a221o_1 _1922_ (.A1(_1202_),
    .A2(_0976_),
    .B1(_1019_),
    .B2(_1087_),
    .C1(_1155_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _1923_ (.A(_0882_),
    .B(_1076_),
    .Y(_1204_));
 sky130_fd_sc_hd__a221o_1 _1924_ (.A1(_1060_),
    .A2(_1151_),
    .B1(_1204_),
    .B2(_1091_),
    .C1(_1089_),
    .X(_1205_));
 sky130_fd_sc_hd__or2_1 _1925_ (.A(_1203_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__or4_1 _1926_ (.A(_1172_),
    .B(_1197_),
    .C(_1201_),
    .D(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__nor3_1 _1927_ (.A(_0901_),
    .B(_0882_),
    .C(_0979_),
    .Y(_1208_));
 sky130_fd_sc_hd__a2111o_1 _1928_ (.A1(_1047_),
    .A2(_1095_),
    .B1(_1175_),
    .C1(_1208_),
    .D1(_1083_),
    .X(_1209_));
 sky130_fd_sc_hd__or4_1 _1929_ (.A(_1057_),
    .B(_1073_),
    .C(_1106_),
    .D(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a221o_1 _1930_ (.A1(_0921_),
    .A2(_0977_),
    .B1(_1048_),
    .B2(_1081_),
    .C1(_1187_),
    .X(_1211_));
 sky130_fd_sc_hd__or4_1 _1931_ (.A(_1064_),
    .B(_1126_),
    .C(_1129_),
    .D(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__or3_1 _1932_ (.A(_1207_),
    .B(_1210_),
    .C(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(_1213_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _1934_ (.A(_0816_),
    .B(_1076_),
    .Y(_1214_));
 sky130_fd_sc_hd__a22o_1 _1935_ (.A1(_1214_),
    .A2(_0976_),
    .B1(_1019_),
    .B2(_1059_),
    .X(_1215_));
 sky130_fd_sc_hd__a2111o_1 _1936_ (.A1(_1048_),
    .A2(_1087_),
    .B1(_1177_),
    .C1(_1191_),
    .D1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__or2_1 _1937_ (.A(_1078_),
    .B(_1129_),
    .X(_1217_));
 sky130_fd_sc_hd__or4_1 _1938_ (.A(_1120_),
    .B(_1141_),
    .C(_1167_),
    .D(_1196_),
    .X(_1218_));
 sky130_fd_sc_hd__or4_1 _1939_ (.A(_1056_),
    .B(_1070_),
    .C(_1098_),
    .D(_1109_),
    .X(_1219_));
 sky130_fd_sc_hd__or4_1 _1940_ (.A(_1061_),
    .B(_1123_),
    .C(_1157_),
    .D(_1183_),
    .X(_1220_));
 sky130_fd_sc_hd__a211o_1 _1941_ (.A1(_0846_),
    .A2(_1091_),
    .B1(_1104_),
    .C1(_1153_),
    .X(_1221_));
 sky130_fd_sc_hd__or4_1 _1942_ (.A(_1107_),
    .B(_1139_),
    .C(_1220_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__or3_1 _1943_ (.A(_1218_),
    .B(_1219_),
    .C(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__or4_1 _1944_ (.A(_1206_),
    .B(_1216_),
    .C(_1217_),
    .D(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _1945_ (.A(_1224_),
    .X(_0024_));
 sky130_fd_sc_hd__or3_1 _1946_ (.A(_1192_),
    .B(_1201_),
    .C(_1217_),
    .X(_1225_));
 sky130_fd_sc_hd__or4_1 _1947_ (.A(_1110_),
    .B(_1193_),
    .C(_1194_),
    .D(_1215_),
    .X(_1226_));
 sky130_fd_sc_hd__or4_1 _1948_ (.A(_1061_),
    .B(_1132_),
    .C(_1145_),
    .D(_1163_),
    .X(_1227_));
 sky130_fd_sc_hd__a2bb2o_1 _1949_ (.A1_N(_1029_),
    .A2_N(_1036_),
    .B1(_1133_),
    .B2(_1011_),
    .X(_1228_));
 sky130_fd_sc_hd__a21o_1 _1950_ (.A1(_1055_),
    .A2(_1181_),
    .B1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__a221o_1 _1951_ (.A1(_0831_),
    .A2(_0977_),
    .B1(_0966_),
    .B2(_1229_),
    .C1(_1170_),
    .X(_1230_));
 sky130_fd_sc_hd__or3_1 _1952_ (.A(_1050_),
    .B(_1227_),
    .C(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__or4_1 _1953_ (.A(_1072_),
    .B(_1096_),
    .C(_1101_),
    .D(_1124_),
    .X(_1232_));
 sky130_fd_sc_hd__or4_1 _1954_ (.A(_1154_),
    .B(_1176_),
    .C(_1205_),
    .D(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__or4_1 _1955_ (.A(_1225_),
    .B(_1226_),
    .C(_1231_),
    .D(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _1956_ (.A(_1234_),
    .X(_0025_));
 sky130_fd_sc_hd__and2b_1 _1957_ (.A_N(\pulse_slower.currentEnableState[1] ),
    .B(net98),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _1958_ (.A(_1235_),
    .X(\pulse_slower.nextEnableState[1] ));
 sky130_fd_sc_hd__inv_2 _1959_ (.A(net11),
    .Y(\instructionLoader.interruptInjector.nmiSync.in ));
 sky130_fd_sc_hd__inv_2 _1960_ (.A(net10),
    .Y(\instructionLoader.interruptInjector.interruptRequest ));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(net1),
    .B(_0950_),
    .Y(net40));
 sky130_fd_sc_hd__and2_2 _1962_ (.A(clknet_4_4_0_clk),
    .B(\pulse_slower.nextEnableState[0] ),
    .X(_1236_));
 sky130_fd_sc_hd__buf_1 _1963_ (.A(_1236_),
    .X(net41));
 sky130_fd_sc_hd__a41oi_4 _1964_ (.A1(_0909_),
    .A2(_0885_),
    .A3(_0865_),
    .A4(_0852_),
    .B1(_0821_),
    .Y(_1237_));
 sky130_fd_sc_hd__a311oi_2 _1965_ (.A1(_0844_),
    .A2(_0882_),
    .A3(_0852_),
    .B1(_0871_),
    .C1(_0917_),
    .Y(_1238_));
 sky130_fd_sc_hd__a311oi_2 _1966_ (.A1(_0844_),
    .A2(_0815_),
    .A3(_0818_),
    .B1(_0901_),
    .C1(_0917_),
    .Y(_1239_));
 sky130_fd_sc_hd__and2_1 _1967_ (.A(\demux.isAddressing ),
    .B(_0947_),
    .X(_1240_));
 sky130_fd_sc_hd__buf_4 _1968_ (.A(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__a2111o_1 _1969_ (.A1(_0875_),
    .A2(_1237_),
    .B1(_1238_),
    .C1(_1239_),
    .D1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__or2_1 _1970_ (.A(\demux.state_machine.timeState[0] ),
    .B(\demux.state_machine.timeState[4] ),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_4 _1971_ (.A(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_1 _1972_ (.A(_1003_),
    .B(_0913_),
    .Y(_1245_));
 sky130_fd_sc_hd__o21ai_1 _1973_ (.A1(_0847_),
    .A2(_0873_),
    .B1(_0877_),
    .Y(_1246_));
 sky130_fd_sc_hd__or4bb_1 _1974_ (.A(_1166_),
    .B(_0910_),
    .C_N(_1245_),
    .D_N(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__a21oi_2 _1975_ (.A1(_0855_),
    .A2(_0860_),
    .B1(_0827_),
    .Y(_1248_));
 sky130_fd_sc_hd__or2_2 _1976_ (.A(_0828_),
    .B(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__or4_1 _1977_ (.A(_1121_),
    .B(_0943_),
    .C(_1131_),
    .D(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_1 _1978_ (.A1(_0877_),
    .A2(_0915_),
    .B1(_0930_),
    .B2(_1004_),
    .X(_1251_));
 sky130_fd_sc_hd__a221o_1 _1979_ (.A1(_1244_),
    .A2(_1247_),
    .B1(_1250_),
    .B2(_1001_),
    .C1(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__a21oi_1 _1980_ (.A1(_0988_),
    .A2(_0993_),
    .B1(_0948_),
    .Y(_1253_));
 sky130_fd_sc_hd__o21ai_1 _1981_ (.A1(_1077_),
    .A2(_1173_),
    .B1(_0995_),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _1982_ (.A(_1253_),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__o211a_1 _1983_ (.A1(_1242_),
    .A2(_1252_),
    .B1(_1255_),
    .C1(_0998_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_8 _1984_ (.A(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__a22o_1 _1985_ (.A1(_0897_),
    .A2(_0912_),
    .B1(_0920_),
    .B2(_0876_),
    .X(_1258_));
 sky130_fd_sc_hd__and3b_2 _1986_ (.A_N(_0832_),
    .B(_0939_),
    .C(_0940_),
    .X(_1259_));
 sky130_fd_sc_hd__and2_1 _1987_ (.A(_0932_),
    .B(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__a22o_1 _1988_ (.A1(_0897_),
    .A2(_1079_),
    .B1(_1260_),
    .B2(_0833_),
    .X(_1261_));
 sky130_fd_sc_hd__o21ai_4 _1989_ (.A1(_1258_),
    .A2(_1261_),
    .B1(_0948_),
    .Y(_1262_));
 sky130_fd_sc_hd__clkbuf_4 _1990_ (.A(_0932_),
    .X(_1263_));
 sky130_fd_sc_hd__o21a_1 _1991_ (.A1(_0927_),
    .A2(_1143_),
    .B1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__inv_2 _1992_ (.A(\demux.state_machine.timeState[6] ),
    .Y(_1265_));
 sky130_fd_sc_hd__nor3_1 _1993_ (.A(_1265_),
    .B(_0871_),
    .C(_0865_),
    .Y(_1266_));
 sky130_fd_sc_hd__and3_2 _1994_ (.A(\demux.state_machine.timeState[1] ),
    .B(_0891_),
    .C(_1084_),
    .X(_1267_));
 sky130_fd_sc_hd__inv_2 _1995_ (.A(\demux.state_machine.timeState[0] ),
    .Y(_1268_));
 sky130_fd_sc_hd__or4_1 _1996_ (.A(_1268_),
    .B(_0832_),
    .C(_0827_),
    .D(_0858_),
    .X(_1269_));
 sky130_fd_sc_hd__or3b_1 _1997_ (.A(_1266_),
    .B(_1267_),
    .C_N(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__a21oi_4 _1998_ (.A1(_0818_),
    .A2(_0861_),
    .B1(_0901_),
    .Y(_1271_));
 sky130_fd_sc_hd__o31a_1 _1999_ (.A1(_0868_),
    .A2(_1131_),
    .A3(_1271_),
    .B1(_1263_),
    .X(_1272_));
 sky130_fd_sc_hd__buf_4 _2000_ (.A(_1268_),
    .X(_1273_));
 sky130_fd_sc_hd__a311oi_4 _2001_ (.A1(_0815_),
    .A2(_0818_),
    .A3(_0825_),
    .B1(_0866_),
    .C1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__and4b_1 _2002_ (.A_N(_0835_),
    .B(_0834_),
    .C(_0833_),
    .D(_0832_),
    .X(_1275_));
 sky130_fd_sc_hd__and3_1 _2003_ (.A(_0896_),
    .B(_0939_),
    .C(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a211o_1 _2004_ (.A1(_0897_),
    .A2(_0913_),
    .B1(_1274_),
    .C1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__nor4_1 _2005_ (.A(_1264_),
    .B(_1270_),
    .C(_1272_),
    .D(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__and2_1 _2006_ (.A(_0932_),
    .B(_0926_),
    .X(_1279_));
 sky130_fd_sc_hd__a221oi_4 _2007_ (.A1(_1003_),
    .A2(_0840_),
    .B1(_1150_),
    .B2(_0897_),
    .C1(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__a21oi_2 _2008_ (.A1(_1003_),
    .A2(_0904_),
    .B1(_1241_),
    .Y(_1281_));
 sky130_fd_sc_hd__or2_1 _2009_ (.A(\demux.state_machine.timeState[0] ),
    .B(_0896_),
    .X(_1282_));
 sky130_fd_sc_hd__and2b_1 _2010_ (.A_N(_0993_),
    .B(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__o21a_1 _2011_ (.A1(_0988_),
    .A2(\demux.state_machine.currentAddress[6] ),
    .B1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__or3_4 _2012_ (.A(\demux.state_machine.timeState[0] ),
    .B(_0896_),
    .C(\demux.state_machine.timeState[4] ),
    .X(_1285_));
 sky130_fd_sc_hd__a22o_1 _2013_ (.A1(_0932_),
    .A2(_0991_),
    .B1(_1285_),
    .B2(\demux.state_machine.currentAddress[1] ),
    .X(_1286_));
 sky130_fd_sc_hd__a211o_1 _2014_ (.A1(_0985_),
    .A2(_1244_),
    .B1(_1286_),
    .C1(_0948_),
    .X(_1287_));
 sky130_fd_sc_hd__nor2_1 _2015_ (.A(_1284_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__a31o_2 _2016_ (.A1(_1278_),
    .A2(_1280_),
    .A3(_1281_),
    .B1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a21oi_4 _2017_ (.A1(_0888_),
    .A2(net52),
    .B1(_0917_),
    .Y(_1290_));
 sky130_fd_sc_hd__o21a_1 _2018_ (.A1(_0912_),
    .A2(_1079_),
    .B1(_1003_),
    .X(_1291_));
 sky130_fd_sc_hd__a211o_1 _2019_ (.A1(\branch_ff.branchForward ),
    .A2(_1290_),
    .B1(_1291_),
    .C1(_1261_),
    .X(_1292_));
 sky130_fd_sc_hd__and4_1 _2020_ (.A(_0952_),
    .B(_1262_),
    .C(_1289_),
    .D(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__buf_2 _2021_ (.A(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__a32o_1 _2022_ (.A1(_0897_),
    .A2(_0985_),
    .A3(_0986_),
    .B1(net54),
    .B2(\demux.state_machine.currentAddress[1] ),
    .X(_1295_));
 sky130_fd_sc_hd__a211o_1 _2023_ (.A1(_0988_),
    .A2(net54),
    .B1(_1295_),
    .C1(_0995_),
    .X(_1296_));
 sky130_fd_sc_hd__a21o_1 _2024_ (.A1(_1214_),
    .A2(_1296_),
    .B1(_0948_),
    .X(_1297_));
 sky130_fd_sc_hd__a21oi_2 _2025_ (.A1(_0885_),
    .A2(_0865_),
    .B1(_1076_),
    .Y(_1298_));
 sky130_fd_sc_hd__o21a_1 _2026_ (.A1(_1189_),
    .A2(_1298_),
    .B1(_1263_),
    .X(_1299_));
 sky130_fd_sc_hd__or3_1 _2027_ (.A(_1241_),
    .B(_1299_),
    .C(_1258_),
    .X(_1300_));
 sky130_fd_sc_hd__o2111a_1 _2028_ (.A1(net13),
    .A2(_0950_),
    .B1(_1297_),
    .C1(_1300_),
    .D1(\pulse_slower.nextEnableState[0] ),
    .X(_1301_));
 sky130_fd_sc_hd__a211oi_4 _2029_ (.A1(_1262_),
    .A2(_1289_),
    .B1(_0960_),
    .C1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__clkbuf_4 _2030_ (.A(_0952_),
    .X(_1303_));
 sky130_fd_sc_hd__a21boi_1 _2031_ (.A1(_1303_),
    .A2(_1292_),
    .B1_N(_1301_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(\branch_ff.branchBackward ),
    .B(_1290_),
    .Y(_1305_));
 sky130_fd_sc_hd__o21a_1 _2033_ (.A1(_0876_),
    .A2(_0879_),
    .B1(_0912_),
    .X(_1306_));
 sky130_fd_sc_hd__or2_1 _2034_ (.A(_0941_),
    .B(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__inv_2 _2035_ (.A(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__o21ai_1 _2036_ (.A1(_1097_),
    .A2(_1248_),
    .B1(_1004_),
    .Y(_1309_));
 sky130_fd_sc_hd__a211o_1 _2037_ (.A1(_0959_),
    .A2(net42),
    .B1(_0951_),
    .C1(_1241_),
    .X(_1310_));
 sky130_fd_sc_hd__a31o_1 _2038_ (.A1(_1305_),
    .A2(_1308_),
    .A3(_1309_),
    .B1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__nor4_1 _2039_ (.A(_1302_),
    .B(_1294_),
    .C(_1304_),
    .D(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _2040_ (.A(_1303_),
    .B(_1292_),
    .Y(_1313_));
 sky130_fd_sc_hd__and2_2 _2041_ (.A(_1313_),
    .B(_1302_),
    .X(_1314_));
 sky130_fd_sc_hd__a21boi_4 _2042_ (.A1(_1262_),
    .A2(_1289_),
    .B1_N(_1304_),
    .Y(_1315_));
 sky130_fd_sc_hd__and3_2 _2043_ (.A(_1301_),
    .B(_1262_),
    .C(_1289_),
    .X(_1316_));
 sky130_fd_sc_hd__and2_1 _2044_ (.A(_0952_),
    .B(_1292_),
    .X(_1317_));
 sky130_fd_sc_hd__and2_2 _2045_ (.A(_1317_),
    .B(_1302_),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _2046_ (.A1(\internalDataflow.accRegToDB[6] ),
    .A2(_1316_),
    .B1(_1318_),
    .B2(\demux.PSR_V ),
    .X(_1319_));
 sky130_fd_sc_hd__a221o_1 _2047_ (.A1(net8),
    .A2(_1314_),
    .B1(_1315_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[22] ),
    .C1(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__a211o_1 _2048_ (.A1(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .A2(_1294_),
    .B1(net134),
    .C1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__nor2_1 _2049_ (.A(_1257_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__nand2_1 _2050_ (.A(_1005_),
    .B(_0927_),
    .Y(_1323_));
 sky130_fd_sc_hd__nand2_2 _2051_ (.A(_1005_),
    .B(_0905_),
    .Y(_1324_));
 sky130_fd_sc_hd__buf_4 _2052_ (.A(_1310_),
    .X(_1325_));
 sky130_fd_sc_hd__a31oi_4 _2053_ (.A1(_1323_),
    .A2(_1280_),
    .A3(_1324_),
    .B1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a31o_1 _2054_ (.A1(_1323_),
    .A2(_1280_),
    .A3(_1324_),
    .B1(_1325_),
    .X(_1327_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(_1256_),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__clkbuf_4 _2056_ (.A(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__and3_2 _2057_ (.A(_0891_),
    .B(_1084_),
    .C(_1285_),
    .X(_1330_));
 sky130_fd_sc_hd__nor4_1 _2058_ (.A(\demux.state_machine.currentAddress[11] ),
    .B(_0988_),
    .C(\demux.state_machine.currentAddress[4] ),
    .D(_0948_),
    .Y(_1331_));
 sky130_fd_sc_hd__o2bb2a_1 _2059_ (.A1_N(_1173_),
    .A2_N(_0995_),
    .B1(_1331_),
    .B2(_1273_),
    .X(_1332_));
 sky130_fd_sc_hd__or4_1 _2060_ (.A(_1138_),
    .B(_1058_),
    .C(_0867_),
    .D(_1204_),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_1 _2061_ (.A1(_1003_),
    .A2(_1333_),
    .B1(_1241_),
    .Y(_1334_));
 sky130_fd_sc_hd__a2111oi_1 _2062_ (.A1(_0959_),
    .A2(net42),
    .B1(_1332_),
    .C1(_1334_),
    .D1(_0951_),
    .Y(_1335_));
 sky130_fd_sc_hd__a21o_1 _2063_ (.A1(_1263_),
    .A2(_1150_),
    .B1(_0941_),
    .X(_1336_));
 sky130_fd_sc_hd__o31a_1 _2064_ (.A1(_1152_),
    .A2(_0913_),
    .A3(_1094_),
    .B1(_1263_),
    .X(_1337_));
 sky130_fd_sc_hd__o41a_1 _2065_ (.A1(_0868_),
    .A2(_1143_),
    .A3(_1131_),
    .A4(_1271_),
    .B1(_1263_),
    .X(_1338_));
 sky130_fd_sc_hd__o41a_1 _2066_ (.A1(_0847_),
    .A2(_0856_),
    .A3(_1202_),
    .A4(_1237_),
    .B1(_1263_),
    .X(_1339_));
 sky130_fd_sc_hd__nor4_1 _2067_ (.A(_1336_),
    .B(_1337_),
    .C(_1338_),
    .D(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a2111o_1 _2068_ (.A1(_0959_),
    .A2(net42),
    .B1(net51),
    .C1(_1241_),
    .D1(_0951_),
    .X(_1341_));
 sky130_fd_sc_hd__or2b_1 _2069_ (.A(net135),
    .B_N(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__or4_1 _2070_ (.A(_1182_),
    .B(_1128_),
    .C(_0910_),
    .D(_1097_),
    .X(_1343_));
 sky130_fd_sc_hd__o21ai_1 _2071_ (.A1(_0987_),
    .A2(_1077_),
    .B1(_0876_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2_1 _2072_ (.A(_1273_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__a22o_2 _2073_ (.A1(_1003_),
    .A2(_1343_),
    .B1(_1345_),
    .B2(_1241_),
    .X(_1346_));
 sky130_fd_sc_hd__or4_1 _2074_ (.A(_1263_),
    .B(\demux.state_machine.currentAddress[11] ),
    .C(\demux.state_machine.currentAddress[1] ),
    .D(\demux.state_machine.currentAddress[7] ),
    .X(_1347_));
 sky130_fd_sc_hd__a211o_1 _2075_ (.A1(\demux.state_machine.currentAddress[5] ),
    .A2(_1077_),
    .B1(\demux.state_machine.currentAddress[10] ),
    .C1(_1273_),
    .X(_1348_));
 sky130_fd_sc_hd__a211o_2 _2076_ (.A1(_1347_),
    .A2(_1348_),
    .B1(\demux.state_machine.currentAddress[3] ),
    .C1(_0948_),
    .X(_1349_));
 sky130_fd_sc_hd__a31oi_4 _2077_ (.A1(_0998_),
    .A2(_1346_),
    .A3(_1349_),
    .B1(net49),
    .Y(_1350_));
 sky130_fd_sc_hd__o21a_1 _2078_ (.A1(_1336_),
    .A2(_1337_),
    .B1(_0982_),
    .X(_1351_));
 sky130_fd_sc_hd__or2_1 _2079_ (.A(\branch_ff.branchForward ),
    .B(\branch_ff.branchBackward ),
    .X(_1352_));
 sky130_fd_sc_hd__a22o_1 _2080_ (.A1(_1051_),
    .A2(_1084_),
    .B1(_1122_),
    .B2(_0939_),
    .X(_1353_));
 sky130_fd_sc_hd__o311a_1 _2081_ (.A1(\demux.state_machine.timeState[4] ),
    .A2(\demux.state_machine.timeState[6] ),
    .A3(\demux.state_machine.timeState[1] ),
    .B1(_1051_),
    .C1(_0890_),
    .X(_1354_));
 sky130_fd_sc_hd__a2111o_1 _2082_ (.A1(_0876_),
    .A2(_1353_),
    .B1(_1354_),
    .C1(_0918_),
    .D1(_0916_),
    .X(_1355_));
 sky130_fd_sc_hd__a31o_1 _2083_ (.A1(_0897_),
    .A2(_0904_),
    .A3(_1352_),
    .B1(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__or2_1 _2084_ (.A(_0847_),
    .B(_0873_),
    .X(_1357_));
 sky130_fd_sc_hd__or2_2 _2085_ (.A(_0943_),
    .B(_1166_),
    .X(_1358_));
 sky130_fd_sc_hd__o41a_1 _2086_ (.A1(_0915_),
    .A2(_1357_),
    .A3(_1249_),
    .A4(_1358_),
    .B1(_0876_),
    .X(_1359_));
 sky130_fd_sc_hd__and3_1 _2087_ (.A(_0896_),
    .B(_0939_),
    .C(_1084_),
    .X(_1360_));
 sky130_fd_sc_hd__and3_1 _2088_ (.A(\demux.state_machine.timeState[6] ),
    .B(_0891_),
    .C(_1084_),
    .X(_1361_));
 sky130_fd_sc_hd__a2111o_1 _2089_ (.A1(_0875_),
    .A2(_0930_),
    .B1(_1266_),
    .C1(_1360_),
    .D1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__or3_1 _2090_ (.A(_0924_),
    .B(_1242_),
    .C(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__inv_2 _2091_ (.A(_1253_),
    .Y(_1364_));
 sky130_fd_sc_hd__o32a_1 _2092_ (.A1(_1356_),
    .A2(_1359_),
    .A3(_1363_),
    .B1(_1295_),
    .B2(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__o21a_2 _2093_ (.A1(_1351_),
    .A2(_1365_),
    .B1(_0998_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(_1342_),
    .A1(_1350_),
    .S(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__and2b_1 _2095_ (.A_N(net135),
    .B(_1341_),
    .X(_1368_));
 sky130_fd_sc_hd__a31o_1 _2096_ (.A1(_0997_),
    .A2(_1346_),
    .A3(_1349_),
    .B1(_1335_),
    .X(_1369_));
 sky130_fd_sc_hd__and3b_1 _2097_ (.A_N(_1366_),
    .B(_1368_),
    .C(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_4 _2098_ (.A(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__a211o_4 _2099_ (.A1(_1303_),
    .A2(_1330_),
    .B1(_1367_),
    .C1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__and3b_2 _2100_ (.A_N(_1366_),
    .B(_1342_),
    .C(_1369_),
    .X(_1373_));
 sky130_fd_sc_hd__and3b_2 _2101_ (.A_N(_1366_),
    .B(_1342_),
    .C(_1350_),
    .X(_1374_));
 sky130_fd_sc_hd__nor2_2 _2102_ (.A(_1370_),
    .B(_1367_),
    .Y(_1375_));
 sky130_fd_sc_hd__a221o_1 _2103_ (.A1(\internalDataflow.stackBusModule.busInputs[46] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[6] ),
    .C1(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__and3_2 _2104_ (.A(_1366_),
    .B(_1341_),
    .C(_1350_),
    .X(_1377_));
 sky130_fd_sc_hd__and4b_2 _2105_ (.A_N(net50),
    .B(_1350_),
    .C(_1303_),
    .D(_1366_),
    .X(_1378_));
 sky130_fd_sc_hd__a22o_1 _2106_ (.A1(\internalDataflow.addressLowBusModule.busInputs[30] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[38] ),
    .X(_1379_));
 sky130_fd_sc_hd__a211o_1 _2107_ (.A1(\internalDataflow.stackBusModule.busInputs[38] ),
    .A2(_1371_),
    .B1(_1376_),
    .C1(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__o21a_1 _2108_ (.A1(_1102_),
    .A2(_0944_),
    .B1(_1004_),
    .X(_1381_));
 sky130_fd_sc_hd__a21oi_2 _2109_ (.A1(\branch_ff.branchBackward ),
    .A2(_1290_),
    .B1(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__or2_2 _2110_ (.A(_1325_),
    .B(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_4 _2111_ (.A(_1241_),
    .X(_1384_));
 sky130_fd_sc_hd__a31o_1 _2112_ (.A1(_0983_),
    .A2(_0905_),
    .A3(_1352_),
    .B1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__o211a_2 _2113_ (.A1(_0982_),
    .A2(_1295_),
    .B1(_1385_),
    .C1(_0998_),
    .X(_1386_));
 sky130_fd_sc_hd__nor3_2 _2114_ (.A(_1326_),
    .B(_1383_),
    .C(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a21oi_2 _2115_ (.A1(_1382_),
    .A2(_1328_),
    .B1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__o21a_1 _2116_ (.A1(_0912_),
    .A2(_1168_),
    .B1(\demux.state_machine.timeState[5] ),
    .X(_1389_));
 sky130_fd_sc_hd__a21o_1 _2117_ (.A1(_0882_),
    .A2(_0861_),
    .B1(_0830_),
    .X(_1390_));
 sky130_fd_sc_hd__nor2_1 _2118_ (.A(_0937_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a2111o_1 _2119_ (.A1(_0875_),
    .A2(_0911_),
    .B1(_1389_),
    .C1(_1391_),
    .D1(_0934_),
    .X(_1392_));
 sky130_fd_sc_hd__o21a_1 _2120_ (.A1(_0831_),
    .A2(_0837_),
    .B1(_1244_),
    .X(_1393_));
 sky130_fd_sc_hd__a221o_1 _2121_ (.A1(_0936_),
    .A2(_1144_),
    .B1(_0872_),
    .B2(_0875_),
    .C1(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__a22o_1 _2122_ (.A1(_0936_),
    .A2(_0927_),
    .B1(_0847_),
    .B2(\demux.state_machine.timeState[0] ),
    .X(_1395_));
 sky130_fd_sc_hd__o21a_1 _2123_ (.A1(_0870_),
    .A2(_1131_),
    .B1(_1243_),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _2124_ (.A1(_1259_),
    .A2(_0945_),
    .B1(_1150_),
    .B2(_0936_),
    .X(_1397_));
 sky130_fd_sc_hd__a2111o_1 _2125_ (.A1(_0875_),
    .A2(_0848_),
    .B1(_1395_),
    .C1(_1396_),
    .D1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__a22o_1 _2126_ (.A1(_0936_),
    .A2(_1121_),
    .B1(_0868_),
    .B2(_1243_),
    .X(_1399_));
 sky130_fd_sc_hd__or2_1 _2127_ (.A(\demux.state_machine.timeState[1] ),
    .B(\demux.state_machine.timeState[5] ),
    .X(_1400_));
 sky130_fd_sc_hd__a221o_1 _2128_ (.A1(_0839_),
    .A2(_1243_),
    .B1(_1400_),
    .B2(_1071_),
    .C1(_1240_),
    .X(_1401_));
 sky130_fd_sc_hd__a2111o_1 _2129_ (.A1(_0879_),
    .A2(_0912_),
    .B1(_0922_),
    .C1(_1399_),
    .D1(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__or4_1 _2130_ (.A(_1392_),
    .B(_1394_),
    .C(_1398_),
    .D(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__o31a_1 _2131_ (.A1(_0863_),
    .A2(_0867_),
    .A3(_1097_),
    .B1(_0876_),
    .X(_1404_));
 sky130_fd_sc_hd__o41ai_2 _2132_ (.A1(_0823_),
    .A2(_0828_),
    .A3(_1202_),
    .A4(_1404_),
    .B1(_1244_),
    .Y(_1405_));
 sky130_fd_sc_hd__or2_1 _2133_ (.A(_0937_),
    .B(_0928_),
    .X(_1406_));
 sky130_fd_sc_hd__and3b_1 _2134_ (.A_N(_1403_),
    .B(_1405_),
    .C(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(_0873_),
    .B(_1244_),
    .Y(_1408_));
 sky130_fd_sc_hd__or3_1 _2136_ (.A(_1004_),
    .B(_0877_),
    .C(_0879_),
    .X(_1409_));
 sky130_fd_sc_hd__o21ai_2 _2137_ (.A1(_0899_),
    .A2(_1409_),
    .B1(_0905_),
    .Y(_1410_));
 sky130_fd_sc_hd__o21a_1 _2138_ (.A1(_0912_),
    .A2(_1168_),
    .B1(\demux.state_machine.timeState[1] ),
    .X(_1411_));
 sky130_fd_sc_hd__a221o_1 _2139_ (.A1(\demux.state_machine.timeState[5] ),
    .A2(_1079_),
    .B1(_1071_),
    .B2(_0879_),
    .C1(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__and2b_1 _2140_ (.A_N(_0896_),
    .B(\demux.state_machine.timeState[6] ),
    .X(_1413_));
 sky130_fd_sc_hd__o21ai_1 _2141_ (.A1(_0875_),
    .A2(_1413_),
    .B1(\demux.state_machine.currentAddress[6] ),
    .Y(_1414_));
 sky130_fd_sc_hd__o21a_1 _2142_ (.A1(_1263_),
    .A2(_1414_),
    .B1(_1241_),
    .X(_1415_));
 sky130_fd_sc_hd__inv_2 _2143_ (.A(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__a221o_1 _2144_ (.A1(\demux.state_machine.currentAddress[7] ),
    .A2(_0993_),
    .B1(_0989_),
    .B2(_0988_),
    .C1(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__o311a_2 _2145_ (.A1(_1384_),
    .A2(_1381_),
    .A3(_1412_),
    .B1(_1417_),
    .C1(_0998_),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_1 _2146_ (.A(\demux.state_machine.currentAddress[6] ),
    .B(_1283_),
    .Y(_1419_));
 sky130_fd_sc_hd__o21ai_2 _2147_ (.A1(\demux.state_machine.currentAddress[7] ),
    .A2(_0985_),
    .B1(_1004_),
    .Y(_1420_));
 sky130_fd_sc_hd__a31o_1 _2148_ (.A1(_1384_),
    .A2(_1419_),
    .A3(_1420_),
    .B1(_0960_),
    .X(_1421_));
 sky130_fd_sc_hd__a311o_4 _2149_ (.A1(_1407_),
    .A2(_1408_),
    .A3(_1410_),
    .B1(_1418_),
    .C1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__a31o_1 _2150_ (.A1(_1407_),
    .A2(_1408_),
    .A3(_1410_),
    .B1(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__nand2_2 _2151_ (.A(_1423_),
    .B(_1418_),
    .Y(_1424_));
 sky130_fd_sc_hd__o21a_1 _2152_ (.A1(_1267_),
    .A2(_1361_),
    .B1(_1303_),
    .X(_1425_));
 sky130_fd_sc_hd__o21ai_1 _2153_ (.A1(_1102_),
    .A2(_0930_),
    .B1(_1001_),
    .Y(_1426_));
 sky130_fd_sc_hd__o21ai_2 _2154_ (.A1(_1259_),
    .A2(_1079_),
    .B1(_1003_),
    .Y(_1427_));
 sky130_fd_sc_hd__and3_1 _2155_ (.A(_1245_),
    .B(_1426_),
    .C(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__and2_1 _2156_ (.A(_1425_),
    .B(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__xnor2_1 _2157_ (.A(_1423_),
    .B(_1418_),
    .Y(_1430_));
 sky130_fd_sc_hd__or2_2 _2158_ (.A(_1429_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__o221a_1 _2159_ (.A1(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(net8),
    .C1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a32o_1 _2160_ (.A1(_1372_),
    .A2(_1380_),
    .A3(_1388_),
    .B1(_1432_),
    .B2(net47),
    .X(_1433_));
 sky130_fd_sc_hd__o2bb2a_2 _2161_ (.A1_N(_1322_),
    .A2_N(_1326_),
    .B1(_1329_),
    .B2(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _2162_ (.A(\demux.state_machine.currentAddress[11] ),
    .B(\demux.state_machine.currentAddress[3] ),
    .X(_1435_));
 sky130_fd_sc_hd__or4_1 _2163_ (.A(_0988_),
    .B(\demux.state_machine.currentAddress[4] ),
    .C(\demux.state_machine.currentAddress[10] ),
    .D(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__a21oi_1 _2164_ (.A1(_0987_),
    .A2(_0993_),
    .B1(_0982_),
    .Y(_1437_));
 sky130_fd_sc_hd__a21bo_1 _2165_ (.A1(_1006_),
    .A2(_1436_),
    .B1_N(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _2166_ (.A(\branch_ff.branchForward ),
    .B(_1290_),
    .Y(_1439_));
 sky130_fd_sc_hd__o21ai_1 _2167_ (.A1(_0930_),
    .A2(_1358_),
    .B1(_1005_),
    .Y(_1440_));
 sky130_fd_sc_hd__or3_2 _2168_ (.A(_1003_),
    .B(_0879_),
    .C(_0945_),
    .X(_1441_));
 sky130_fd_sc_hd__a22o_1 _2169_ (.A1(_1071_),
    .A2(_1285_),
    .B1(_1441_),
    .B2(_1168_),
    .X(_1442_));
 sky130_fd_sc_hd__a211o_1 _2170_ (.A1(_1005_),
    .A2(_1102_),
    .B1(_1267_),
    .C1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a21o_1 _2171_ (.A1(_1005_),
    .A2(_0910_),
    .B1(_1384_),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _2172_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__a22o_1 _2173_ (.A1(_1005_),
    .A2(\demux.state_machine.currentAddress[7] ),
    .B1(_0993_),
    .B2(_0985_),
    .X(_1446_));
 sky130_fd_sc_hd__a31o_1 _2174_ (.A1(_1273_),
    .A2(_0988_),
    .A3(_0945_),
    .B1(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__o21a_1 _2175_ (.A1(_0987_),
    .A2(\demux.state_machine.currentAddress[6] ),
    .B1(_1283_),
    .X(_1448_));
 sky130_fd_sc_hd__nor3_1 _2176_ (.A(_0982_),
    .B(_1447_),
    .C(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__a31o_1 _2177_ (.A1(_1439_),
    .A2(_1440_),
    .A3(_1445_),
    .B1(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_1 _2178_ (.A(_0982_),
    .B(_1324_),
    .Y(_1451_));
 sky130_fd_sc_hd__and2_1 _2179_ (.A(_1004_),
    .B(_1237_),
    .X(_1452_));
 sky130_fd_sc_hd__and2_1 _2180_ (.A(_1004_),
    .B(_0868_),
    .X(_1453_));
 sky130_fd_sc_hd__or4_1 _2181_ (.A(_1264_),
    .B(_1279_),
    .C(_1452_),
    .D(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__or3_1 _2182_ (.A(_1161_),
    .B(_1131_),
    .C(_0915_),
    .X(_1455_));
 sky130_fd_sc_hd__o31a_1 _2183_ (.A1(_1357_),
    .A2(_1249_),
    .A3(_1455_),
    .B1(_1004_),
    .X(_1456_));
 sky130_fd_sc_hd__or3_1 _2184_ (.A(_1307_),
    .B(_1330_),
    .C(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__or4b_1 _2185_ (.A(_1451_),
    .B(_1454_),
    .C(_1457_),
    .D_N(_1305_),
    .X(_1458_));
 sky130_fd_sc_hd__and4_1 _2186_ (.A(_0998_),
    .B(_1438_),
    .C(_1450_),
    .D(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__buf_2 _2187_ (.A(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _2188_ (.A(_1434_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__and2_1 _2189_ (.A(_1006_),
    .B(_0905_),
    .X(_1462_));
 sky130_fd_sc_hd__a221o_1 _2190_ (.A1(_1006_),
    .A2(_1102_),
    .B1(_1168_),
    .B2(_0983_),
    .C1(_1330_),
    .X(_1463_));
 sky130_fd_sc_hd__a211o_1 _2191_ (.A1(_1001_),
    .A2(_0913_),
    .B1(_1462_),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_2 _2192_ (.A(_1303_),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _2193_ (.A(_1274_),
    .B(_1453_),
    .Y(_1466_));
 sky130_fd_sc_hd__nor2_2 _2194_ (.A(_1325_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__inv_2 _2195_ (.A(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__and2_1 _2196_ (.A(_0888_),
    .B(net53),
    .X(_1469_));
 sky130_fd_sc_hd__and3b_1 _2197_ (.A_N(_1469_),
    .B(_1352_),
    .C(_1001_),
    .X(_1470_));
 sky130_fd_sc_hd__or4b_1 _2198_ (.A(_0913_),
    .B(_1298_),
    .C(_1248_),
    .D_N(_1390_),
    .X(_1471_));
 sky130_fd_sc_hd__o32a_1 _2199_ (.A1(_0873_),
    .A2(_0910_),
    .A3(_1471_),
    .B1(_1360_),
    .B2(_1006_),
    .X(_1472_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(_1006_),
    .B(_1455_),
    .X(_1473_));
 sky130_fd_sc_hd__or2_1 _2201_ (.A(_1264_),
    .B(_1336_),
    .X(_1474_));
 sky130_fd_sc_hd__a211o_1 _2202_ (.A1(_1006_),
    .A2(_1358_),
    .B1(_1473_),
    .C1(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__or4_1 _2203_ (.A(_1384_),
    .B(_1266_),
    .C(_1267_),
    .D(_1306_),
    .X(_1476_));
 sky130_fd_sc_hd__a221o_1 _2204_ (.A1(\demux.state_machine.currentAddress[6] ),
    .A2(_1283_),
    .B1(_1285_),
    .B2(_0988_),
    .C1(_1287_),
    .X(_1477_));
 sky130_fd_sc_hd__and2_2 _2205_ (.A(_0998_),
    .B(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__o41a_2 _2206_ (.A1(_1470_),
    .A2(_1472_),
    .A3(_1475_),
    .A4(_1476_),
    .B1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__inv_2 _2207_ (.A(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _2208_ (.A(_1372_),
    .B(_1380_),
    .Y(_1481_));
 sky130_fd_sc_hd__a21oi_4 _2209_ (.A1(_1257_),
    .A2(_1481_),
    .B1(_1322_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux2_1 _2210_ (.A0(_1468_),
    .A1(_1480_),
    .S(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__a31oi_2 _2211_ (.A1(_1384_),
    .A2(_1419_),
    .A3(_1420_),
    .B1(_0960_),
    .Y(_1484_));
 sky130_fd_sc_hd__a311o_1 _2212_ (.A1(_0876_),
    .A2(_0888_),
    .A3(net53),
    .B1(_0936_),
    .C1(_1263_),
    .X(_1485_));
 sky130_fd_sc_hd__and3_1 _2213_ (.A(_0891_),
    .B(_1275_),
    .C(_1244_),
    .X(_1486_));
 sky130_fd_sc_hd__a21o_1 _2214_ (.A1(_0905_),
    .A2(_1485_),
    .B1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__or4bb_2 _2215_ (.A(_1403_),
    .B(_1487_),
    .C_N(_1406_),
    .D_N(_1405_),
    .X(_1488_));
 sky130_fd_sc_hd__o21ai_2 _2216_ (.A1(_1003_),
    .A2(\demux.state_machine.timeState[1] ),
    .B1(_1102_),
    .Y(_1489_));
 sky130_fd_sc_hd__a21o_1 _2217_ (.A1(_1427_),
    .A2(_1489_),
    .B1(_1310_),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _2218_ (.A(_0917_),
    .B(_0937_),
    .Y(_1491_));
 sky130_fd_sc_hd__o211a_1 _2219_ (.A1(\demux.state_machine.timeState[5] ),
    .A2(_0945_),
    .B1(_1084_),
    .C1(_0891_),
    .X(_1492_));
 sky130_fd_sc_hd__a221o_1 _2220_ (.A1(_0897_),
    .A2(_0912_),
    .B1(_1168_),
    .B2(\demux.state_machine.timeState[1] ),
    .C1(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__a221o_1 _2221_ (.A1(_1491_),
    .A2(_0913_),
    .B1(_0930_),
    .B2(_0876_),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__and3_1 _2222_ (.A(_1273_),
    .B(\demux.state_machine.currentAddress[12] ),
    .C(_1491_),
    .X(_1495_));
 sky130_fd_sc_hd__a32o_1 _2223_ (.A1(_1273_),
    .A2(\demux.state_machine.currentAddress[1] ),
    .A3(_0945_),
    .B1(_0993_),
    .B2(_0985_),
    .X(_1496_));
 sky130_fd_sc_hd__a211o_1 _2224_ (.A1(_0991_),
    .A2(_0993_),
    .B1(_1495_),
    .C1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__o32ai_4 _2225_ (.A1(_1241_),
    .A2(_1290_),
    .A3(_1494_),
    .B1(_1497_),
    .B2(_1416_),
    .Y(_1498_));
 sky130_fd_sc_hd__o211ai_1 _2226_ (.A1(\demux.state_machine.currentAddress[5] ),
    .A2(_0987_),
    .B1(_1384_),
    .C1(_1004_),
    .Y(_1499_));
 sky130_fd_sc_hd__a21o_1 _2227_ (.A1(_1498_),
    .A2(_1499_),
    .B1(_0960_),
    .X(_1500_));
 sky130_fd_sc_hd__and4_1 _2228_ (.A(_1484_),
    .B(_1488_),
    .C(_1490_),
    .D(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_4 _2229_ (.A(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__nor2_1 _2230_ (.A(_0961_),
    .B(_1498_),
    .Y(_0118_));
 sky130_fd_sc_hd__a211oi_2 _2231_ (.A1(_1484_),
    .A2(_1488_),
    .B1(_1490_),
    .C1(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__a21oi_2 _2232_ (.A1(_1427_),
    .A2(_1489_),
    .B1(_1310_),
    .Y(_0120_));
 sky130_fd_sc_hd__or2_1 _2233_ (.A(_0120_),
    .B(_1500_),
    .X(_0121_));
 sky130_fd_sc_hd__nor3b_4 _2234_ (.A(_1502_),
    .B(_0119_),
    .C_N(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2b_2 _2235_ (.A_N(_1425_),
    .B(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__a21oi_1 _2236_ (.A1(_1484_),
    .A2(_1488_),
    .B1(_0118_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor2_2 _2237_ (.A(_0124_),
    .B(_0121_),
    .Y(_0125_));
 sky130_fd_sc_hd__a22o_1 _2238_ (.A1(\internalDataflow.addressLowBusModule.busInputs[38] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[30] ),
    .X(_0126_));
 sky130_fd_sc_hd__nor3b_4 _2239_ (.A(_0120_),
    .B(_1500_),
    .C_N(_0124_),
    .Y(_0127_));
 sky130_fd_sc_hd__a22o_1 _2240_ (.A1(\internalDataflow.addressLowBusModule.busInputs[22] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net8),
    .X(_0128_));
 sky130_fd_sc_hd__or3_2 _2241_ (.A(_0122_),
    .B(_0126_),
    .C(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__and2_2 _2242_ (.A(_0123_),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_1465_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__a21o_1 _2244_ (.A1(_1465_),
    .A2(_1483_),
    .B1(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _2245_ (.A(_1461_),
    .B(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_2 _2246_ (.A(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__nand2_1 _2247_ (.A(_1461_),
    .B(_0132_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_2 _2248_ (.A(_0134_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__a221o_1 _2249_ (.A1(\internalDataflow.stackBusModule.busInputs[45] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[5] ),
    .C1(_1375_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _2250_ (.A1(\internalDataflow.addressLowBusModule.busInputs[29] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[37] ),
    .X(_0138_));
 sky130_fd_sc_hd__a21o_1 _2251_ (.A1(\internalDataflow.stackBusModule.busInputs[37] ),
    .A2(_1371_),
    .B1(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__o21a_1 _2252_ (.A1(_0137_),
    .A2(_0139_),
    .B1(_1372_),
    .X(_0140_));
 sky130_fd_sc_hd__o221a_1 _2253_ (.A1(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(net7),
    .C1(_1431_),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _2254_ (.A1(_1388_),
    .A2(_0140_),
    .B1(_0141_),
    .B2(net47),
    .X(_0142_));
 sky130_fd_sc_hd__a21o_1 _2255_ (.A1(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .A2(_1315_),
    .B1(net48),
    .X(_0143_));
 sky130_fd_sc_hd__a221o_1 _2256_ (.A1(\internalDataflow.accRegToDB[5] ),
    .A2(_1316_),
    .B1(_1314_),
    .B2(net7),
    .C1(_1318_),
    .X(_0144_));
 sky130_fd_sc_hd__a211o_1 _2257_ (.A1(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .A2(_1294_),
    .B1(_0143_),
    .C1(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_2 _2258_ (.A0(_0142_),
    .A1(_0145_),
    .S(_1329_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_1 _2259_ (.A(_1460_),
    .B(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__inv_2 _2260_ (.A(_1257_),
    .Y(_0148_));
 sky130_fd_sc_hd__mux2_2 _2261_ (.A0(_0140_),
    .A1(_0145_),
    .S(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2262_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _2263_ (.A1(\internalDataflow.addressLowBusModule.busInputs[37] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[29] ),
    .X(_0151_));
 sky130_fd_sc_hd__a221o_1 _2264_ (.A1(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net7),
    .C1(_0122_),
    .X(_0152_));
 sky130_fd_sc_hd__o21a_4 _2265_ (.A1(_0151_),
    .A2(_0152_),
    .B1(_0123_),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _2266_ (.A(_1465_),
    .Y(_0154_));
 sky130_fd_sc_hd__mux2_1 _2267_ (.A0(_0150_),
    .A1(_0153_),
    .S(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _2268_ (.A(_0147_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__or2_1 _2269_ (.A(_0147_),
    .B(_0155_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _2270_ (.A(_0156_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a221o_1 _2271_ (.A1(\internalDataflow.stackBusModule.busInputs[44] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[4] ),
    .C1(_1375_),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _2272_ (.A1(\internalDataflow.addressLowBusModule.busInputs[28] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[36] ),
    .X(_0160_));
 sky130_fd_sc_hd__a21o_1 _2273_ (.A1(\internalDataflow.stackBusModule.busInputs[36] ),
    .A2(_1371_),
    .B1(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__o21a_1 _2274_ (.A1(_0159_),
    .A2(_0161_),
    .B1(_1372_),
    .X(_0162_));
 sky130_fd_sc_hd__o221a_1 _2275_ (.A1(\internalDataflow.addressHighBusModule.busInputs[20] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(_0954_),
    .C1(_1431_),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _2276_ (.A1(_1388_),
    .A2(_0162_),
    .B1(_0163_),
    .B2(_1387_),
    .X(_0164_));
 sky130_fd_sc_hd__nor3_1 _2277_ (.A(\demux.reset ),
    .B(\demux.setInterruptFlag ),
    .C(\demux.nmi ),
    .Y(_0165_));
 sky130_fd_sc_hd__a31o_1 _2278_ (.A1(_0983_),
    .A2(_1079_),
    .A3(_0165_),
    .B1(_1260_),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _2279_ (.A1(\internalDataflow.addressLowBusModule.busInputs[20] ),
    .A2(_1315_),
    .B1(_0166_),
    .B2(_1318_),
    .X(_0167_));
 sky130_fd_sc_hd__a221o_1 _2280_ (.A1(\internalDataflow.accRegToDB[4] ),
    .A2(_1316_),
    .B1(_1314_),
    .B2(net6),
    .C1(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__a211o_1 _2281_ (.A1(\internalDataflow.addressHighBusModule.busInputs[20] ),
    .A2(_1294_),
    .B1(net134),
    .C1(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_2 _2282_ (.A0(_0164_),
    .A1(_0169_),
    .S(_1329_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _2283_ (.A(_1460_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_2 _2284_ (.A0(_0162_),
    .A1(_0169_),
    .S(_0148_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _2286_ (.A1(\internalDataflow.addressLowBusModule.busInputs[36] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[28] ),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _2287_ (.A1(\internalDataflow.addressLowBusModule.busInputs[20] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net6),
    .X(_0175_));
 sky130_fd_sc_hd__or3_2 _2288_ (.A(_0122_),
    .B(_0174_),
    .C(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_2 _2289_ (.A(_0123_),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(_0173_),
    .A1(_0177_),
    .S(_0154_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _2291_ (.A(_0171_),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _2292_ (.A(_0171_),
    .B(_0178_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2b_2 _2293_ (.A_N(_0179_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _2294_ (.A(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__a22o_1 _2295_ (.A1(\internalDataflow.accRegToDB[3] ),
    .A2(_1316_),
    .B1(_1318_),
    .B2(\internalDataflow.dataBusModule.busInputs[43] ),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _2296_ (.A1(\internalDataflow.addressHighBusModule.busInputs[19] ),
    .A2(_1294_),
    .B1(_1314_),
    .B2(net5),
    .X(_0184_));
 sky130_fd_sc_hd__a2111o_1 _2297_ (.A1(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .A2(_1315_),
    .B1(_0183_),
    .C1(_0184_),
    .D1(net48),
    .X(_0185_));
 sky130_fd_sc_hd__nor2_1 _2298_ (.A(_1257_),
    .B(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__a21o_1 _2299_ (.A1(_1382_),
    .A2(_1329_),
    .B1(_1387_),
    .X(_0187_));
 sky130_fd_sc_hd__a221o_1 _2300_ (.A1(\internalDataflow.stackBusModule.busInputs[43] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[3] ),
    .C1(_1375_),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _2301_ (.A1(\internalDataflow.addressLowBusModule.busInputs[27] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[35] ),
    .X(_0189_));
 sky130_fd_sc_hd__a21o_1 _2302_ (.A1(\internalDataflow.stackBusModule.busInputs[35] ),
    .A2(_1371_),
    .B1(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__o21ai_2 _2303_ (.A1(_0188_),
    .A2(_0190_),
    .B1(_1372_),
    .Y(_0191_));
 sky130_fd_sc_hd__o221a_1 _2304_ (.A1(\internalDataflow.addressHighBusModule.busInputs[19] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(_0957_),
    .C1(_1431_),
    .X(_0192_));
 sky130_fd_sc_hd__a2bb2o_1 _2305_ (.A1_N(_0187_),
    .A2_N(_0191_),
    .B1(_0192_),
    .B2(net47),
    .X(_0193_));
 sky130_fd_sc_hd__o2bb2a_2 _2306_ (.A1_N(_1326_),
    .A2_N(_0186_),
    .B1(_0193_),
    .B2(_1329_),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _2307_ (.A(_1460_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__a21oi_4 _2308_ (.A1(_1257_),
    .A2(_0191_),
    .B1(_0186_),
    .Y(_0196_));
 sky130_fd_sc_hd__mux2_1 _2309_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _2310_ (.A1(\internalDataflow.addressLowBusModule.busInputs[35] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[27] ),
    .X(_0198_));
 sky130_fd_sc_hd__a221o_1 _2311_ (.A1(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(_0957_),
    .C1(_0122_),
    .X(_0199_));
 sky130_fd_sc_hd__o21a_2 _2312_ (.A1(_0198_),
    .A2(_0199_),
    .B1(_0123_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(_0197_),
    .A1(_0200_),
    .S(_0154_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _2314_ (.A(_0195_),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__nor2_1 _2315_ (.A(_0195_),
    .B(_0201_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_2 _2316_ (.A(_0202_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__a22o_1 _2317_ (.A1(\internalDataflow.accRegToDB[2] ),
    .A2(_1316_),
    .B1(_1318_),
    .B2(\instructionLoader.interruptInjector.processStatusRegIFlag ),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_1 _2318_ (.A1(\internalDataflow.addressHighBusModule.busInputs[18] ),
    .A2(_1294_),
    .B1(_1314_),
    .B2(net4),
    .X(_0206_));
 sky130_fd_sc_hd__a2111o_1 _2319_ (.A1(\internalDataflow.addressLowBusModule.busInputs[18] ),
    .A2(_1315_),
    .B1(_0205_),
    .C1(_0206_),
    .D1(net48),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_1 _2320_ (.A(_1257_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__a221o_1 _2321_ (.A1(\internalDataflow.stackBusModule.busInputs[42] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[2] ),
    .C1(_1375_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _2322_ (.A(\internalDataflow.stackBusModule.busInputs[34] ),
    .B(_1371_),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _2323_ (.A1(\internalDataflow.addressLowBusModule.busInputs[26] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[34] ),
    .X(_0211_));
 sky130_fd_sc_hd__o31a_1 _2324_ (.A1(_0209_),
    .A2(_0210_),
    .A3(_0211_),
    .B1(_1372_),
    .X(_0212_));
 sky130_fd_sc_hd__o221a_1 _2325_ (.A1(\internalDataflow.addressHighBusModule.busInputs[18] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(net4),
    .C1(_1431_),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _2326_ (.A1(_1388_),
    .A2(_0212_),
    .B1(_0213_),
    .B2(net47),
    .X(_0214_));
 sky130_fd_sc_hd__o2bb2a_2 _2327_ (.A1_N(_1326_),
    .A2_N(_0208_),
    .B1(_0214_),
    .B2(_1329_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_2 _2328_ (.A(_1460_),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ba_2 _2329_ (.A1(_0148_),
    .A2(_0212_),
    .B1_N(_0208_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__and3b_1 _2331_ (.A_N(\demux.nmi ),
    .B(_1425_),
    .C(_0122_),
    .X(_0219_));
 sky130_fd_sc_hd__a221o_1 _2332_ (.A1(\internalDataflow.addressLowBusModule.busInputs[34] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[26] ),
    .C1(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__a221o_4 _2333_ (.A1(\internalDataflow.addressLowBusModule.busInputs[18] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net4),
    .C1(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_2 _2334_ (.A0(_0218_),
    .A1(_0221_),
    .S(_0154_),
    .X(_0222_));
 sky130_fd_sc_hd__xor2_4 _2335_ (.A(_0216_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__inv_2 _2336_ (.A(\internalDataflow.stackBusModule.busInputs[40] ),
    .Y(_0224_));
 sky130_fd_sc_hd__or4_1 _2337_ (.A(_0224_),
    .B(_1366_),
    .C(_1368_),
    .D(_1350_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _2338_ (.A(\internalDataflow.accRegToDB[0] ),
    .Y(_0226_));
 sky130_fd_sc_hd__or4_1 _2339_ (.A(_0226_),
    .B(_1366_),
    .C(_1368_),
    .D(_1369_),
    .X(_0227_));
 sky130_fd_sc_hd__o211ai_1 _2340_ (.A1(_1371_),
    .A2(_1367_),
    .B1(_0225_),
    .C1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__and4_1 _2341_ (.A(\internalDataflow.addressLowBusModule.busInputs[24] ),
    .B(_1366_),
    .C(_1341_),
    .D(_1350_),
    .X(_0229_));
 sky130_fd_sc_hd__a221o_1 _2342_ (.A1(\internalDataflow.stackBusModule.busInputs[32] ),
    .A2(_1371_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[32] ),
    .C1(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__o21a_1 _2343_ (.A1(_0228_),
    .A2(_0230_),
    .B1(_1372_),
    .X(_0231_));
 sky130_fd_sc_hd__a32o_1 _2344_ (.A1(net2),
    .A2(_1313_),
    .A3(_1302_),
    .B1(_1316_),
    .B2(\internalDataflow.accRegToDB[0] ),
    .X(_0232_));
 sky130_fd_sc_hd__a32o_1 _2345_ (.A1(\demux.PSR_C ),
    .A2(_1317_),
    .A3(_1302_),
    .B1(_1294_),
    .B2(\internalDataflow.addressHighBusModule.busInputs[16] ),
    .X(_0233_));
 sky130_fd_sc_hd__a2111o_1 _2346_ (.A1(\internalDataflow.addressLowBusModule.busInputs[16] ),
    .A2(_1315_),
    .B1(_0232_),
    .C1(_0233_),
    .D1(net134),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _2347_ (.A(_1256_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__o21a_2 _2348_ (.A1(_0148_),
    .A2(_0231_),
    .B1(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__and4_1 _2350_ (.A(_1265_),
    .B(_1303_),
    .C(_1267_),
    .D(_0122_),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _2351_ (.A1(\internalDataflow.addressLowBusModule.busInputs[32] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[24] ),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _2352_ (.A1(\internalDataflow.addressLowBusModule.busInputs[16] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net2),
    .X(_0240_));
 sky130_fd_sc_hd__or3_4 _2353_ (.A(_0238_),
    .B(_0239_),
    .C(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_1 _2354_ (.A(_0154_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__inv_2 _2355_ (.A(_1460_),
    .Y(_0243_));
 sky130_fd_sc_hd__o211a_1 _2356_ (.A1(_0228_),
    .A2(_0230_),
    .B1(_1372_),
    .C1(_1388_),
    .X(_0244_));
 sky130_fd_sc_hd__o21bai_1 _2357_ (.A1(_1325_),
    .A2(_1428_),
    .B1_N(_1425_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand3_1 _2358_ (.A(_1114_),
    .B(_1423_),
    .C(_1418_),
    .Y(_0246_));
 sky130_fd_sc_hd__or2_1 _2359_ (.A(\internalDataflow.addressHighBusModule.busInputs[16] ),
    .B(_1422_),
    .X(_0247_));
 sky130_fd_sc_hd__o2111a_1 _2360_ (.A1(_1430_),
    .A2(_0245_),
    .B1(_0246_),
    .C1(_0247_),
    .D1(_1387_),
    .X(_0248_));
 sky130_fd_sc_hd__o32ai_4 _2361_ (.A1(_1329_),
    .A2(_0244_),
    .A3(_0248_),
    .B1(_0235_),
    .B2(_1327_),
    .Y(_0249_));
 sky130_fd_sc_hd__nor2_1 _2362_ (.A(_0243_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__a211o_1 _2363_ (.A1(_1465_),
    .A2(_0237_),
    .B1(_0242_),
    .C1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__a32o_1 _2364_ (.A1(_0983_),
    .A2(_0917_),
    .A3(_0987_),
    .B1(_0993_),
    .B2(_0985_),
    .X(_0252_));
 sky130_fd_sc_hd__a221o_1 _2365_ (.A1(_1006_),
    .A2(_0987_),
    .B1(\free_carry_ff.freeCarry ),
    .B2(_0252_),
    .C1(_1364_),
    .X(_0253_));
 sky130_fd_sc_hd__a221o_1 _2366_ (.A1(_1071_),
    .A2(_1244_),
    .B1(_1285_),
    .B2(_1168_),
    .C1(_1444_),
    .X(_0254_));
 sky130_fd_sc_hd__or3b_1 _2367_ (.A(_0254_),
    .B(_1274_),
    .C_N(_1440_),
    .X(_0255_));
 sky130_fd_sc_hd__or4_1 _2368_ (.A(_1121_),
    .B(_1200_),
    .C(_0853_),
    .D(_1174_),
    .X(_0256_));
 sky130_fd_sc_hd__o311a_1 _2369_ (.A1(_0868_),
    .A2(_1143_),
    .A3(_0256_),
    .B1(\demux.PSR_C ),
    .C1(_1006_),
    .X(_0257_));
 sky130_fd_sc_hd__or3b_1 _2370_ (.A(_0255_),
    .B(_0257_),
    .C_N(_1439_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _2371_ (.A(_0998_),
    .B(_0253_),
    .C(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _2372_ (.A(_1465_),
    .B(_0241_),
    .X(_0260_));
 sky130_fd_sc_hd__o211a_1 _2373_ (.A1(_0154_),
    .A2(_0237_),
    .B1(_0260_),
    .C1(_0250_),
    .X(_0261_));
 sky130_fd_sc_hd__a21o_2 _2374_ (.A1(_0251_),
    .A2(_0259_),
    .B1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__a32o_1 _2375_ (.A1(\demux.PSR_Z ),
    .A2(_1317_),
    .A3(_1302_),
    .B1(\internalDataflow.accRegToDB[1] ),
    .B2(_1316_),
    .X(_0263_));
 sky130_fd_sc_hd__a32o_1 _2376_ (.A1(net3),
    .A2(_1313_),
    .A3(_1302_),
    .B1(_1294_),
    .B2(\internalDataflow.addressHighBusModule.busInputs[17] ),
    .X(_0264_));
 sky130_fd_sc_hd__a2111o_1 _2377_ (.A1(\internalDataflow.addressLowBusModule.busInputs[17] ),
    .A2(_1315_),
    .B1(_0263_),
    .C1(_0264_),
    .D1(net48),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _2378_ (.A(_1257_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a22o_1 _2379_ (.A1(\internalDataflow.stackBusModule.busInputs[41] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[1] ),
    .X(_0267_));
 sky130_fd_sc_hd__and2_1 _2380_ (.A(\internalDataflow.stackBusModule.busInputs[33] ),
    .B(_1371_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _2381_ (.A1(\internalDataflow.addressLowBusModule.busInputs[25] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[33] ),
    .X(_0269_));
 sky130_fd_sc_hd__o41ai_2 _2382_ (.A1(_1375_),
    .A2(_0267_),
    .A3(_0268_),
    .A4(_0269_),
    .B1(_1372_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _2383_ (.A(_0187_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o22a_1 _2384_ (.A1(\internalDataflow.addressHighBusModule.busInputs[17] ),
    .A2(_1422_),
    .B1(_1424_),
    .B2(net3),
    .X(_0272_));
 sky130_fd_sc_hd__a31o_1 _2385_ (.A1(net47),
    .A2(_1431_),
    .A3(_0272_),
    .B1(_1329_),
    .X(_0273_));
 sky130_fd_sc_hd__o2bb2a_2 _2386_ (.A1_N(_1326_),
    .A2_N(_0266_),
    .B1(_0271_),
    .B2(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__and2_2 _2387_ (.A(_1460_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__a21oi_4 _2388_ (.A1(_1257_),
    .A2(net44),
    .B1(_0266_),
    .Y(_0276_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(_1467_),
    .A1(_1479_),
    .S(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _2390_ (.A1(\internalDataflow.addressLowBusModule.busInputs[25] ),
    .A2(_0125_),
    .B1(_0127_),
    .B2(net3),
    .X(_0278_));
 sky130_fd_sc_hd__or2b_1 _2391_ (.A(\demux.nmi ),
    .B_N(\demux.reset ),
    .X(_0279_));
 sky130_fd_sc_hd__a32o_1 _2392_ (.A1(_1425_),
    .A2(_0122_),
    .A3(_0279_),
    .B1(net46),
    .B2(\internalDataflow.addressLowBusModule.busInputs[33] ),
    .X(_0280_));
 sky130_fd_sc_hd__a211o_2 _2393_ (.A1(\internalDataflow.addressLowBusModule.busInputs[17] ),
    .A2(_1502_),
    .B1(_0278_),
    .C1(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_2 _2394_ (.A0(_0277_),
    .A1(_0281_),
    .S(_0154_),
    .X(_0282_));
 sky130_fd_sc_hd__xor2_4 _2395_ (.A(_0275_),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _2396_ (.A(_0275_),
    .B(_0282_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_2 _2397_ (.A1(_0262_),
    .A2(_0283_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _2398_ (.A(_0216_),
    .B(_0222_),
    .X(_0286_));
 sky130_fd_sc_hd__a21o_1 _2399_ (.A1(_0223_),
    .A2(_0285_),
    .B1(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _2400_ (.A1(_0204_),
    .A2(_0287_),
    .B1(_0202_),
    .X(_0288_));
 sky130_fd_sc_hd__a21o_1 _2401_ (.A1(_0182_),
    .A2(_0288_),
    .B1(_0179_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _2402_ (.A(_0158_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__and2_1 _2403_ (.A(_0156_),
    .B(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__o21a_1 _2404_ (.A1(_0136_),
    .A2(_0291_),
    .B1(_0134_),
    .X(_0292_));
 sky130_fd_sc_hd__a221o_1 _2405_ (.A1(\internalDataflow.stackBusModule.busInputs[47] ),
    .A2(_1373_),
    .B1(_1374_),
    .B2(\internalDataflow.accRegToDB[7] ),
    .C1(_1375_),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _2406_ (.A1(\internalDataflow.addressLowBusModule.busInputs[31] ),
    .A2(_1377_),
    .B1(_1378_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[39] ),
    .X(_0294_));
 sky130_fd_sc_hd__a211o_1 _2407_ (.A1(\internalDataflow.stackBusModule.busInputs[39] ),
    .A2(_1371_),
    .B1(_0293_),
    .C1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__nand2_2 _2408_ (.A(_1372_),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _2409_ (.A(\internalDataflow.addressHighBusModule.busInputs[23] ),
    .Y(_0297_));
 sky130_fd_sc_hd__nand3_1 _2410_ (.A(_1429_),
    .B(_1422_),
    .C(_1424_),
    .Y(_0298_));
 sky130_fd_sc_hd__o221a_1 _2411_ (.A1(_0297_),
    .A2(_1422_),
    .B1(_1424_),
    .B2(_0968_),
    .C1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(_0296_),
    .A1(_0299_),
    .S(net47),
    .X(_0300_));
 sky130_fd_sc_hd__inv_2 _2413_ (.A(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__a22o_1 _2414_ (.A1(\internalDataflow.accRegToDB[7] ),
    .A2(_1316_),
    .B1(_1318_),
    .B2(\demux.PSR_N ),
    .X(_0302_));
 sky130_fd_sc_hd__a221o_1 _2415_ (.A1(\internalDataflow.addressHighBusModule.busInputs[23] ),
    .A2(_1294_),
    .B1(_1314_),
    .B2(_1012_),
    .C1(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a211o_1 _2416_ (.A1(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .A2(_1315_),
    .B1(_0303_),
    .C1(net48),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_4 _2417_ (.A0(_0301_),
    .A1(_0304_),
    .S(_1329_),
    .X(_0305_));
 sky130_fd_sc_hd__nand2_1 _2418_ (.A(_1460_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _2419_ (.A(_1257_),
    .B(_0304_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21oi_4 _2420_ (.A1(_1257_),
    .A2(_0296_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(_1468_),
    .A1(_1480_),
    .S(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _2422_ (.A1(\internalDataflow.addressLowBusModule.busInputs[39] ),
    .A2(net46),
    .B1(_0125_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[31] ),
    .X(_0310_));
 sky130_fd_sc_hd__a221o_1 _2423_ (.A1(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .A2(_1502_),
    .B1(_0127_),
    .B2(net9),
    .C1(_0122_),
    .X(_0311_));
 sky130_fd_sc_hd__o21a_2 _2424_ (.A1(_0310_),
    .A2(_0311_),
    .B1(_0123_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_1 _2425_ (.A(_1465_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21o_1 _2426_ (.A1(_1465_),
    .A2(_0309_),
    .B1(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__or2_2 _2427_ (.A(_0306_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _2428_ (.A(_0292_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__and2_1 _2429_ (.A(_0306_),
    .B(_0314_),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _2430_ (.A(_0292_),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__o21ai_2 _2431_ (.A1(_0868_),
    .A2(_1143_),
    .B1(_1007_),
    .Y(_0319_));
 sky130_fd_sc_hd__nor2_1 _2432_ (.A(_1325_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__nand2_2 _2433_ (.A(\internalDataflow.dataBusModule.busInputs[43] ),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _2434_ (.A(net14),
    .Y(_0322_));
 sky130_fd_sc_hd__nor2_4 _2435_ (.A(_1273_),
    .B(_1325_),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _2436_ (.A(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_2 _2437_ (.A(_1325_),
    .B(_0319_),
    .X(_0325_));
 sky130_fd_sc_hd__o311a_1 _2438_ (.A1(_0866_),
    .A2(_0844_),
    .A3(_0324_),
    .B1(_0325_),
    .C1(\demux.PSR_V ),
    .X(_0326_));
 sky130_fd_sc_hd__o21a_1 _2439_ (.A1(_1168_),
    .A2(_1094_),
    .B1(_0983_),
    .X(_0327_));
 sky130_fd_sc_hd__a21oi_1 _2440_ (.A1(_1008_),
    .A2(_0873_),
    .B1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__or2_1 _2441_ (.A(_1325_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(_1482_),
    .A1(_0326_),
    .S(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__a31o_1 _2443_ (.A1(_0322_),
    .A2(net89),
    .A3(_0999_),
    .B1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__a41o_1 _2444_ (.A1(_0316_),
    .A2(_0318_),
    .A3(_0320_),
    .A4(_0321_),
    .B1(_0331_),
    .X(\internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ));
 sky130_fd_sc_hd__clkbuf_4 _2445_ (.A(_1303_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _2446_ (.A(_0332_),
    .B(_0327_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _2447_ (.A(\demux.state_machine.timeState[5] ),
    .B(\demux.setInterruptFlag ),
    .C(_1079_),
    .X(_0334_));
 sky130_fd_sc_hd__a21o_1 _2448_ (.A1(_0982_),
    .A2(_0334_),
    .B1(_0819_),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _2449_ (.A(_0332_),
    .B(_0327_),
    .Y(_0336_));
 sky130_fd_sc_hd__and2_1 _2450_ (.A(\internalDataflow.dataBusModule.busInputs[43] ),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o21ai_1 _2451_ (.A1(_0842_),
    .A2(_0908_),
    .B1(_0323_),
    .Y(_0338_));
 sky130_fd_sc_hd__mux2_1 _2452_ (.A0(_0335_),
    .A1(_0337_),
    .S(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__a21o_1 _2453_ (.A1(_0196_),
    .A2(_0333_),
    .B1(_0339_),
    .X(\internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ));
 sky130_fd_sc_hd__nand2_1 _2454_ (.A(_0982_),
    .B(_0334_),
    .Y(_0340_));
 sky130_fd_sc_hd__nor2_1 _2455_ (.A(_0981_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__a21oi_1 _2456_ (.A1(_1008_),
    .A2(_0846_),
    .B1(_0334_),
    .Y(_0342_));
 sky130_fd_sc_hd__o211a_1 _2457_ (.A1(_1325_),
    .A2(_0342_),
    .B1(_0336_),
    .C1(\instructionLoader.interruptInjector.processStatusRegIFlag ),
    .X(_0343_));
 sky130_fd_sc_hd__a211o_1 _2458_ (.A1(_0217_),
    .A2(_0333_),
    .B1(_0341_),
    .C1(_0343_),
    .X(\internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ));
 sky130_fd_sc_hd__or4_1 _2459_ (.A(_0149_),
    .B(_0172_),
    .C(_0196_),
    .D(_0217_),
    .X(_0344_));
 sky130_fd_sc_hd__a221o_1 _2460_ (.A1(_0983_),
    .A2(_1150_),
    .B1(_1237_),
    .B2(_1002_),
    .C1(_0918_),
    .X(_0345_));
 sky130_fd_sc_hd__a211o_1 _2461_ (.A1(_1002_),
    .A2(_1353_),
    .B1(_1239_),
    .C1(_1238_),
    .X(_0346_));
 sky130_fd_sc_hd__a211o_1 _2462_ (.A1(_1008_),
    .A2(_0840_),
    .B1(_0345_),
    .C1(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__o21a_1 _2463_ (.A1(_1359_),
    .A2(_0347_),
    .B1(_0332_),
    .X(_0348_));
 sky130_fd_sc_hd__or4b_1 _2464_ (.A(_1482_),
    .B(_0344_),
    .C(_0308_),
    .D_N(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _2465_ (.A(\demux.PSR_Z ),
    .B(_0336_),
    .Y(_0350_));
 sky130_fd_sc_hd__o2bb2a_1 _2466_ (.A1_N(_0276_),
    .A2_N(_0333_),
    .B1(_0348_),
    .B2(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__o31ai_1 _2467_ (.A1(_0276_),
    .A2(_0236_),
    .A3(_0349_),
    .B1(_0351_),
    .Y(\internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ));
 sky130_fd_sc_hd__o21a_1 _2468_ (.A1(_1274_),
    .A2(_1454_),
    .B1(_0332_),
    .X(_0352_));
 sky130_fd_sc_hd__o31a_1 _2469_ (.A1(_1097_),
    .A2(_1298_),
    .A3(_1358_),
    .B1(_1007_),
    .X(_0353_));
 sky130_fd_sc_hd__a211o_1 _2470_ (.A1(_1168_),
    .A2(_1441_),
    .B1(_1330_),
    .C1(_1267_),
    .X(_0354_));
 sky130_fd_sc_hd__o21a_1 _2471_ (.A1(_0847_),
    .A2(_0868_),
    .B1(_1006_),
    .X(_0355_));
 sky130_fd_sc_hd__a221o_1 _2472_ (.A1(_1071_),
    .A2(_1285_),
    .B1(_1409_),
    .B2(_1102_),
    .C1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _2473_ (.A(_1273_),
    .B(_1390_),
    .Y(_0357_));
 sky130_fd_sc_hd__a2111o_1 _2474_ (.A1(_1007_),
    .A2(_1249_),
    .B1(_1444_),
    .C1(_0356_),
    .D1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__or4_2 _2475_ (.A(_1474_),
    .B(_0353_),
    .C(_0354_),
    .D(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_2 _2476_ (.A(_1462_),
    .B(_1290_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ai_4 _2477_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_1478_),
    .Y(_0361_));
 sky130_fd_sc_hd__a31o_1 _2478_ (.A1(_0315_),
    .A2(_0318_),
    .A3(_0321_),
    .B1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a21oi_1 _2479_ (.A1(_0909_),
    .A2(_0852_),
    .B1(_1076_),
    .Y(_0363_));
 sky130_fd_sc_hd__o31a_4 _2480_ (.A1(_1121_),
    .A2(_1144_),
    .A3(_0363_),
    .B1(_0323_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _2481_ (.A(_0250_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21oi_1 _2482_ (.A1(_0204_),
    .A2(_0287_),
    .B1(_0202_),
    .Y(_0366_));
 sky130_fd_sc_hd__xor2_4 _2483_ (.A(_0262_),
    .B(_0283_),
    .X(_0367_));
 sky130_fd_sc_hd__xor2_4 _2484_ (.A(_0223_),
    .B(_0285_),
    .X(_0368_));
 sky130_fd_sc_hd__o22ai_2 _2485_ (.A1(_0204_),
    .A2(_0287_),
    .B1(_0367_),
    .B2(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__a21oi_1 _2486_ (.A1(_0366_),
    .A2(_0369_),
    .B1(_0181_),
    .Y(_0370_));
 sky130_fd_sc_hd__o21ai_1 _2487_ (.A1(_0179_),
    .A2(_0370_),
    .B1(_0158_),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_2 _2488_ (.A1(_0156_),
    .A2(_0371_),
    .B1(_0136_),
    .X(_0372_));
 sky130_fd_sc_hd__nand3_1 _2489_ (.A(_0136_),
    .B(_0156_),
    .C(_0371_),
    .Y(_0373_));
 sky130_fd_sc_hd__or3_1 _2490_ (.A(_0158_),
    .B(_0179_),
    .C(_0370_),
    .X(_0374_));
 sky130_fd_sc_hd__and2_2 _2491_ (.A(_0371_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__a21o_2 _2492_ (.A1(_0372_),
    .A2(_0373_),
    .B1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__inv_2 _2493_ (.A(_0317_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_2 _2494_ (.A(_0315_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _2495_ (.A1(_0134_),
    .A2(_0372_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__nand3_2 _2496_ (.A(_0134_),
    .B(_0372_),
    .C(_0378_),
    .Y(_0380_));
 sky130_fd_sc_hd__and3_1 _2497_ (.A(_0376_),
    .B(_0379_),
    .C(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _2498_ (.A(\internalDataflow.dataBusModule.busInputs[43] ),
    .B(_0320_),
    .X(_0382_));
 sky130_fd_sc_hd__a31o_2 _2499_ (.A1(_0134_),
    .A2(_0315_),
    .A3(_0372_),
    .B1(_0317_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(_0382_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__o2bb2a_2 _2501_ (.A1_N(_0362_),
    .A2_N(_0365_),
    .B1(_0381_),
    .B2(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__and3b_1 _2502_ (.A_N(_0352_),
    .B(\demux.PSR_C ),
    .C(_0336_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ai_1 _2503_ (.A1(_0907_),
    .A2(_0921_),
    .B1(_0323_),
    .Y(_0387_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(_0335_),
    .A1(_0386_),
    .S(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a221o_1 _2505_ (.A1(_0236_),
    .A2(_0333_),
    .B1(_0352_),
    .B2(_0385_),
    .C1(_0388_),
    .X(\internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ));
 sky130_fd_sc_hd__inv_2 _2506_ (.A(\internalDataflow.stackBusModule.busInputs[32] ),
    .Y(_0389_));
 sky130_fd_sc_hd__o21a_1 _2507_ (.A1(_0831_),
    .A2(_1108_),
    .B1(_1008_),
    .X(_0390_));
 sky130_fd_sc_hd__o21a_1 _2508_ (.A1(_0910_),
    .A2(_1097_),
    .B1(_1002_),
    .X(_0391_));
 sky130_fd_sc_hd__o21a_4 _2509_ (.A1(_0390_),
    .A2(_0391_),
    .B1(_0332_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(_0389_),
    .A1(_0249_),
    .S(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _2511_ (.A(_0393_),
    .Y(_0026_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(net104),
    .A1(_0274_),
    .S(_0392_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_0394_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(net93),
    .A1(_0215_),
    .S(_0392_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_0395_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(net106),
    .A1(_0194_),
    .S(_0392_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_0396_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(net114),
    .A1(_0170_),
    .S(_0392_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_0397_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(net99),
    .A1(_0146_),
    .S(_0392_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_0398_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net109),
    .A1(_1434_),
    .S(_0392_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_0399_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net131),
    .A1(_0305_),
    .S(_0392_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(_0400_),
    .X(_0033_));
 sky130_fd_sc_hd__o31a_1 _2526_ (.A1(_1121_),
    .A2(_1144_),
    .A3(_0873_),
    .B1(_1008_),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _2527_ (.A(_1452_),
    .B(_1475_),
    .C(_0354_),
    .D(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__o31ai_2 _2528_ (.A1(_0358_),
    .A2(_0360_),
    .A3(_0402_),
    .B1(_1478_),
    .Y(_0403_));
 sky130_fd_sc_hd__and2b_1 _2529_ (.A_N(_0261_),
    .B(_0251_),
    .X(_0404_));
 sky130_fd_sc_hd__xor2_1 _2530_ (.A(_0404_),
    .B(_0259_),
    .X(_0405_));
 sky130_fd_sc_hd__inv_2 _2531_ (.A(_0361_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_2 _2532_ (.A(_1271_),
    .B(_0323_),
    .Y(_0407_));
 sky130_fd_sc_hd__and3_2 _2533_ (.A(_1007_),
    .B(_0332_),
    .C(_1131_),
    .X(_0408_));
 sky130_fd_sc_hd__and3_1 _2534_ (.A(_1007_),
    .B(_1303_),
    .C(_1271_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_2 _2535_ (.A(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__a221o_1 _2536_ (.A1(_0275_),
    .A2(_0364_),
    .B1(_0408_),
    .B2(_0251_),
    .C1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__and3_2 _2537_ (.A(_1007_),
    .B(_1303_),
    .C(_1202_),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _2538_ (.A(_0404_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _2539_ (.A1(_0261_),
    .A2(_0407_),
    .B1(_0411_),
    .B2(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__a221o_1 _2540_ (.A1(net80),
    .A2(_0403_),
    .B1(_0405_),
    .B2(_0406_),
    .C1(_0414_),
    .X(_0034_));
 sky130_fd_sc_hd__o21a_1 _2541_ (.A1(_0275_),
    .A2(_0282_),
    .B1(_0408_),
    .X(_0415_));
 sky130_fd_sc_hd__a221o_1 _2542_ (.A1(_0216_),
    .A2(_0364_),
    .B1(_0412_),
    .B2(_0283_),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__a211o_1 _2543_ (.A1(_0284_),
    .A2(_0410_),
    .B1(_0416_),
    .C1(_0406_),
    .X(_0417_));
 sky130_fd_sc_hd__or3_1 _2544_ (.A(_0288_),
    .B(_0321_),
    .C(_0369_),
    .X(_0418_));
 sky130_fd_sc_hd__xor2_1 _2545_ (.A(_0367_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _2546_ (.A(_0406_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__a22o_1 _2547_ (.A1(net96),
    .A2(net45),
    .B1(_0417_),
    .B2(_0420_),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _2548_ (.A(_0223_),
    .B(_0412_),
    .X(_0421_));
 sky130_fd_sc_hd__o21a_1 _2549_ (.A1(_0216_),
    .A2(_0222_),
    .B1(_0408_),
    .X(_0422_));
 sky130_fd_sc_hd__a221o_1 _2550_ (.A1(_0195_),
    .A2(_0364_),
    .B1(_0410_),
    .B2(_0286_),
    .C1(_0406_),
    .X(_0423_));
 sky130_fd_sc_hd__o32a_1 _2551_ (.A1(_0421_),
    .A2(_0422_),
    .A3(_0423_),
    .B1(_0368_),
    .B2(_0361_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _2552_ (.A(_1466_),
    .B(_0325_),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _2553_ (.A(_0367_),
    .B(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__nor2_1 _2554_ (.A(_0367_),
    .B(_0425_),
    .Y(_0427_));
 sky130_fd_sc_hd__or4_1 _2555_ (.A(_0288_),
    .B(_0369_),
    .C(_0426_),
    .D(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__xnor2_1 _2556_ (.A(_0368_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(_0424_),
    .A1(_0429_),
    .S(_0382_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(_0430_),
    .A1(\internalDataflow.addressLowBusModule.busInputs[26] ),
    .S(net45),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _2559_ (.A(_0431_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(_0367_),
    .A1(_0425_),
    .S(_0368_),
    .X(_0432_));
 sky130_fd_sc_hd__nor2_1 _2561_ (.A(_0427_),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a21oi_1 _2562_ (.A1(_0204_),
    .A2(_0287_),
    .B1(_0361_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _2563_ (.A(_0204_),
    .B(_0287_),
    .X(_0435_));
 sky130_fd_sc_hd__o211a_1 _2564_ (.A1(_0418_),
    .A2(_0433_),
    .B1(_0434_),
    .C1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(_1131_),
    .B(_0323_),
    .Y(_0437_));
 sky130_fd_sc_hd__a2bb2o_1 _2566_ (.A1_N(_0203_),
    .A2_N(_0437_),
    .B1(_0364_),
    .B2(_0171_),
    .X(_0438_));
 sky130_fd_sc_hd__a211o_1 _2567_ (.A1(_0204_),
    .A2(_0412_),
    .B1(_0410_),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__o211a_1 _2568_ (.A1(_0202_),
    .A2(_0407_),
    .B1(_0439_),
    .C1(_0361_),
    .X(_0440_));
 sky130_fd_sc_hd__a211o_1 _2569_ (.A1(net82),
    .A2(net45),
    .B1(_0436_),
    .C1(_0440_),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _2570_ (.A(_0181_),
    .B(_0366_),
    .C(_0369_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _2571_ (.A(_0182_),
    .B(_0288_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _2572_ (.A1(_0181_),
    .A2(_0366_),
    .B1(_0361_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _2573_ (.A(_1202_),
    .B(_0323_),
    .Y(_0444_));
 sky130_fd_sc_hd__nor2_1 _2574_ (.A(_0181_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a221o_1 _2575_ (.A1(_0147_),
    .A2(_0364_),
    .B1(_0408_),
    .B2(_0180_),
    .C1(_0410_),
    .X(_0446_));
 sky130_fd_sc_hd__o22a_1 _2576_ (.A1(_0179_),
    .A2(_0407_),
    .B1(_0445_),
    .B2(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__a21oi_1 _2577_ (.A1(_0442_),
    .A2(_0443_),
    .B1(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__o2bb2a_1 _2578_ (.A1_N(\internalDataflow.addressLowBusModule.busInputs[28] ),
    .A2_N(net45),
    .B1(_0448_),
    .B2(_0382_),
    .X(_0449_));
 sky130_fd_sc_hd__o31ai_1 _2579_ (.A1(_0321_),
    .A2(_0370_),
    .A3(_0441_),
    .B1(_0449_),
    .Y(_0038_));
 sky130_fd_sc_hd__a41oi_4 _2580_ (.A1(_0376_),
    .A2(_0379_),
    .A3(_0380_),
    .A4(_0383_),
    .B1(_0375_),
    .Y(_0450_));
 sky130_fd_sc_hd__a31o_1 _2581_ (.A1(_0375_),
    .A2(_0381_),
    .A3(_0383_),
    .B1(_0321_),
    .X(_0451_));
 sky130_fd_sc_hd__or2_1 _2582_ (.A(_0158_),
    .B(_0289_),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _2583_ (.A(_0156_),
    .B(_0410_),
    .Y(_0453_));
 sky130_fd_sc_hd__a32o_1 _2584_ (.A1(_1434_),
    .A2(_1460_),
    .A3(_0364_),
    .B1(_0408_),
    .B2(_0157_),
    .X(_0454_));
 sky130_fd_sc_hd__a211o_1 _2585_ (.A1(_0158_),
    .A2(_0412_),
    .B1(_0410_),
    .C1(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__a32o_1 _2586_ (.A1(_0290_),
    .A2(_0406_),
    .A3(_0452_),
    .B1(_0453_),
    .B2(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__a22oi_1 _2587_ (.A1(net112),
    .A2(net45),
    .B1(_0456_),
    .B2(_0321_),
    .Y(_0457_));
 sky130_fd_sc_hd__o21ai_1 _2588_ (.A1(_0450_),
    .A2(_0451_),
    .B1(_0457_),
    .Y(_0039_));
 sky130_fd_sc_hd__o21ai_1 _2589_ (.A1(_0136_),
    .A2(_0291_),
    .B1(_0406_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_1 _2590_ (.A1(_0136_),
    .A2(_0291_),
    .B1(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _2591_ (.A(_0136_),
    .B(_0444_),
    .Y(_0460_));
 sky130_fd_sc_hd__a32o_1 _2592_ (.A1(_1460_),
    .A2(_0305_),
    .A3(_0364_),
    .B1(_0408_),
    .B2(_0135_),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _2593_ (.A(_0134_),
    .B(_0410_),
    .Y(_0462_));
 sky130_fd_sc_hd__o311a_1 _2594_ (.A1(_0410_),
    .A2(_0460_),
    .A3(_0461_),
    .B1(_0462_),
    .C1(_0361_),
    .X(_0463_));
 sky130_fd_sc_hd__or3_1 _2595_ (.A(_0382_),
    .B(_0459_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__a21boi_1 _2596_ (.A1(_0134_),
    .A2(_0372_),
    .B1_N(_0378_),
    .Y(_0465_));
 sky130_fd_sc_hd__and3b_1 _2597_ (.A_N(_0378_),
    .B(_0372_),
    .C(_0134_),
    .X(_0466_));
 sky130_fd_sc_hd__nor2_1 _2598_ (.A(_1466_),
    .B(_0325_),
    .Y(_0467_));
 sky130_fd_sc_hd__o2111a_1 _2599_ (.A1(_0465_),
    .A2(_0466_),
    .B1(_0383_),
    .C1(_0467_),
    .D1(_0376_),
    .X(_0468_));
 sky130_fd_sc_hd__nand3_1 _2600_ (.A(_0375_),
    .B(_0372_),
    .C(_0373_),
    .Y(_0469_));
 sky130_fd_sc_hd__o211a_1 _2601_ (.A1(_0450_),
    .A2(_0468_),
    .B1(_0469_),
    .C1(_0376_),
    .X(_0470_));
 sky130_fd_sc_hd__a211o_1 _2602_ (.A1(_0376_),
    .A2(_0469_),
    .B1(_0468_),
    .C1(_0450_),
    .X(_0471_));
 sky130_fd_sc_hd__or3b_1 _2603_ (.A(_0470_),
    .B(_0321_),
    .C_N(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _2604_ (.A1(net129),
    .A2(net45),
    .B1(_0464_),
    .B2(_0472_),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _2605_ (.A(_0425_),
    .B(_0469_),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_1 _2606_ (.A(_0465_),
    .B(_0466_),
    .Y(_0474_));
 sky130_fd_sc_hd__a31o_1 _2607_ (.A1(_0376_),
    .A2(_0383_),
    .A3(_0473_),
    .B1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_1 _2608_ (.A(_0292_),
    .B(_0378_),
    .Y(_0476_));
 sky130_fd_sc_hd__a21o_1 _2609_ (.A1(_0292_),
    .A2(_0378_),
    .B1(_0361_),
    .X(_0477_));
 sky130_fd_sc_hd__nand2_1 _2610_ (.A(_0259_),
    .B(_0364_),
    .Y(_0478_));
 sky130_fd_sc_hd__o221a_1 _2611_ (.A1(_0378_),
    .A2(_0444_),
    .B1(_0437_),
    .B2(_0317_),
    .C1(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(_0315_),
    .A1(_0479_),
    .S(_0407_),
    .X(_0480_));
 sky130_fd_sc_hd__o21a_1 _2613_ (.A1(_0476_),
    .A2(_0477_),
    .B1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(_0475_),
    .A1(_0481_),
    .S(_0321_),
    .X(_0482_));
 sky130_fd_sc_hd__a21bo_1 _2615_ (.A1(net83),
    .A2(net45),
    .B1_N(_0482_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _2616_ (.A(_1406_),
    .B(_1405_),
    .Y(_0483_));
 sky130_fd_sc_hd__a211o_1 _2617_ (.A1(_1001_),
    .A2(_0911_),
    .B1(_1391_),
    .C1(_0934_),
    .X(_0484_));
 sky130_fd_sc_hd__a211o_1 _2618_ (.A1(_1001_),
    .A2(_0848_),
    .B1(_1395_),
    .C1(_1396_),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _2619_ (.A1(_1491_),
    .A2(_1150_),
    .B1(_1285_),
    .B2(_1259_),
    .X(_0486_));
 sky130_fd_sc_hd__a211o_1 _2620_ (.A1(_1001_),
    .A2(_1094_),
    .B1(_1394_),
    .C1(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__or4_1 _2621_ (.A(_0483_),
    .B(_0484_),
    .C(_0485_),
    .D(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__a221o_1 _2622_ (.A1(_0877_),
    .A2(_0921_),
    .B1(_1244_),
    .B2(_0839_),
    .C1(_1399_),
    .X(_0489_));
 sky130_fd_sc_hd__or3_1 _2623_ (.A(_1384_),
    .B(_1486_),
    .C(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__or2_1 _2624_ (.A(_0879_),
    .B(_1400_),
    .X(_0491_));
 sky130_fd_sc_hd__or3_1 _2625_ (.A(\demux.state_machine.timeState[3] ),
    .B(_1285_),
    .C(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__or3_1 _2626_ (.A(_1007_),
    .B(_0936_),
    .C(_1400_),
    .X(_0493_));
 sky130_fd_sc_hd__or2_1 _2627_ (.A(_1001_),
    .B(_0491_),
    .X(_0494_));
 sky130_fd_sc_hd__o21a_1 _2628_ (.A1(_0983_),
    .A2(_0494_),
    .B1(_0913_),
    .X(_0495_));
 sky130_fd_sc_hd__a221o_1 _2629_ (.A1(_1079_),
    .A2(_0492_),
    .B1(_0493_),
    .B2(_1102_),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__a2111o_1 _2630_ (.A1(_0905_),
    .A2(_1441_),
    .B1(_0488_),
    .C1(_0490_),
    .D1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__a221o_1 _2631_ (.A1(_1435_),
    .A2(_0993_),
    .B1(_1244_),
    .B2(\demux.state_machine.currentAddress[7] ),
    .C1(_0994_),
    .X(_0498_));
 sky130_fd_sc_hd__a21oi_1 _2632_ (.A1(\demux.state_machine.currentAddress[6] ),
    .A2(_1441_),
    .B1(_0982_),
    .Y(_0499_));
 sky130_fd_sc_hd__or3b_1 _2633_ (.A(_0498_),
    .B(_1495_),
    .C_N(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a221o_1 _2634_ (.A1(_0985_),
    .A2(_1244_),
    .B1(_1285_),
    .B2(_0987_),
    .C1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_4 _2635_ (.A(_0999_),
    .B(_0497_),
    .C(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__inv_2 _2636_ (.A(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21o_1 _2637_ (.A1(net97),
    .A2(_0503_),
    .B1(_0241_),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _2638_ (.A1(net79),
    .A2(_0503_),
    .B1(_0281_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _2639_ (.A1(net75),
    .A2(_0503_),
    .B1(_0221_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(net122),
    .A1(_0200_),
    .S(_0502_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_0504_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(net28),
    .A1(_0177_),
    .S(_0502_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(_0505_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(net111),
    .A1(_0153_),
    .S(_0502_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(_0506_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(net123),
    .A1(_0130_),
    .S(_0502_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _2647_ (.A(_0507_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(net31),
    .A1(_0312_),
    .S(_0502_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _2649_ (.A(_0508_),
    .X(_0049_));
 sky130_fd_sc_hd__o31a_1 _2650_ (.A1(_0868_),
    .A2(_0870_),
    .A3(_1202_),
    .B1(_1002_),
    .X(_0509_));
 sky130_fd_sc_hd__o31a_1 _2651_ (.A1(_0839_),
    .A2(_1058_),
    .A3(_1128_),
    .B1(_1008_),
    .X(_0510_));
 sky130_fd_sc_hd__o31a_4 _2652_ (.A1(_0345_),
    .A2(_0509_),
    .A3(_0510_),
    .B1(_0332_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(_0226_),
    .A1(_0249_),
    .S(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__inv_2 _2654_ (.A(_0512_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(\internalDataflow.accRegToDB[1] ),
    .A1(_0274_),
    .S(_0511_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _2656_ (.A(_0513_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(\internalDataflow.accRegToDB[2] ),
    .A1(_0215_),
    .S(_0511_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _2658_ (.A(_0514_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(\internalDataflow.accRegToDB[3] ),
    .A1(_0194_),
    .S(_0511_),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_0515_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(\internalDataflow.accRegToDB[4] ),
    .A1(_0170_),
    .S(_0511_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_0516_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(\internalDataflow.accRegToDB[5] ),
    .A1(_0146_),
    .S(_0511_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_0517_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(\internalDataflow.accRegToDB[6] ),
    .A1(_1434_),
    .S(_0511_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_0518_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(\internalDataflow.accRegToDB[7] ),
    .A1(_0305_),
    .S(_0511_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _2668_ (.A(_0519_),
    .X(_0057_));
 sky130_fd_sc_hd__nand2_1 _2669_ (.A(_0939_),
    .B(_0940_),
    .Y(_0520_));
 sky130_fd_sc_hd__o22ai_4 _2670_ (.A1(\demux.nmi ),
    .A2(\instructionLoader.interruptInjector.irqGenerated ),
    .B1(net43),
    .B2(\instructionLoader.interruptInjector.resetDetected ),
    .Y(_0521_));
 sky130_fd_sc_hd__o21ai_2 _2671_ (.A1(_0520_),
    .A2(_0324_),
    .B1(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__o21a_1 _2672_ (.A1(_1469_),
    .A2(_0898_),
    .B1(_0877_),
    .X(_0523_));
 sky130_fd_sc_hd__o31a_1 _2673_ (.A1(_1005_),
    .A2(_0936_),
    .A3(_0523_),
    .B1(_0905_),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _2674_ (.A(_1394_),
    .B(_1398_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _2675_ (.A(\demux.state_machine.timeState[5] ),
    .B(\demux.state_machine.timeState[3] ),
    .X(_0526_));
 sky130_fd_sc_hd__a221o_1 _2676_ (.A1(_1071_),
    .A2(_0491_),
    .B1(_0526_),
    .B2(_1079_),
    .C1(_1411_),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _2677_ (.A(_1392_),
    .B(_0525_),
    .C(_0490_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__nand2_1 _2678_ (.A(_1005_),
    .B(_0985_),
    .Y(_0529_));
 sky130_fd_sc_hd__and2_1 _2679_ (.A(_0877_),
    .B(_0933_),
    .X(_0530_));
 sky130_fd_sc_hd__o21ai_1 _2680_ (.A1(_1005_),
    .A2(_0530_),
    .B1(\demux.state_machine.currentAddress[7] ),
    .Y(_0531_));
 sky130_fd_sc_hd__a31oi_1 _2681_ (.A1(_0529_),
    .A2(_0499_),
    .A3(_0531_),
    .B1(_0961_),
    .Y(_0532_));
 sky130_fd_sc_hd__o31a_2 _2682_ (.A1(_0483_),
    .A2(_0524_),
    .A3(_0528_),
    .B1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__nand2_1 _2683_ (.A(_0521_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__buf_2 _2684_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_4 _2685_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__inv_2 _2686_ (.A(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_2 _2687_ (.A(_0522_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__a21bo_1 _2688_ (.A1(_1001_),
    .A2(_0933_),
    .B1_N(_1414_),
    .X(_0539_));
 sky130_fd_sc_hd__o211a_1 _2689_ (.A1(\demux.state_machine.currentAddress[6] ),
    .A2(\demux.state_machine.currentAddress[7] ),
    .B1(_0539_),
    .C1(_1273_),
    .X(_0540_));
 sky130_fd_sc_hd__or3_1 _2690_ (.A(_0934_),
    .B(_1385_),
    .C(_1412_),
    .X(_0541_));
 sky130_fd_sc_hd__o221ai_4 _2691_ (.A1(_0982_),
    .A2(_0540_),
    .B1(_0541_),
    .B2(_1290_),
    .C1(_0999_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _2692_ (.A(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__clkbuf_4 _2693_ (.A(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\internalDataflow.addressLowBusModule.busInputs[16] ),
    .A1(_0241_),
    .S(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__xnor2_1 _2695_ (.A(_0538_),
    .B(_0545_),
    .Y(_0058_));
 sky130_fd_sc_hd__nor2_4 _2696_ (.A(_0538_),
    .B(_0543_),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _2697_ (.A(\internalDataflow.addressLowBusModule.busInputs[16] ),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _2698_ (.A(\internalDataflow.addressLowBusModule.busInputs[17] ),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_1 _2699_ (.A1(_0521_),
    .A2(_0533_),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__and3_1 _2700_ (.A(_0548_),
    .B(_0521_),
    .C(_0533_),
    .X(_0550_));
 sky130_fd_sc_hd__nor2_1 _2701_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__xnor2_1 _2702_ (.A(_0547_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__clkbuf_4 _2703_ (.A(_0542_),
    .X(_0553_));
 sky130_fd_sc_hd__and2_2 _2704_ (.A(_0538_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_4 _2705_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _2706_ (.A(_0536_),
    .X(_0556_));
 sky130_fd_sc_hd__buf_2 _2707_ (.A(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_4 _2708_ (.A(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__and2_1 _2709_ (.A(_0522_),
    .B(_0557_),
    .X(_0559_));
 sky130_fd_sc_hd__a21o_1 _2710_ (.A1(_0241_),
    .A2(_0558_),
    .B1(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__and2_1 _2711_ (.A(_0281_),
    .B(_0241_),
    .X(_0561_));
 sky130_fd_sc_hd__nor2_1 _2712_ (.A(_0281_),
    .B(_0241_),
    .Y(_0562_));
 sky130_fd_sc_hd__nor2_1 _2713_ (.A(_0561_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__xnor2_1 _2714_ (.A(_0560_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(_0553_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__a221o_1 _2716_ (.A1(_0546_),
    .A2(_0552_),
    .B1(_0555_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[17] ),
    .C1(_0565_),
    .X(_0059_));
 sky130_fd_sc_hd__o22a_1 _2717_ (.A1(_0559_),
    .A2(_0561_),
    .B1(_0562_),
    .B2(_0537_),
    .X(_0566_));
 sky130_fd_sc_hd__xor2_1 _2718_ (.A(_0221_),
    .B(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__xor2_1 _2719_ (.A(\internalDataflow.addressLowBusModule.busInputs[18] ),
    .B(_0535_),
    .X(_0568_));
 sky130_fd_sc_hd__o21bai_2 _2720_ (.A1(_0547_),
    .A2(_0550_),
    .B1_N(_0549_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__or2_1 _2722_ (.A(_0568_),
    .B(_0569_),
    .X(_0571_));
 sky130_fd_sc_hd__a32o_1 _2723_ (.A1(_0546_),
    .A2(_0570_),
    .A3(_0571_),
    .B1(_0555_),
    .B2(\internalDataflow.addressLowBusModule.busInputs[18] ),
    .X(_0572_));
 sky130_fd_sc_hd__a21o_1 _2724_ (.A1(_0544_),
    .A2(_0567_),
    .B1(_0572_),
    .X(_0060_));
 sky130_fd_sc_hd__and3b_1 _2725_ (.A_N(_0221_),
    .B(_0559_),
    .C(_0562_),
    .X(_0573_));
 sky130_fd_sc_hd__a31o_1 _2726_ (.A1(_0221_),
    .A2(_0537_),
    .A3(_0561_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__xor2_1 _2727_ (.A(_0200_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__and2_1 _2728_ (.A(\internalDataflow.addressLowBusModule.busInputs[18] ),
    .B(_0535_),
    .X(_0576_));
 sky130_fd_sc_hd__and2_1 _2729_ (.A(_0568_),
    .B(_0569_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_1 _2730_ (.A(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .B(_0558_),
    .Y(_0578_));
 sky130_fd_sc_hd__and2_1 _2731_ (.A(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .B(_0535_),
    .X(_0579_));
 sky130_fd_sc_hd__nor2_1 _2732_ (.A(_0578_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__o21ai_1 _2733_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__o31a_1 _2734_ (.A1(_0576_),
    .A2(_0577_),
    .A3(_0580_),
    .B1(_0553_),
    .X(_0582_));
 sky130_fd_sc_hd__a22o_1 _2735_ (.A1(_0544_),
    .A2(_0575_),
    .B1(_0581_),
    .B2(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(_0583_),
    .A1(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .S(_0554_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _2737_ (.A(_0584_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _2738_ (.A(\internalDataflow.addressLowBusModule.busInputs[20] ),
    .B(_0535_),
    .X(_0585_));
 sky130_fd_sc_hd__nor2_1 _2739_ (.A(\internalDataflow.addressLowBusModule.busInputs[20] ),
    .B(_0535_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _2740_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _2741_ (.A(\internalDataflow.addressLowBusModule.busInputs[19] ),
    .B(_0534_),
    .X(_0588_));
 sky130_fd_sc_hd__a311o_1 _2742_ (.A1(_0568_),
    .A2(_0569_),
    .A3(_0588_),
    .B1(_0579_),
    .C1(_0576_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _2743_ (.A(_0587_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a211o_1 _2744_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0538_),
    .C1(_0544_),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _2745_ (.A(_0200_),
    .B(_0221_),
    .C(_0561_),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _2746_ (.A1(_0176_),
    .A2(_0592_),
    .B1(_0558_),
    .X(_0593_));
 sky130_fd_sc_hd__nor2_1 _2747_ (.A(_0177_),
    .B(_0592_),
    .Y(_0594_));
 sky130_fd_sc_hd__and4bb_1 _2748_ (.A_N(_0200_),
    .B_N(_0221_),
    .C(_0522_),
    .D(_0562_),
    .X(_0595_));
 sky130_fd_sc_hd__xnor2_1 _2749_ (.A(_0177_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__o22a_1 _2750_ (.A1(_0593_),
    .A2(_0594_),
    .B1(_0596_),
    .B2(_0537_),
    .X(_0597_));
 sky130_fd_sc_hd__o2bb2a_1 _2751_ (.A1_N(\internalDataflow.addressLowBusModule.busInputs[20] ),
    .A2_N(_0555_),
    .B1(_0597_),
    .B2(_0553_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ai_1 _2752_ (.A1(_0590_),
    .A2(_0591_),
    .B1(_0598_),
    .Y(_0062_));
 sky130_fd_sc_hd__or2_1 _2753_ (.A(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0535_),
    .X(_0599_));
 sky130_fd_sc_hd__nand2_1 _2754_ (.A(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0558_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _2755_ (.A(_0599_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__a21o_1 _2756_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0585_),
    .X(_0602_));
 sky130_fd_sc_hd__xnor2_1 _2757_ (.A(_0601_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _2758_ (.A(_0595_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_2 _2759_ (.A1(_0177_),
    .A2(_0604_),
    .B1(_0536_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _2760_ (.A(_0593_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__xor2_1 _2761_ (.A(_0153_),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__nor2_1 _2762_ (.A(_0553_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__a221o_1 _2763_ (.A1(net133),
    .A2(_0555_),
    .B1(_0603_),
    .B2(_0546_),
    .C1(_0608_),
    .X(_0063_));
 sky130_fd_sc_hd__a31o_1 _2764_ (.A1(_0153_),
    .A2(_0176_),
    .A3(_0592_),
    .B1(_0558_),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_1 _2765_ (.A(_0153_),
    .B(_0558_),
    .Y(_0610_));
 sky130_fd_sc_hd__and3_1 _2766_ (.A(_0605_),
    .B(_0609_),
    .C(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__xor2_1 _2767_ (.A(_0130_),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__and2_1 _2768_ (.A(\internalDataflow.addressLowBusModule.busInputs[22] ),
    .B(_0535_),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_1 _2769_ (.A(\internalDataflow.addressLowBusModule.busInputs[22] ),
    .B(_0536_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _2770_ (.A(_0613_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__and2_1 _2771_ (.A(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .B(_0535_),
    .X(_0616_));
 sky130_fd_sc_hd__a311o_1 _2772_ (.A1(_0587_),
    .A2(_0589_),
    .A3(_0599_),
    .B1(_0616_),
    .C1(_0585_),
    .X(_0617_));
 sky130_fd_sc_hd__a21boi_1 _2773_ (.A1(_0615_),
    .A2(_0617_),
    .B1_N(_0546_),
    .Y(_0618_));
 sky130_fd_sc_hd__o21a_1 _2774_ (.A1(_0615_),
    .A2(_0617_),
    .B1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__a221o_1 _2775_ (.A1(net120),
    .A2(_0555_),
    .B1(_0612_),
    .B2(_0544_),
    .C1(_0619_),
    .X(_0064_));
 sky130_fd_sc_hd__a41o_1 _2776_ (.A1(_0129_),
    .A2(_0153_),
    .A3(_0176_),
    .A4(_0592_),
    .B1(_0536_),
    .X(_0620_));
 sky130_fd_sc_hd__o21ai_1 _2777_ (.A1(_0130_),
    .A2(_0153_),
    .B1(_0536_),
    .Y(_0621_));
 sky130_fd_sc_hd__and3_1 _2778_ (.A(_0605_),
    .B(_0620_),
    .C(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__xor2_1 _2779_ (.A(_0312_),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _2780_ (.A(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .B(_0535_),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_1 _2781_ (.A(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .B(_0558_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _2782_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a21oi_1 _2783_ (.A1(_0615_),
    .A2(_0617_),
    .B1(_0613_),
    .Y(_0627_));
 sky130_fd_sc_hd__or2_1 _2784_ (.A(_0626_),
    .B(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__a21oi_1 _2785_ (.A1(_0626_),
    .A2(_0627_),
    .B1(_0544_),
    .Y(_0629_));
 sky130_fd_sc_hd__a22o_1 _2786_ (.A1(_0544_),
    .A2(_0623_),
    .B1(_0628_),
    .B2(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(_0630_),
    .A1(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .S(_0554_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _2788_ (.A(_0631_),
    .X(_0065_));
 sky130_fd_sc_hd__nand2_4 _2789_ (.A(_1383_),
    .B(_1386_),
    .Y(_0632_));
 sky130_fd_sc_hd__nor2_2 _2790_ (.A(_1326_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__and3_2 _2791_ (.A(_1383_),
    .B(_1386_),
    .C(_1329_),
    .X(_0634_));
 sky130_fd_sc_hd__o2111a_1 _2792_ (.A1(_1430_),
    .A2(_0245_),
    .B1(_0246_),
    .C1(_0247_),
    .D1(_0632_),
    .X(_0635_));
 sky130_fd_sc_hd__a221o_2 _2793_ (.A1(_0231_),
    .A2(_0633_),
    .B1(_0634_),
    .B2(_0234_),
    .C1(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__o21a_1 _2794_ (.A1(_1007_),
    .A2(_1400_),
    .B1(_1168_),
    .X(_0637_));
 sky130_fd_sc_hd__inv_2 _2795_ (.A(_0820_),
    .Y(_0638_));
 sky130_fd_sc_hd__o211a_1 _2796_ (.A1(_1007_),
    .A2(_0491_),
    .B1(_1084_),
    .C1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__a221o_1 _2797_ (.A1(\demux.state_machine.timeState[3] ),
    .A2(_1079_),
    .B1(_0494_),
    .B2(_1102_),
    .C1(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__or3_1 _2798_ (.A(_0489_),
    .B(_0637_),
    .C(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _2799_ (.A(_1384_),
    .B(_1487_),
    .C(_0488_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__a221o_1 _2800_ (.A1(_0985_),
    .A2(_1283_),
    .B1(_1441_),
    .B2(_0987_),
    .C1(_0500_),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _2801_ (.A(_0999_),
    .B(_0642_),
    .C(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_8 _2802_ (.A(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(net102),
    .A1(_0636_),
    .S(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _2804_ (.A(_0646_),
    .X(_0066_));
 sky130_fd_sc_hd__inv_2 _2805_ (.A(net44),
    .Y(_0647_));
 sky130_fd_sc_hd__and3_1 _2806_ (.A(_1431_),
    .B(_0272_),
    .C(_0632_),
    .X(_0648_));
 sky130_fd_sc_hd__a221o_2 _2807_ (.A1(_0647_),
    .A2(_0633_),
    .B1(_0634_),
    .B2(_0265_),
    .C1(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(net17),
    .A1(_0649_),
    .S(_0645_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _2809_ (.A(_0650_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _2810_ (.A(_0207_),
    .B(_0634_),
    .X(_0651_));
 sky130_fd_sc_hd__a221o_2 _2811_ (.A1(_0213_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0212_),
    .C1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(net108),
    .A1(_0652_),
    .S(_0645_),
    .X(_0653_));
 sky130_fd_sc_hd__clkbuf_1 _2813_ (.A(_0653_),
    .X(_0068_));
 sky130_fd_sc_hd__or2_1 _2814_ (.A(_1326_),
    .B(_0632_),
    .X(_0654_));
 sky130_fd_sc_hd__a2bb2o_1 _2815_ (.A1_N(_0191_),
    .A2_N(_0654_),
    .B1(_0632_),
    .B2(_0192_),
    .X(_0655_));
 sky130_fd_sc_hd__a21o_1 _2816_ (.A1(_0185_),
    .A2(_0634_),
    .B1(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(net91),
    .A1(_0656_),
    .S(_0645_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_1 _2818_ (.A(_0657_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _2819_ (.A1(_0163_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0162_),
    .X(_0658_));
 sky130_fd_sc_hd__a21o_2 _2820_ (.A1(_0169_),
    .A2(_0634_),
    .B1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(net127),
    .A1(_0659_),
    .S(_0645_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _2822_ (.A(_0660_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _2823_ (.A(_0145_),
    .B(_0634_),
    .X(_0661_));
 sky130_fd_sc_hd__a221o_2 _2824_ (.A1(_0141_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0140_),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _2825_ (.A0(net115),
    .A1(_0662_),
    .S(_0645_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _2826_ (.A(_0663_),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _2827_ (.A(_1481_),
    .B(_0654_),
    .Y(_0664_));
 sky130_fd_sc_hd__a221o_2 _2828_ (.A1(_1432_),
    .A2(_0632_),
    .B1(_0634_),
    .B2(_1321_),
    .C1(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(net124),
    .A1(_0665_),
    .S(_0645_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_1 _2830_ (.A(_0666_),
    .X(_0072_));
 sky130_fd_sc_hd__inv_2 _2831_ (.A(_0299_),
    .Y(_0667_));
 sky130_fd_sc_hd__nor2_1 _2832_ (.A(_0296_),
    .B(_0654_),
    .Y(_0668_));
 sky130_fd_sc_hd__a221o_2 _2833_ (.A1(_0667_),
    .A2(_0632_),
    .B1(_0634_),
    .B2(_0304_),
    .C1(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _2834_ (.A0(net121),
    .A1(_0669_),
    .S(_0645_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _2835_ (.A(_0670_),
    .X(_0073_));
 sky130_fd_sc_hd__or3_1 _2836_ (.A(\instructionLoader.interruptInjector.processStatusRegIFlag ),
    .B(\demux.setInterruptFlag ),
    .C(_0961_),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_1 _2837_ (.A1(\instructionLoader.interruptInjector.resetDetected ),
    .A2(_0999_),
    .B1(_0671_),
    .B2(\demux.reset ),
    .X(_0074_));
 sky130_fd_sc_hd__or3_1 _2838_ (.A(_0837_),
    .B(_1152_),
    .C(_1190_),
    .X(_0672_));
 sky130_fd_sc_hd__a22o_1 _2839_ (.A1(_1002_),
    .A2(_0867_),
    .B1(_0672_),
    .B2(_1008_),
    .X(_0673_));
 sky130_fd_sc_hd__and2_1 _2840_ (.A(_0332_),
    .B(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_4 _2841_ (.A(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(_0224_),
    .A1(_0249_),
    .S(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__inv_2 _2843_ (.A(_0676_),
    .Y(_0075_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(net128),
    .A1(_0274_),
    .S(_0675_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_0677_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(net105),
    .A1(_0215_),
    .S(_0675_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_0678_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(net110),
    .A1(_0194_),
    .S(_0675_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _2849_ (.A(_0679_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(net107),
    .A1(_0170_),
    .S(_0675_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _2851_ (.A(_0680_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(net103),
    .A1(_0146_),
    .S(_0675_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_1 _2853_ (.A(_0681_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(net100),
    .A1(_1434_),
    .S(_0675_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _2855_ (.A(_0682_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\internalDataflow.stackBusModule.busInputs[47] ),
    .A1(_0305_),
    .S(_0675_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _2857_ (.A(_0683_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _2858_ (.A(\internalDataflow.addressLowBusModule.busInputs[32] ),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _2859_ (.A(_1489_),
    .Y(_0685_));
 sky130_fd_sc_hd__a211o_1 _2860_ (.A1(_1008_),
    .A2(_1204_),
    .B1(_0685_),
    .C1(_0916_),
    .X(_0686_));
 sky130_fd_sc_hd__o31a_4 _2861_ (.A1(_0924_),
    .A2(_1362_),
    .A3(_0686_),
    .B1(_0332_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(_0684_),
    .A1(_0249_),
    .S(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _2863_ (.A(_0688_),
    .Y(_0083_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(\internalDataflow.addressLowBusModule.busInputs[33] ),
    .A1(_0274_),
    .S(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _2865_ (.A(_0689_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(\internalDataflow.addressLowBusModule.busInputs[34] ),
    .A1(_0215_),
    .S(_0687_),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _2867_ (.A(_0690_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\internalDataflow.addressLowBusModule.busInputs[35] ),
    .A1(_0194_),
    .S(_0687_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_0691_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\internalDataflow.addressLowBusModule.busInputs[36] ),
    .A1(_0170_),
    .S(_0687_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _2871_ (.A(_0692_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\internalDataflow.addressLowBusModule.busInputs[37] ),
    .A1(_0146_),
    .S(_0687_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _2873_ (.A(_0693_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\internalDataflow.addressLowBusModule.busInputs[38] ),
    .A1(_1434_),
    .S(_0687_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_0694_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\internalDataflow.addressLowBusModule.busInputs[39] ),
    .A1(_0305_),
    .S(_0687_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_0695_),
    .X(_0090_));
 sky130_fd_sc_hd__xor2_1 _2878_ (.A(\internalDataflow.addressHighBusModule.busInputs[16] ),
    .B(_0536_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _2879_ (.A(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .B(_0536_),
    .X(_0697_));
 sky130_fd_sc_hd__a311o_1 _2880_ (.A1(_0615_),
    .A2(_0617_),
    .A3(_0624_),
    .B1(_0697_),
    .C1(_0613_),
    .X(_0698_));
 sky130_fd_sc_hd__or2_1 _2881_ (.A(_0696_),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_1 _2882_ (.A(_0696_),
    .B(_0698_),
    .Y(_0700_));
 sky130_fd_sc_hd__xnor2_1 _2883_ (.A(_0312_),
    .B(_0537_),
    .Y(_0701_));
 sky130_fd_sc_hd__and4_1 _2884_ (.A(_0605_),
    .B(_0620_),
    .C(_0621_),
    .D(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__nand2_1 _2885_ (.A(_0636_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__or2_1 _2886_ (.A(_0636_),
    .B(_0702_),
    .X(_0704_));
 sky130_fd_sc_hd__a32o_1 _2887_ (.A1(_0544_),
    .A2(_0703_),
    .A3(_0704_),
    .B1(_0555_),
    .B2(\internalDataflow.addressHighBusModule.busInputs[16] ),
    .X(_0705_));
 sky130_fd_sc_hd__a31o_1 _2888_ (.A1(_0546_),
    .A2(_0699_),
    .A3(_0700_),
    .B1(_0705_),
    .X(_0091_));
 sky130_fd_sc_hd__xnor2_1 _2889_ (.A(_0312_),
    .B(_0636_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _2890_ (.A(_0702_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__xnor2_1 _2891_ (.A(_0649_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _2892_ (.A(\internalDataflow.addressHighBusModule.busInputs[16] ),
    .B(_0536_),
    .Y(_0709_));
 sky130_fd_sc_hd__nor2_1 _2893_ (.A(\internalDataflow.addressHighBusModule.busInputs[17] ),
    .B(_0536_),
    .Y(_0710_));
 sky130_fd_sc_hd__and2_1 _2894_ (.A(\internalDataflow.addressHighBusModule.busInputs[17] ),
    .B(_0556_),
    .X(_0711_));
 sky130_fd_sc_hd__nor2_1 _2895_ (.A(_0710_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__a21oi_1 _2896_ (.A1(_0709_),
    .A2(_0700_),
    .B1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__and3_1 _2897_ (.A(_0709_),
    .B(_0700_),
    .C(_0712_),
    .X(_0714_));
 sky130_fd_sc_hd__or2_1 _2898_ (.A(_0713_),
    .B(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(_0708_),
    .A1(_0715_),
    .S(_0553_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(_0716_),
    .A1(\internalDataflow.addressHighBusModule.busInputs[17] ),
    .S(_0554_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _2901_ (.A(_0717_),
    .X(_0092_));
 sky130_fd_sc_hd__a21oi_1 _2902_ (.A1(_0709_),
    .A2(_0700_),
    .B1(_0710_),
    .Y(_0718_));
 sky130_fd_sc_hd__xor2_1 _2903_ (.A(\internalDataflow.addressHighBusModule.busInputs[18] ),
    .B(_0556_),
    .X(_0719_));
 sky130_fd_sc_hd__o21ai_1 _2904_ (.A1(_0711_),
    .A2(_0718_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__o31a_1 _2905_ (.A1(_0711_),
    .A2(_0719_),
    .A3(_0718_),
    .B1(_0546_),
    .X(_0721_));
 sky130_fd_sc_hd__and2_1 _2906_ (.A(_0556_),
    .B(_0649_),
    .X(_0722_));
 sky130_fd_sc_hd__nor2_1 _2907_ (.A(_0556_),
    .B(_0649_),
    .Y(_0723_));
 sky130_fd_sc_hd__or3_1 _2908_ (.A(_0707_),
    .B(_0722_),
    .C(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__xor2_1 _2909_ (.A(_0652_),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nor2_1 _2910_ (.A(_0553_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__a221o_1 _2911_ (.A1(net130),
    .A2(_0555_),
    .B1(_0720_),
    .B2(_0721_),
    .C1(_0726_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _2912_ (.A(_0537_),
    .B(_0652_),
    .Y(_0727_));
 sky130_fd_sc_hd__or2_1 _2913_ (.A(_0537_),
    .B(_0652_),
    .X(_0728_));
 sky130_fd_sc_hd__a21oi_1 _2914_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0724_),
    .Y(_0729_));
 sky130_fd_sc_hd__xor2_1 _2915_ (.A(_0656_),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nor2_1 _2916_ (.A(\internalDataflow.addressHighBusModule.busInputs[19] ),
    .B(_0556_),
    .Y(_0731_));
 sky130_fd_sc_hd__and2_1 _2917_ (.A(\internalDataflow.addressHighBusModule.busInputs[19] ),
    .B(_0556_),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _2918_ (.A(_0731_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__a21boi_2 _2919_ (.A1(\internalDataflow.addressHighBusModule.busInputs[18] ),
    .A2(_0556_),
    .B1_N(_0720_),
    .Y(_0734_));
 sky130_fd_sc_hd__xnor2_1 _2920_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(_0730_),
    .A1(_0735_),
    .S(_0553_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_0736_),
    .A1(\internalDataflow.addressHighBusModule.busInputs[19] ),
    .S(_0554_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_0737_),
    .X(_0094_));
 sky130_fd_sc_hd__nand2_1 _2924_ (.A(\internalDataflow.addressHighBusModule.busInputs[20] ),
    .B(_0556_),
    .Y(_0738_));
 sky130_fd_sc_hd__or2_1 _2925_ (.A(\internalDataflow.addressHighBusModule.busInputs[20] ),
    .B(_0556_),
    .X(_0739_));
 sky130_fd_sc_hd__and2_1 _2926_ (.A(_0738_),
    .B(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__o21bai_2 _2927_ (.A1(_0731_),
    .A2(_0734_),
    .B1_N(_0732_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _2928_ (.A(_0740_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__o21a_1 _2929_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0546_),
    .X(_0743_));
 sky130_fd_sc_hd__nand2_1 _2930_ (.A(_0557_),
    .B(_0656_),
    .Y(_0744_));
 sky130_fd_sc_hd__or2_1 _2931_ (.A(_0557_),
    .B(_0656_),
    .X(_0745_));
 sky130_fd_sc_hd__and3_1 _2932_ (.A(_0729_),
    .B(_0744_),
    .C(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__o21ai_1 _2933_ (.A1(_0659_),
    .A2(_0746_),
    .B1(_0544_),
    .Y(_0747_));
 sky130_fd_sc_hd__a21oi_1 _2934_ (.A1(_0659_),
    .A2(_0746_),
    .B1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__a221o_1 _2935_ (.A1(net132),
    .A2(_0555_),
    .B1(_0742_),
    .B2(_0743_),
    .C1(_0748_),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _2936_ (.A(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .B(_0557_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _2937_ (.A(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .B(_0558_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(_0749_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__a21bo_1 _2939_ (.A1(_0740_),
    .A2(_0741_),
    .B1_N(_0738_),
    .X(_0752_));
 sky130_fd_sc_hd__xnor2_1 _2940_ (.A(_0751_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__xnor2_1 _2941_ (.A(_0537_),
    .B(_0659_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _2942_ (.A(_0746_),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _2943_ (.A(_0662_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__or2_1 _2944_ (.A(_0662_),
    .B(_0755_),
    .X(_0757_));
 sky130_fd_sc_hd__a21oi_1 _2945_ (.A1(_0756_),
    .A2(_0757_),
    .B1(_0553_),
    .Y(_0758_));
 sky130_fd_sc_hd__a221o_1 _2946_ (.A1(net125),
    .A2(_0555_),
    .B1(_0753_),
    .B2(_0546_),
    .C1(_0758_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _2947_ (.A(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .B(_0557_),
    .Y(_0759_));
 sky130_fd_sc_hd__or2_1 _2948_ (.A(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .B(_0558_),
    .X(_0760_));
 sky130_fd_sc_hd__and2_1 _2949_ (.A(_0759_),
    .B(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__and2_1 _2950_ (.A(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .B(_0557_),
    .X(_0762_));
 sky130_fd_sc_hd__a21oi_1 _2951_ (.A1(_0749_),
    .A2(_0752_),
    .B1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__xnor2_1 _2952_ (.A(_0761_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__xnor2_1 _2953_ (.A(_0557_),
    .B(_0662_),
    .Y(_0765_));
 sky130_fd_sc_hd__nor2_1 _2954_ (.A(_0755_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__o21ai_1 _2955_ (.A1(_0665_),
    .A2(_0766_),
    .B1(_0544_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21oi_1 _2956_ (.A1(_0665_),
    .A2(_0766_),
    .B1(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__a221o_1 _2957_ (.A1(net119),
    .A2(_0555_),
    .B1(_0764_),
    .B2(_0546_),
    .C1(_0768_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _2958_ (.A(_0557_),
    .B(_0665_),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _2959_ (.A(_0558_),
    .B(_0665_),
    .Y(_0770_));
 sky130_fd_sc_hd__or4_1 _2960_ (.A(_0755_),
    .B(_0765_),
    .C(_0769_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__xnor2_1 _2961_ (.A(_0669_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__nor2_1 _2962_ (.A(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .B(_0557_),
    .Y(_0773_));
 sky130_fd_sc_hd__o21a_1 _2963_ (.A1(_0773_),
    .A2(_0763_),
    .B1(_0759_),
    .X(_0774_));
 sky130_fd_sc_hd__xnor2_1 _2964_ (.A(\internalDataflow.addressHighBusModule.busInputs[23] ),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__xnor2_1 _2965_ (.A(_0537_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_0772_),
    .A1(_0776_),
    .S(_0553_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_0777_),
    .A1(\internalDataflow.addressHighBusModule.busInputs[23] ),
    .S(_0554_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_0778_),
    .X(_0098_));
 sky130_fd_sc_hd__or2b_1 _2969_ (.A(_1297_),
    .B_N(_1254_),
    .X(_0779_));
 sky130_fd_sc_hd__or3_1 _2970_ (.A(_1384_),
    .B(_1260_),
    .C(_1330_),
    .X(_0780_));
 sky130_fd_sc_hd__a221o_1 _2971_ (.A1(_1002_),
    .A2(_0929_),
    .B1(_1282_),
    .B2(_1102_),
    .C1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__and3_1 _2972_ (.A(_0999_),
    .B(_0779_),
    .C(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_8 _2973_ (.A(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(net126),
    .A1(_0236_),
    .S(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_1 _2975_ (.A(_0784_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(net33),
    .A1(_0276_),
    .S(_0783_),
    .X(_0785_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_0785_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(net34),
    .A1(_0217_),
    .S(_0783_),
    .X(_0786_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_0786_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(net88),
    .A1(_0196_),
    .S(_0783_),
    .X(_0787_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_0787_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(net116),
    .A1(_0172_),
    .S(_0783_),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_0788_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(net117),
    .A1(_0149_),
    .S(_0783_),
    .X(_0789_));
 sky130_fd_sc_hd__clkbuf_1 _2985_ (.A(_0789_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(net38),
    .A1(_1482_),
    .S(_0783_),
    .X(_0790_));
 sky130_fd_sc_hd__clkbuf_1 _2987_ (.A(_0790_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(net87),
    .A1(_0308_),
    .S(_0783_),
    .X(_0791_));
 sky130_fd_sc_hd__clkbuf_1 _2989_ (.A(_0791_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_1 _2990_ (.A(_0981_),
    .B(_0340_),
    .X(_0792_));
 sky130_fd_sc_hd__or4b_1 _2991_ (.A(\instructionLoader.interruptInjector.processStatusRegIFlag ),
    .B(\demux.setInterruptFlag ),
    .C(\instructionLoader.interruptInjector.irqGenerated ),
    .D_N(\instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ),
    .X(_0793_));
 sky130_fd_sc_hd__a21bo_1 _2992_ (.A1(net90),
    .A2(_0792_),
    .B1_N(_0793_),
    .X(_0107_));
 sky130_fd_sc_hd__or3b_1 _2993_ (.A(\demux.nmi ),
    .B(\instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ),
    .C_N(\instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ),
    .X(_0794_));
 sky130_fd_sc_hd__a21bo_1 _2994_ (.A1(\demux.nmi ),
    .A2(_0792_),
    .B1_N(_0794_),
    .X(_0108_));
 sky130_fd_sc_hd__a21oi_1 _2995_ (.A1(_0999_),
    .A2(_1022_),
    .B1(net92),
    .Y(_0795_));
 sky130_fd_sc_hd__nor2_1 _2996_ (.A(_0341_),
    .B(_0795_),
    .Y(_0109_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(net14),
    .A1(net89),
    .S(_0981_),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_0796_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _2999_ (.A(\demux.nmi ),
    .B(_0671_),
    .X(_0797_));
 sky130_fd_sc_hd__a22o_1 _3000_ (.A1(\demux.nmi ),
    .A2(_0341_),
    .B1(_0797_),
    .B2(net77),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _3001_ (.A(\instructionLoader.interruptInjector.resetDetected ),
    .B(_0981_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_0798_),
    .X(_0112_));
 sky130_fd_sc_hd__a211o_1 _3003_ (.A1(_0529_),
    .A2(_1437_),
    .B1(_0961_),
    .C1(_1281_),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(_0385_),
    .A1(net118),
    .S(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_1 _3005_ (.A(_0800_),
    .X(_0113_));
 sky130_fd_sc_hd__nand2_1 _3006_ (.A(_0905_),
    .B(_0323_),
    .Y(_0801_));
 sky130_fd_sc_hd__and4_1 _3007_ (.A(_0968_),
    .B(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .C(_0905_),
    .D(_0323_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _3008_ (.A1(net94),
    .A2(_0801_),
    .B1(_0802_),
    .B2(_0385_),
    .X(_0114_));
 sky130_fd_sc_hd__a21o_1 _3009_ (.A1(_0947_),
    .A2(_0996_),
    .B1(_0961_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(_0979_),
    .A1(_0803_),
    .S(\demux.isAddressing ),
    .X(_0804_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_0804_),
    .X(_0115_));
 sky130_fd_sc_hd__or3_1 _3012_ (.A(_0968_),
    .B(\internalDataflow.addressLowBusModule.busInputs[23] ),
    .C(_0801_),
    .X(_0805_));
 sky130_fd_sc_hd__a2bb2o_1 _3013_ (.A1_N(_0385_),
    .A2_N(_0805_),
    .B1(_0801_),
    .B2(net95),
    .X(_0116_));
 sky130_fd_sc_hd__o31a_1 _3014_ (.A1(_0915_),
    .A2(_1249_),
    .A3(_1358_),
    .B1(_1002_),
    .X(_0806_));
 sky130_fd_sc_hd__a21bo_1 _3015_ (.A1(_1002_),
    .A2(_0847_),
    .B1_N(_0328_),
    .X(_0807_));
 sky130_fd_sc_hd__o31a_1 _3016_ (.A1(_0806_),
    .A2(_0347_),
    .A3(_0807_),
    .B1(_0332_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _3017_ (.A0(\demux.PSR_N ),
    .A1(_0308_),
    .S(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_1 _3018_ (.A(_0809_),
    .X(_0117_));
 sky130_fd_sc_hd__dfstp_1 _3019_ (.CLK(clknet_4_7_0_clk),
    .D(_0000_),
    .SET_B(net68),
    .Q(\demux.state_machine.currentAddress[0] ));
 sky130_fd_sc_hd__dfrtp_2 _3020_ (.CLK(clknet_4_6_0_clk),
    .D(_0004_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3021_ (.CLK(clknet_4_7_0_clk),
    .D(_0005_),
    .RESET_B(net68),
    .Q(\demux.state_machine.currentAddress[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3022_ (.CLK(clknet_4_7_0_clk),
    .D(_0006_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3023_ (.CLK(clknet_4_6_0_clk),
    .D(_0007_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3024_ (.CLK(clknet_4_7_0_clk),
    .D(_0008_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3025_ (.CLK(clknet_4_7_0_clk),
    .D(_0009_),
    .RESET_B(net68),
    .Q(\demux.state_machine.currentAddress[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3026_ (.CLK(clknet_4_7_0_clk),
    .D(_0010_),
    .RESET_B(net68),
    .Q(\demux.state_machine.currentAddress[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3027_ (.CLK(clknet_4_7_0_clk),
    .D(_0011_),
    .RESET_B(net68),
    .Q(\demux.state_machine.currentAddress[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3028_ (.CLK(clknet_4_7_0_clk),
    .D(_0012_),
    .RESET_B(net68),
    .Q(\demux.state_machine.currentAddress[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3029_ (.CLK(clknet_4_7_0_clk),
    .D(_0001_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3030_ (.CLK(clknet_4_6_0_clk),
    .D(_0002_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3031_ (.CLK(clknet_4_7_0_clk),
    .D(_0003_),
    .RESET_B(net67),
    .Q(\demux.state_machine.currentAddress[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3032_ (.CLK(clknet_4_3_0_clk),
    .D(_0026_),
    .RESET_B(net60),
    .Q(\internalDataflow.stackBusModule.busInputs[32] ));
 sky130_fd_sc_hd__dfrtp_1 _3033_ (.CLK(clknet_4_2_0_clk),
    .D(_0027_),
    .RESET_B(net58),
    .Q(\internalDataflow.stackBusModule.busInputs[33] ));
 sky130_fd_sc_hd__dfrtp_1 _3034_ (.CLK(clknet_4_8_0_clk),
    .D(_0028_),
    .RESET_B(net62),
    .Q(\internalDataflow.stackBusModule.busInputs[34] ));
 sky130_fd_sc_hd__dfrtp_1 _3035_ (.CLK(clknet_4_2_0_clk),
    .D(_0029_),
    .RESET_B(net58),
    .Q(\internalDataflow.stackBusModule.busInputs[35] ));
 sky130_fd_sc_hd__dfrtp_1 _3036_ (.CLK(clknet_4_2_0_clk),
    .D(_0030_),
    .RESET_B(net58),
    .Q(\internalDataflow.stackBusModule.busInputs[36] ));
 sky130_fd_sc_hd__dfrtp_1 _3037_ (.CLK(clknet_4_3_0_clk),
    .D(_0031_),
    .RESET_B(net59),
    .Q(\internalDataflow.stackBusModule.busInputs[37] ));
 sky130_fd_sc_hd__dfrtp_1 _3038_ (.CLK(clknet_4_3_0_clk),
    .D(_0032_),
    .RESET_B(net58),
    .Q(\internalDataflow.stackBusModule.busInputs[38] ));
 sky130_fd_sc_hd__dfrtp_1 _3039_ (.CLK(clknet_4_8_0_clk),
    .D(_0033_),
    .RESET_B(net62),
    .Q(\internalDataflow.stackBusModule.busInputs[39] ));
 sky130_fd_sc_hd__dfrtp_1 _3040_ (.CLK(clknet_4_4_0_clk),
    .D(\pulse_slower.nextEnableState[0] ),
    .RESET_B(net60),
    .Q(\pulse_slower.currentEnableState[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3041_ (.CLK(clknet_4_4_0_clk),
    .D(\pulse_slower.nextEnableState[1] ),
    .RESET_B(net60),
    .Q(\pulse_slower.currentEnableState[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3042_ (.CLK(clknet_4_1_0_clk),
    .D(_0034_),
    .RESET_B(net60),
    .Q(\internalDataflow.addressLowBusModule.busInputs[24] ));
 sky130_fd_sc_hd__dfrtp_1 _3043_ (.CLK(clknet_4_0_0_clk),
    .D(_0035_),
    .RESET_B(net57),
    .Q(\internalDataflow.addressLowBusModule.busInputs[25] ));
 sky130_fd_sc_hd__dfrtp_1 _3044_ (.CLK(clknet_4_0_0_clk),
    .D(_0036_),
    .RESET_B(net57),
    .Q(\internalDataflow.addressLowBusModule.busInputs[26] ));
 sky130_fd_sc_hd__dfrtp_1 _3045_ (.CLK(clknet_4_0_0_clk),
    .D(_0037_),
    .RESET_B(net57),
    .Q(\internalDataflow.addressLowBusModule.busInputs[27] ));
 sky130_fd_sc_hd__dfrtp_1 _3046_ (.CLK(clknet_4_1_0_clk),
    .D(_0038_),
    .RESET_B(net57),
    .Q(\internalDataflow.addressLowBusModule.busInputs[28] ));
 sky130_fd_sc_hd__dfrtp_1 _3047_ (.CLK(clknet_4_1_0_clk),
    .D(_0039_),
    .RESET_B(net60),
    .Q(\internalDataflow.addressLowBusModule.busInputs[29] ));
 sky130_fd_sc_hd__dfrtp_2 _3048_ (.CLK(clknet_4_1_0_clk),
    .D(_0040_),
    .RESET_B(net60),
    .Q(\internalDataflow.addressLowBusModule.busInputs[30] ));
 sky130_fd_sc_hd__dfrtp_1 _3049_ (.CLK(clknet_4_0_0_clk),
    .D(_0041_),
    .RESET_B(net57),
    .Q(\internalDataflow.addressLowBusModule.busInputs[31] ));
 sky130_fd_sc_hd__dfrtp_1 _3050_ (.CLK(clknet_4_4_0_clk),
    .D(_0042_),
    .RESET_B(net60),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _3051_ (.CLK(clknet_4_0_0_clk),
    .D(_0043_),
    .RESET_B(net57),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _3052_ (.CLK(clknet_4_1_0_clk),
    .D(_0044_),
    .RESET_B(net61),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _3053_ (.CLK(clknet_4_8_0_clk),
    .D(_0045_),
    .RESET_B(net62),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _3054_ (.CLK(clknet_4_14_0_clk),
    .D(_0046_),
    .RESET_B(net70),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _3055_ (.CLK(clknet_4_4_0_clk),
    .D(_0047_),
    .RESET_B(net69),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _3056_ (.CLK(clknet_4_0_0_clk),
    .D(_0048_),
    .RESET_B(net57),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _3057_ (.CLK(clknet_4_13_0_clk),
    .D(_0049_),
    .RESET_B(net70),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _3058_ (.CLK(clknet_4_3_0_clk),
    .D(_0050_),
    .RESET_B(net63),
    .Q(\internalDataflow.accRegToDB[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3059_ (.CLK(clknet_4_8_0_clk),
    .D(_0051_),
    .RESET_B(net62),
    .Q(\internalDataflow.accRegToDB[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3060_ (.CLK(clknet_4_8_0_clk),
    .D(_0052_),
    .RESET_B(net62),
    .Q(\internalDataflow.accRegToDB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3061_ (.CLK(clknet_4_8_0_clk),
    .D(_0053_),
    .RESET_B(net62),
    .Q(\internalDataflow.accRegToDB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3062_ (.CLK(clknet_4_2_0_clk),
    .D(_0054_),
    .RESET_B(net62),
    .Q(\internalDataflow.accRegToDB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3063_ (.CLK(clknet_4_9_0_clk),
    .D(_0055_),
    .RESET_B(net63),
    .Q(\internalDataflow.accRegToDB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3064_ (.CLK(clknet_4_8_0_clk),
    .D(_0056_),
    .RESET_B(net63),
    .Q(\internalDataflow.accRegToDB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3065_ (.CLK(clknet_4_8_0_clk),
    .D(_0057_),
    .RESET_B(net62),
    .Q(\internalDataflow.accRegToDB[7] ));
 sky130_fd_sc_hd__dfrtp_2 _3066_ (.CLK(clknet_4_9_0_clk),
    .D(_0058_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[16] ));
 sky130_fd_sc_hd__dfrtp_4 _3067_ (.CLK(clknet_4_13_0_clk),
    .D(_0059_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3068_ (.CLK(clknet_4_9_0_clk),
    .D(_0060_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[18] ));
 sky130_fd_sc_hd__dfrtp_4 _3069_ (.CLK(clknet_4_9_0_clk),
    .D(_0061_),
    .RESET_B(net63),
    .Q(\internalDataflow.addressLowBusModule.busInputs[19] ));
 sky130_fd_sc_hd__dfrtp_2 _3070_ (.CLK(clknet_4_11_0_clk),
    .D(_0062_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[20] ));
 sky130_fd_sc_hd__dfrtp_4 _3071_ (.CLK(clknet_4_11_0_clk),
    .D(_0063_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3072_ (.CLK(clknet_4_12_0_clk),
    .D(_0064_),
    .RESET_B(net65),
    .Q(\internalDataflow.addressLowBusModule.busInputs[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3073_ (.CLK(clknet_4_13_0_clk),
    .D(_0065_),
    .RESET_B(net70),
    .Q(\internalDataflow.addressLowBusModule.busInputs[23] ));
 sky130_fd_sc_hd__dfrtp_1 _3074_ (.CLK(clknet_4_10_0_clk),
    .D(_0066_),
    .RESET_B(net64),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_2 _3075_ (.CLK(clknet_4_13_0_clk),
    .D(_0067_),
    .RESET_B(net70),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _3076_ (.CLK(clknet_4_2_0_clk),
    .D(_0068_),
    .RESET_B(net58),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _3077_ (.CLK(clknet_4_10_0_clk),
    .D(_0069_),
    .RESET_B(net64),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _3078_ (.CLK(clknet_4_5_0_clk),
    .D(_0070_),
    .RESET_B(net69),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _3079_ (.CLK(clknet_4_10_0_clk),
    .D(_0071_),
    .RESET_B(net64),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _3080_ (.CLK(clknet_4_10_0_clk),
    .D(_0072_),
    .RESET_B(net64),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _3081_ (.CLK(clknet_4_14_0_clk),
    .D(_0073_),
    .RESET_B(net71),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_4 _3082_ (.CLK(clknet_4_13_0_clk),
    .D(_0074_),
    .RESET_B(net70),
    .Q(\demux.reset ));
 sky130_fd_sc_hd__dfrtp_1 _3083_ (.CLK(clknet_4_3_0_clk),
    .D(_0075_),
    .RESET_B(net59),
    .Q(\internalDataflow.stackBusModule.busInputs[40] ));
 sky130_fd_sc_hd__dfrtp_1 _3084_ (.CLK(clknet_4_2_0_clk),
    .D(_0076_),
    .RESET_B(net59),
    .Q(\internalDataflow.stackBusModule.busInputs[41] ));
 sky130_fd_sc_hd__dfrtp_1 _3085_ (.CLK(clknet_4_8_0_clk),
    .D(_0077_),
    .RESET_B(net62),
    .Q(\internalDataflow.stackBusModule.busInputs[42] ));
 sky130_fd_sc_hd__dfrtp_1 _3086_ (.CLK(clknet_4_8_0_clk),
    .D(_0078_),
    .RESET_B(net63),
    .Q(\internalDataflow.stackBusModule.busInputs[43] ));
 sky130_fd_sc_hd__dfrtp_1 _3087_ (.CLK(clknet_4_2_0_clk),
    .D(_0079_),
    .RESET_B(net59),
    .Q(\internalDataflow.stackBusModule.busInputs[44] ));
 sky130_fd_sc_hd__dfrtp_1 _3088_ (.CLK(clknet_4_9_0_clk),
    .D(_0080_),
    .RESET_B(net63),
    .Q(\internalDataflow.stackBusModule.busInputs[45] ));
 sky130_fd_sc_hd__dfrtp_1 _3089_ (.CLK(clknet_4_3_0_clk),
    .D(_0081_),
    .RESET_B(net59),
    .Q(\internalDataflow.stackBusModule.busInputs[46] ));
 sky130_fd_sc_hd__dfrtp_1 _3090_ (.CLK(clknet_4_8_0_clk),
    .D(_0082_),
    .RESET_B(net62),
    .Q(\internalDataflow.stackBusModule.busInputs[47] ));
 sky130_fd_sc_hd__dfrtp_1 _3091_ (.CLK(clknet_4_3_0_clk),
    .D(_0083_),
    .RESET_B(net61),
    .Q(\internalDataflow.addressLowBusModule.busInputs[32] ));
 sky130_fd_sc_hd__dfrtp_1 _3092_ (.CLK(clknet_4_2_0_clk),
    .D(_0084_),
    .RESET_B(net58),
    .Q(\internalDataflow.addressLowBusModule.busInputs[33] ));
 sky130_fd_sc_hd__dfrtp_1 _3093_ (.CLK(clknet_4_2_0_clk),
    .D(_0085_),
    .RESET_B(net58),
    .Q(\internalDataflow.addressLowBusModule.busInputs[34] ));
 sky130_fd_sc_hd__dfrtp_1 _3094_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .RESET_B(net58),
    .Q(\internalDataflow.addressLowBusModule.busInputs[35] ));
 sky130_fd_sc_hd__dfrtp_1 _3095_ (.CLK(clknet_4_2_0_clk),
    .D(_0087_),
    .RESET_B(net58),
    .Q(\internalDataflow.addressLowBusModule.busInputs[36] ));
 sky130_fd_sc_hd__dfrtp_1 _3096_ (.CLK(clknet_4_3_0_clk),
    .D(_0088_),
    .RESET_B(net59),
    .Q(\internalDataflow.addressLowBusModule.busInputs[37] ));
 sky130_fd_sc_hd__dfrtp_1 _3097_ (.CLK(clknet_4_0_0_clk),
    .D(_0089_),
    .RESET_B(net59),
    .Q(\internalDataflow.addressLowBusModule.busInputs[38] ));
 sky130_fd_sc_hd__dfrtp_1 _3098_ (.CLK(clknet_4_2_0_clk),
    .D(_0090_),
    .RESET_B(net58),
    .Q(\internalDataflow.addressLowBusModule.busInputs[39] ));
 sky130_fd_sc_hd__dfrtp_4 _3099_ (.CLK(clknet_4_13_0_clk),
    .D(_0091_),
    .RESET_B(net66),
    .Q(\internalDataflow.addressHighBusModule.busInputs[16] ));
 sky130_fd_sc_hd__dfrtp_2 _3100_ (.CLK(clknet_4_13_0_clk),
    .D(_0092_),
    .RESET_B(net66),
    .Q(\internalDataflow.addressHighBusModule.busInputs[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3101_ (.CLK(clknet_4_11_0_clk),
    .D(_0093_),
    .RESET_B(net66),
    .Q(\internalDataflow.addressHighBusModule.busInputs[18] ));
 sky130_fd_sc_hd__dfrtp_2 _3102_ (.CLK(clknet_4_11_0_clk),
    .D(_0094_),
    .RESET_B(net64),
    .Q(\internalDataflow.addressHighBusModule.busInputs[19] ));
 sky130_fd_sc_hd__dfrtp_4 _3103_ (.CLK(clknet_4_10_0_clk),
    .D(_0095_),
    .RESET_B(net64),
    .Q(\internalDataflow.addressHighBusModule.busInputs[20] ));
 sky130_fd_sc_hd__dfrtp_2 _3104_ (.CLK(clknet_4_10_0_clk),
    .D(_0096_),
    .RESET_B(net64),
    .Q(\internalDataflow.addressHighBusModule.busInputs[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3105_ (.CLK(clknet_4_10_0_clk),
    .D(_0097_),
    .RESET_B(net64),
    .Q(\internalDataflow.addressHighBusModule.busInputs[22] ));
 sky130_fd_sc_hd__dfrtp_2 _3106_ (.CLK(clknet_4_9_0_clk),
    .D(_0098_),
    .RESET_B(net63),
    .Q(\internalDataflow.addressHighBusModule.busInputs[23] ));
 sky130_fd_sc_hd__dfrtp_1 _3107_ (.CLK(clknet_4_0_0_clk),
    .D(_0099_),
    .RESET_B(net57),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _3108_ (.CLK(clknet_4_8_0_clk),
    .D(_0100_),
    .RESET_B(net64),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _3109_ (.CLK(clknet_4_12_0_clk),
    .D(_0101_),
    .RESET_B(net70),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _3110_ (.CLK(clknet_4_11_0_clk),
    .D(_0102_),
    .RESET_B(net66),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _3111_ (.CLK(clknet_4_0_0_clk),
    .D(_0103_),
    .RESET_B(net57),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _3112_ (.CLK(clknet_4_2_0_clk),
    .D(_0104_),
    .RESET_B(net57),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _3113_ (.CLK(clknet_4_5_0_clk),
    .D(_0105_),
    .RESET_B(net69),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _3114_ (.CLK(clknet_4_11_0_clk),
    .D(_0106_),
    .RESET_B(net66),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _3115_ (.CLK(clknet_4_15_0_clk),
    .D(net73),
    .RESET_B(net71),
    .Q(\instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI ));
 sky130_fd_sc_hd__dfrtp_1 _3116_ (.CLK(clknet_4_15_0_clk),
    .D(\instructionLoader.interruptInjector.nmiSync.in ),
    .RESET_B(net71),
    .Q(\instructionLoader.interruptInjector.nmiSync.nextQ2 ));
 sky130_fd_sc_hd__dfrtp_1 _3117_ (.CLK(clknet_4_14_0_clk),
    .D(net74),
    .RESET_B(net71),
    .Q(\instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ ));
 sky130_fd_sc_hd__dfrtp_1 _3118_ (.CLK(clknet_4_14_0_clk),
    .D(\instructionLoader.interruptInjector.interruptRequest ),
    .RESET_B(net71),
    .Q(\instructionLoader.interruptInjector.irqSync.nextQ2 ));
 sky130_fd_sc_hd__dfrtp_4 _3119_ (.CLK(clknet_4_13_0_clk),
    .D(_0107_),
    .RESET_B(net70),
    .Q(\instructionLoader.interruptInjector.irqGenerated ));
 sky130_fd_sc_hd__dfrtp_4 _3120_ (.CLK(clknet_4_14_0_clk),
    .D(_0108_),
    .RESET_B(net71),
    .Q(\demux.nmi ));
 sky130_fd_sc_hd__dfrtp_1 _3121_ (.CLK(clknet_4_13_0_clk),
    .D(_0109_),
    .RESET_B(net70),
    .Q(\demux.setInterruptFlag ));
 sky130_fd_sc_hd__dfrtp_1 _3122_ (.CLK(clknet_4_5_0_clk),
    .D(_0110_),
    .RESET_B(net69),
    .Q(\negEdgeDetector.q1 ));
 sky130_fd_sc_hd__dfrtp_1 _3123_ (.CLK(clknet_4_14_0_clk),
    .D(_0111_),
    .RESET_B(net71),
    .Q(\instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ));
 sky130_fd_sc_hd__dfstp_2 _3124_ (.CLK(clknet_4_12_0_clk),
    .D(_0112_),
    .SET_B(net70),
    .Q(\instructionLoader.interruptInjector.resetDetected ));
 sky130_fd_sc_hd__dfrtp_1 _3125_ (.CLK(clknet_4_4_0_clk),
    .D(_0113_),
    .RESET_B(net69),
    .Q(\free_carry_ff.freeCarry ));
 sky130_fd_sc_hd__dfstp_2 _3126_ (.CLK(clknet_4_6_0_clk),
    .D(_0013_),
    .SET_B(net67),
    .Q(\demux.state_machine.timeState[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3127_ (.CLK(clknet_4_6_0_clk),
    .D(_0014_),
    .RESET_B(net69),
    .Q(\demux.state_machine.timeState[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3128_ (.CLK(clknet_4_5_0_clk),
    .D(_0015_),
    .RESET_B(net69),
    .Q(\demux.state_machine.timeState[2] ));
 sky130_fd_sc_hd__dfrtp_2 _3129_ (.CLK(clknet_4_6_0_clk),
    .D(_0016_),
    .RESET_B(net67),
    .Q(\demux.state_machine.timeState[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3130_ (.CLK(clknet_4_6_0_clk),
    .D(_0017_),
    .RESET_B(net69),
    .Q(\demux.state_machine.timeState[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3131_ (.CLK(clknet_4_5_0_clk),
    .D(_0018_),
    .RESET_B(net69),
    .Q(\demux.state_machine.timeState[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3132_ (.CLK(clknet_4_5_0_clk),
    .D(_0019_),
    .RESET_B(net69),
    .Q(\demux.state_machine.timeState[6] ));
 sky130_fd_sc_hd__dfrtp_2 _3133_ (.CLK(clknet_4_12_0_clk),
    .D(\internalDataflow.psr.processStatusReg.stat_buf_nxt[0] ),
    .RESET_B(net65),
    .Q(\demux.PSR_C ));
 sky130_fd_sc_hd__dfrtp_2 _3134_ (.CLK(clknet_4_12_0_clk),
    .D(\internalDataflow.psr.processStatusReg.stat_buf_nxt[1] ),
    .RESET_B(net65),
    .Q(\demux.PSR_Z ));
 sky130_fd_sc_hd__dfrtp_2 _3135_ (.CLK(clknet_4_12_0_clk),
    .D(\internalDataflow.psr.processStatusReg.stat_buf_nxt[2] ),
    .RESET_B(net70),
    .Q(\instructionLoader.interruptInjector.processStatusRegIFlag ));
 sky130_fd_sc_hd__dfrtp_4 _3136_ (.CLK(clknet_4_12_0_clk),
    .D(\internalDataflow.psr.processStatusReg.stat_buf_nxt[3] ),
    .RESET_B(net65),
    .Q(\internalDataflow.dataBusModule.busInputs[43] ));
 sky130_fd_sc_hd__dfrtp_4 _3137_ (.CLK(clknet_4_4_0_clk),
    .D(\internalDataflow.psr.processStatusReg.stat_buf_nxt[6] ),
    .RESET_B(net60),
    .Q(\demux.PSR_V ));
 sky130_fd_sc_hd__dfrtp_1 _3138_ (.CLK(clknet_4_15_0_clk),
    .D(_0020_),
    .RESET_B(net71),
    .Q(\demux.state_machine.currentInstruction[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3139_ (.CLK(clknet_4_15_0_clk),
    .D(_0021_),
    .RESET_B(net71),
    .Q(\demux.state_machine.currentInstruction[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3140_ (.CLK(clknet_4_15_0_clk),
    .D(_0022_),
    .RESET_B(net72),
    .Q(\demux.state_machine.currentInstruction[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3141_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .RESET_B(net72),
    .Q(\demux.state_machine.currentInstruction[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3142_ (.CLK(clknet_4_15_0_clk),
    .D(_0024_),
    .RESET_B(net72),
    .Q(\demux.state_machine.currentInstruction[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3143_ (.CLK(clknet_4_15_0_clk),
    .D(_0025_),
    .RESET_B(net72),
    .Q(\demux.state_machine.currentInstruction[5] ));
 sky130_fd_sc_hd__dfrtp_2 _3144_ (.CLK(clknet_4_4_0_clk),
    .D(_0114_),
    .RESET_B(net60),
    .Q(\branch_ff.branchForward ));
 sky130_fd_sc_hd__dfstp_1 _3145_ (.CLK(clknet_4_6_0_clk),
    .D(_0115_),
    .SET_B(net67),
    .Q(\demux.isAddressing ));
 sky130_fd_sc_hd__dfrtp_2 _3146_ (.CLK(clknet_4_4_0_clk),
    .D(_0116_),
    .RESET_B(net60),
    .Q(\branch_ff.branchBackward ));
 sky130_fd_sc_hd__dfrtp_1 _3147_ (.CLK(clknet_4_9_0_clk),
    .D(_0117_),
    .RESET_B(net65),
    .Q(\demux.PSR_N ));
 sky130_fd_sc_hd__buf_2 _3148_ (.A(clknet_4_1_0_clk),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net61),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net61),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net12),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net66),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net12),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net72),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net72),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net72),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net12),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\instructionLoader.interruptInjector.nmiSync.nextQ2 ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\internalDataflow.addressLowBusModule.busInputs[27] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\internalDataflow.addressLowBusModule.busInputs[31] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\demux.state_machine.timeState[3] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\demux.state_machine.currentAddress[3] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\demux.state_machine.currentAddress[10] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net39),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net35),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\negEdgeDetector.q1 ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\instructionLoader.interruptInjector.irqGenerated ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net19),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\instructionLoader.interruptInjector.irqSync.nextQ2 ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\demux.setInterruptFlag ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\internalDataflow.stackBusModule.busInputs[34] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\branch_ff.branchForward ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\branch_ff.branchBackward ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\internalDataflow.addressLowBusModule.busInputs[25] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net24),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\pulse_slower.currentEnableState[0] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\internalDataflow.stackBusModule.busInputs[37] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\internalDataflow.stackBusModule.busInputs[46] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\demux.state_machine.currentAddress[5] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net26),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net16),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\internalDataflow.stackBusModule.busInputs[45] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\internalDataflow.stackBusModule.busInputs[33] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\internalDataflow.stackBusModule.busInputs[42] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\internalDataflow.stackBusModule.busInputs[35] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\internalDataflow.stackBusModule.busInputs[44] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net18),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\internalDataflow.stackBusModule.busInputs[38] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\internalDataflow.stackBusModule.busInputs[43] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net29),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\demux.state_machine.currentAddress[8] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\internalDataflow.addressLowBusModule.busInputs[29] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\demux.state_machine.currentAddress[9] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\internalDataflow.stackBusModule.busInputs[36] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net21),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net36),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net37),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\free_carry_ff.freeCarry ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\internalDataflow.addressHighBusModule.busInputs[22] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\internalDataflow.addressLowBusModule.busInputs[22] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net23),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net27),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net30),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net22),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\internalDataflow.addressHighBusModule.busInputs[21] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net32),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net20),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\internalDataflow.stackBusModule.busInputs[41] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\internalDataflow.addressLowBusModule.busInputs[30] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\internalDataflow.addressHighBusModule.busInputs[18] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\internalDataflow.stackBusModule.busInputs[39] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\demux.state_machine.currentAddress[2] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\internalDataflow.addressHighBusModule.busInputs[20] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\internalDataflow.addressLowBusModule.busInputs[21] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net25),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\internalDataflow.addressLowBusModule.busInputs[24] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\demux.state_machine.currentAddress[4] ),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input1 (.A(dataBusEnable),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(interruptRequest),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(nonMaskableInterrupt),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(nrst),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(ready),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(setOverflow),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(dataBusInput[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(dataBusInput[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(dataBusInput[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(dataBusInput[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(dataBusInput[4]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(dataBusInput[5]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(dataBusInput[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(dataBusInput[7]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 max_cap1 (.A(_1312_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 max_cap44 (.A(_0270_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 max_cap46 (.A(_0119_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 max_cap47 (.A(_1387_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 max_cap48 (.A(_1312_),
    .X(net48));
 sky130_fd_sc_hd__buf_1 max_cap49 (.A(net135),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 max_cap50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_1 max_cap52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_1 max_cap54 (.A(_0989_),
    .X(net54));
 sky130_fd_sc_hd__buf_1 max_cap56 (.A(_0947_),
    .X(net56));
 sky130_fd_sc_hd__buf_1 output15 (.A(net15),
    .X(M10ClkOut));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(addressBusHigh[0]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(addressBusHigh[1]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(addressBusHigh[2]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(addressBusHigh[3]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(addressBusHigh[4]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(addressBusHigh[5]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(addressBusHigh[6]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(addressBusHigh[7]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(addressBusLow[0]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(addressBusLow[1]));
 sky130_fd_sc_hd__clkbuf_4 output26 (.A(net26),
    .X(addressBusLow[2]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(addressBusLow[3]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(addressBusLow[4]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(addressBusLow[5]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(addressBusLow[6]));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net31),
    .X(addressBusLow[7]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(dataBusOutput[0]));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net33),
    .X(dataBusOutput[1]));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net34),
    .X(dataBusOutput[2]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(dataBusOutput[3]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(dataBusOutput[4]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(dataBusOutput[5]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(dataBusOutput[6]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(dataBusOutput[7]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(dataBusSelect));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(functionalClockOut));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(readNotWrite));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(sync));
 sky130_fd_sc_hd__buf_1 wire2 (.A(_1335_),
    .X(net135));
 sky130_fd_sc_hd__buf_2 wire45 (.A(_0403_),
    .X(net45));
 sky130_fd_sc_hd__buf_1 wire51 (.A(_1340_),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire53 (.A(_0895_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 wire55 (.A(_0955_),
    .X(net55));
endmodule

