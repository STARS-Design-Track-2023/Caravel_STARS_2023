magic
tech sky130A
magscale 1 2
timestamp 1693969485
<< obsli1 >>
rect 1104 2159 52532 53329
<< obsm1 >>
rect 14 2128 53530 53360
<< metal2 >>
rect 6458 55024 6514 55824
rect 18050 55024 18106 55824
rect 30286 55024 30342 55824
rect 41878 55024 41934 55824
rect 53470 55024 53526 55824
rect 18 0 74 800
rect 11610 0 11666 800
rect 23202 0 23258 800
rect 35438 0 35494 800
rect 47030 0 47086 800
<< obsm2 >>
rect 20 54968 6402 55024
rect 6570 54968 17994 55024
rect 18162 54968 30230 55024
rect 30398 54968 41822 55024
rect 41990 54968 53414 55024
rect 20 856 53524 54968
rect 130 800 11554 856
rect 11722 800 23146 856
rect 23314 800 35382 856
rect 35550 800 46974 856
rect 47142 800 53524 856
<< metal3 >>
rect 0 49648 800 49768
rect 52880 42848 53680 42968
rect 0 37408 800 37528
rect 52880 30608 53680 30728
rect 0 24488 800 24608
rect 52880 17688 53680 17808
rect 0 12248 800 12368
rect 52880 5448 53680 5568
<< obsm3 >>
rect 800 49848 52880 53345
rect 880 49568 52880 49848
rect 800 43048 52880 49568
rect 800 42768 52800 43048
rect 800 37608 52880 42768
rect 880 37328 52880 37608
rect 800 30808 52880 37328
rect 800 30528 52800 30808
rect 800 24688 52880 30528
rect 880 24408 52880 24688
rect 800 17888 52880 24408
rect 800 17608 52800 17888
rect 800 12448 52880 17608
rect 880 12168 52880 12448
rect 800 5648 52880 12168
rect 800 5368 52800 5648
rect 800 2143 52880 5368
<< metal4 >>
rect 4208 2128 4528 53360
rect 19568 2128 19888 53360
rect 34928 2128 35248 53360
rect 50288 2128 50608 53360
<< obsm4 >>
rect 9995 6427 19488 48381
rect 19968 6427 20181 48381
<< labels >>
rlabel metal3 s 52880 5448 53680 5568 6 PWM_o
port 1 nsew signal output
rlabel metal3 s 52880 42848 53680 42968 6 clk
port 2 nsew signal input
rlabel metal2 s 30286 55024 30342 55824 6 modes
port 3 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 octaves
port 4 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 pb[0]
port 5 nsew signal input
rlabel metal2 s 18050 55024 18106 55824 6 pb[10]
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 pb[11]
port 7 nsew signal input
rlabel metal2 s 53470 55024 53526 55824 6 pb[12]
port 8 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 pb[1]
port 9 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 pb[2]
port 10 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 pb[3]
port 11 nsew signal input
rlabel metal3 s 52880 30608 53680 30728 6 pb[4]
port 12 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 pb[5]
port 13 nsew signal input
rlabel metal2 s 41878 55024 41934 55824 6 pb[6]
port 14 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 pb[7]
port 15 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 pb[8]
port 16 nsew signal input
rlabel metal2 s 6458 55024 6514 55824 6 pb[9]
port 17 nsew signal input
rlabel metal3 s 52880 17688 53680 17808 6 reset
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 53360 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 53360 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 53360 6 vssd1
port 20 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 53360 6 vssd1
port 20 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 53680 55824
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7350778
string GDS_FILE /home/designer-25/CUP/openlane/Synthia/runs/23_09_05_20_00/results/signoff/Synthia.magic.gds
string GDS_START 915390
<< end >>

