magic
tech sky130A
magscale 1 2
timestamp 1693932456
<< viali >>
rect 1409 45985 1443 46019
rect 21833 45985 21867 46019
rect 22293 45985 22327 46019
rect 1685 45917 1719 45951
rect 6561 45917 6595 45951
rect 9873 45917 9907 45951
rect 14841 45917 14875 45951
rect 14933 45917 14967 45951
rect 22201 45917 22235 45951
rect 23949 45917 23983 45951
rect 27629 45917 27663 45951
rect 28365 45917 28399 45951
rect 33149 45917 33183 45951
rect 42165 45917 42199 45951
rect 14565 45849 14599 45883
rect 41981 45849 42015 45883
rect 6745 45781 6779 45815
rect 9321 45781 9355 45815
rect 15117 45781 15151 45815
rect 24133 45781 24167 45815
rect 27537 45781 27571 45815
rect 28181 45781 28215 45815
rect 32965 45781 32999 45815
rect 22937 45577 22971 45611
rect 27721 45577 27755 45611
rect 27889 45577 27923 45611
rect 9505 45509 9539 45543
rect 15853 45509 15887 45543
rect 25421 45509 25455 45543
rect 28089 45509 28123 45543
rect 8861 45441 8895 45475
rect 9597 45441 9631 45475
rect 10609 45441 10643 45475
rect 11713 45441 11747 45475
rect 13277 45441 13311 45475
rect 13544 45441 13578 45475
rect 16037 45441 16071 45475
rect 17049 45441 17083 45475
rect 18429 45441 18463 45475
rect 22017 45441 22051 45475
rect 24041 45441 24075 45475
rect 24225 45441 24259 45475
rect 25145 45441 25179 45475
rect 9781 45373 9815 45407
rect 9965 45373 9999 45407
rect 15301 45373 15335 45407
rect 17141 45373 17175 45407
rect 17233 45373 17267 45407
rect 18061 45373 18095 45407
rect 23489 45373 23523 45407
rect 27537 45373 27571 45407
rect 29653 45373 29687 45407
rect 29929 45373 29963 45407
rect 30573 45373 30607 45407
rect 9137 45305 9171 45339
rect 14657 45305 14691 45339
rect 16681 45305 16715 45339
rect 9045 45237 9079 45271
rect 11529 45237 11563 45271
rect 14749 45237 14783 45271
rect 15761 45237 15795 45271
rect 16221 45237 16255 45271
rect 17509 45237 17543 45271
rect 18245 45237 18279 45271
rect 22661 45237 22695 45271
rect 24041 45237 24075 45271
rect 25053 45237 25087 45271
rect 25513 45237 25547 45271
rect 26985 45237 27019 45271
rect 27905 45237 27939 45271
rect 28181 45237 28215 45271
rect 30021 45237 30055 45271
rect 9210 45033 9244 45067
rect 11332 45033 11366 45067
rect 13645 45033 13679 45067
rect 17588 45033 17622 45067
rect 27997 45033 28031 45067
rect 29377 45033 29411 45067
rect 14933 44965 14967 44999
rect 23949 44965 23983 44999
rect 8953 44897 8987 44931
rect 11069 44897 11103 44931
rect 12817 44897 12851 44931
rect 13461 44897 13495 44931
rect 14289 44897 14323 44931
rect 14381 44897 14415 44931
rect 16957 44897 16991 44931
rect 21649 44897 21683 44931
rect 23121 44897 23155 44931
rect 24685 44897 24719 44931
rect 28641 44897 28675 44931
rect 29101 44897 29135 44931
rect 8769 44829 8803 44863
rect 13829 44829 13863 44863
rect 15117 44829 15151 44863
rect 17233 44829 17267 44863
rect 17325 44829 17359 44863
rect 21373 44829 21407 44863
rect 23305 44829 23339 44863
rect 24225 44829 24259 44863
rect 24409 44829 24443 44863
rect 26249 44829 26283 44863
rect 29009 44829 29043 44863
rect 23857 44761 23891 44795
rect 23949 44761 23983 44795
rect 26525 44761 26559 44795
rect 8585 44693 8619 44727
rect 10701 44693 10735 44727
rect 12909 44693 12943 44727
rect 14473 44693 14507 44727
rect 14841 44693 14875 44727
rect 15485 44693 15519 44727
rect 19073 44693 19107 44727
rect 24133 44693 24167 44727
rect 26157 44693 26191 44727
rect 28089 44693 28123 44727
rect 9689 44489 9723 44523
rect 9781 44489 9815 44523
rect 10149 44489 10183 44523
rect 10977 44489 11011 44523
rect 11345 44489 11379 44523
rect 11621 44489 11655 44523
rect 11989 44489 12023 44523
rect 16497 44489 16531 44523
rect 17049 44489 17083 44523
rect 18245 44489 18279 44523
rect 23581 44489 23615 44523
rect 23857 44489 23891 44523
rect 25421 44489 25455 44523
rect 25973 44489 26007 44523
rect 26702 44489 26736 44523
rect 10885 44421 10919 44455
rect 18582 44421 18616 44455
rect 22109 44421 22143 44455
rect 24133 44421 24167 44455
rect 24869 44421 24903 44455
rect 26801 44421 26835 44455
rect 27261 44421 27295 44455
rect 8309 44353 8343 44387
rect 8576 44353 8610 44387
rect 12633 44353 12667 44387
rect 12909 44353 12943 44387
rect 15384 44353 15418 44387
rect 18061 44353 18095 44387
rect 23765 44353 23799 44387
rect 23949 44353 23983 44387
rect 25605 44353 25639 44387
rect 25881 44353 25915 44387
rect 26065 44353 26099 44387
rect 26525 44353 26559 44387
rect 26617 44353 26651 44387
rect 44833 44353 44867 44387
rect 10241 44285 10275 44319
rect 10425 44285 10459 44319
rect 10793 44285 10827 44319
rect 12081 44285 12115 44319
rect 12265 44285 12299 44319
rect 12817 44285 12851 44319
rect 14473 44285 14507 44319
rect 14749 44285 14783 44319
rect 15117 44285 15151 44319
rect 17141 44285 17175 44319
rect 17325 44285 17359 44319
rect 18337 44285 18371 44319
rect 20361 44285 20395 44319
rect 21833 44285 21867 44319
rect 24777 44285 24811 44319
rect 25789 44285 25823 44319
rect 26985 44285 27019 44319
rect 44557 44285 44591 44319
rect 19717 44217 19751 44251
rect 25145 44217 25179 44251
rect 12449 44149 12483 44183
rect 13001 44149 13035 44183
rect 16681 44149 16715 44183
rect 19809 44149 19843 44183
rect 25329 44149 25363 44183
rect 28733 44149 28767 44183
rect 7389 43945 7423 43979
rect 10517 43945 10551 43979
rect 14105 43945 14139 43979
rect 15761 43945 15795 43979
rect 18337 43945 18371 43979
rect 19257 43945 19291 43979
rect 22201 43945 22235 43979
rect 23673 43945 23707 43979
rect 10609 43877 10643 43911
rect 9965 43809 9999 43843
rect 14657 43809 14691 43843
rect 18889 43809 18923 43843
rect 19809 43809 19843 43843
rect 22753 43809 22787 43843
rect 23397 43809 23431 43843
rect 25973 43809 26007 43843
rect 30297 43809 30331 43843
rect 32137 43809 32171 43843
rect 33609 43809 33643 43843
rect 11989 43741 12023 43775
rect 14473 43741 14507 43775
rect 15393 43741 15427 43775
rect 15945 43741 15979 43775
rect 18797 43741 18831 43775
rect 19625 43741 19659 43775
rect 22201 43741 22235 43775
rect 22385 43741 22419 43775
rect 25237 43741 25271 43775
rect 33885 43741 33919 43775
rect 7113 43673 7147 43707
rect 11744 43673 11778 43707
rect 15117 43673 15151 43707
rect 23657 43673 23691 43707
rect 23857 43673 23891 43707
rect 26249 43673 26283 43707
rect 30573 43673 30607 43707
rect 14565 43605 14599 43639
rect 18705 43605 18739 43639
rect 19717 43605 19751 43639
rect 23489 43605 23523 43639
rect 25421 43605 25455 43639
rect 27721 43605 27755 43639
rect 32045 43605 32079 43639
rect 7757 43401 7791 43435
rect 7665 43333 7699 43367
rect 8401 43333 8435 43367
rect 27445 43333 27479 43367
rect 8304 43265 8338 43299
rect 8493 43265 8527 43299
rect 8676 43265 8710 43299
rect 8769 43265 8803 43299
rect 13369 43265 13403 43299
rect 20729 43265 20763 43299
rect 27261 43265 27295 43299
rect 33885 43265 33919 43299
rect 35817 43265 35851 43299
rect 6929 43197 6963 43231
rect 9505 43197 9539 43231
rect 10149 43197 10183 43231
rect 16681 43197 16715 43231
rect 33977 43197 34011 43231
rect 34253 43197 34287 43231
rect 7481 43061 7515 43095
rect 8125 43061 8159 43095
rect 13185 43061 13219 43095
rect 17325 43061 17359 43095
rect 19441 43061 19475 43095
rect 27077 43061 27111 43095
rect 32413 43061 32447 43095
rect 35725 43061 35759 43095
rect 36001 43061 36035 43095
rect 7131 42857 7165 42891
rect 14841 42857 14875 42891
rect 16221 42857 16255 42891
rect 17797 42857 17831 42891
rect 32781 42857 32815 42891
rect 7573 42721 7607 42755
rect 8125 42721 8159 42755
rect 12633 42721 12667 42755
rect 13829 42721 13863 42755
rect 16313 42721 16347 42755
rect 23029 42721 23063 42755
rect 23213 42721 23247 42755
rect 24409 42721 24443 42755
rect 30205 42721 30239 42755
rect 35265 42721 35299 42755
rect 3893 42653 3927 42687
rect 4077 42653 4111 42687
rect 4905 42653 4939 42687
rect 7389 42653 7423 42687
rect 7849 42653 7883 42687
rect 13277 42653 13311 42687
rect 13461 42653 13495 42687
rect 13645 42653 13679 42687
rect 14657 42653 14691 42687
rect 15393 42653 15427 42687
rect 15577 42653 15611 42687
rect 15725 42653 15759 42687
rect 16083 42653 16117 42687
rect 18061 42653 18095 42687
rect 18153 42653 18187 42687
rect 18337 42653 18371 42687
rect 18797 42653 18831 42687
rect 19349 42653 19383 42687
rect 21281 42653 21315 42687
rect 24041 42653 24075 42687
rect 30297 42653 30331 42687
rect 30757 42653 30791 42687
rect 30941 42653 30975 42687
rect 32045 42653 32079 42687
rect 32965 42653 32999 42687
rect 33149 42653 33183 42687
rect 33267 42653 33301 42687
rect 33425 42653 33459 42687
rect 33517 42653 33551 42687
rect 34069 42653 34103 42687
rect 9045 42585 9079 42619
rect 10793 42585 10827 42619
rect 12357 42585 12391 42619
rect 12725 42585 12759 42619
rect 15853 42585 15887 42619
rect 15945 42585 15979 42619
rect 21557 42585 21591 42619
rect 24685 42585 24719 42619
rect 27997 42585 28031 42619
rect 31401 42585 31435 42619
rect 33057 42585 33091 42619
rect 4261 42517 4295 42551
rect 5457 42517 5491 42551
rect 5641 42517 5675 42551
rect 8769 42517 8803 42551
rect 10885 42517 10919 42551
rect 14105 42517 14139 42551
rect 18521 42517 18555 42551
rect 18613 42517 18647 42551
rect 19993 42517 20027 42551
rect 23857 42517 23891 42551
rect 24225 42517 24259 42551
rect 26157 42517 26191 42551
rect 26709 42517 26743 42551
rect 30665 42517 30699 42551
rect 30941 42517 30975 42551
rect 34713 42517 34747 42551
rect 7021 42313 7055 42347
rect 8861 42313 8895 42347
rect 12173 42313 12207 42347
rect 13645 42313 13679 42347
rect 15577 42313 15611 42347
rect 16681 42313 16715 42347
rect 20913 42313 20947 42347
rect 22017 42313 22051 42347
rect 24685 42313 24719 42347
rect 31769 42313 31803 42347
rect 33977 42313 34011 42347
rect 34897 42313 34931 42347
rect 5825 42245 5859 42279
rect 6653 42245 6687 42279
rect 9229 42245 9263 42279
rect 12532 42245 12566 42279
rect 14013 42245 14047 42279
rect 23029 42245 23063 42279
rect 25145 42245 25179 42279
rect 33471 42245 33505 42279
rect 33609 42245 33643 42279
rect 33701 42245 33735 42279
rect 34713 42245 34747 42279
rect 3709 42177 3743 42211
rect 6377 42177 6411 42211
rect 6470 42177 6504 42211
rect 6745 42177 6779 42211
rect 6883 42177 6917 42211
rect 7481 42177 7515 42211
rect 7748 42177 7782 42211
rect 8953 42177 8987 42211
rect 10977 42177 11011 42211
rect 12265 42177 12299 42211
rect 15761 42177 15795 42211
rect 17693 42177 17727 42211
rect 17960 42177 17994 42211
rect 21925 42177 21959 42211
rect 22109 42177 22143 42211
rect 22201 42177 22235 42211
rect 22385 42177 22419 42211
rect 22661 42177 22695 42211
rect 22845 42177 22879 42211
rect 23765 42177 23799 42211
rect 23949 42177 23983 42211
rect 25053 42177 25087 42211
rect 26617 42177 26651 42211
rect 26801 42177 26835 42211
rect 26985 42177 27019 42211
rect 28825 42177 28859 42211
rect 31585 42177 31619 42211
rect 31861 42177 31895 42211
rect 32137 42177 32171 42211
rect 32321 42177 32355 42211
rect 33333 42177 33367 42211
rect 33793 42177 33827 42211
rect 34253 42177 34287 42211
rect 34897 42177 34931 42211
rect 34989 42177 35023 42211
rect 6101 42109 6135 42143
rect 10793 42109 10827 42143
rect 11529 42109 11563 42143
rect 13737 42109 13771 42143
rect 15945 42109 15979 42143
rect 17325 42109 17359 42143
rect 19165 42109 19199 42143
rect 19441 42109 19475 42143
rect 23581 42109 23615 42143
rect 25329 42109 25363 42143
rect 27261 42109 27295 42143
rect 29101 42109 29135 42143
rect 30573 42109 30607 42143
rect 31217 42109 31251 42143
rect 34161 42109 34195 42143
rect 23765 42041 23799 42075
rect 31401 42041 31435 42075
rect 34621 42041 34655 42075
rect 4261 41973 4295 42007
rect 4353 41973 4387 42007
rect 10701 41973 10735 42007
rect 11161 41973 11195 42007
rect 15485 41973 15519 42007
rect 19073 41973 19107 42007
rect 22201 41973 22235 42007
rect 22477 41973 22511 42007
rect 26709 41973 26743 42007
rect 28733 41973 28767 42007
rect 30665 41973 30699 42007
rect 32137 41973 32171 42007
rect 3617 41769 3651 41803
rect 4997 41769 5031 41803
rect 6469 41769 6503 41803
rect 8309 41769 8343 41803
rect 11529 41769 11563 41803
rect 12265 41769 12299 41803
rect 13093 41769 13127 41803
rect 17325 41769 17359 41803
rect 19073 41769 19107 41803
rect 19257 41769 19291 41803
rect 19993 41769 20027 41803
rect 23213 41769 23247 41803
rect 26801 41769 26835 41803
rect 29561 41769 29595 41803
rect 30941 41769 30975 41803
rect 31493 41769 31527 41803
rect 32321 41769 32355 41803
rect 33701 41769 33735 41803
rect 35633 41769 35667 41803
rect 7757 41701 7791 41735
rect 22937 41701 22971 41735
rect 32873 41701 32907 41735
rect 34253 41701 34287 41735
rect 2145 41633 2179 41667
rect 3801 41633 3835 41667
rect 5365 41633 5399 41667
rect 7389 41633 7423 41667
rect 9505 41633 9539 41667
rect 13645 41633 13679 41667
rect 18429 41633 18463 41667
rect 20545 41633 20579 41667
rect 28365 41633 28399 41667
rect 30205 41633 30239 41667
rect 32781 41633 32815 41667
rect 32965 41633 32999 41667
rect 1869 41565 1903 41599
rect 3985 41565 4019 41599
rect 4353 41565 4387 41599
rect 4501 41565 4535 41599
rect 4859 41565 4893 41599
rect 6101 41565 6135 41599
rect 6285 41565 6319 41599
rect 7573 41565 7607 41599
rect 8493 41565 8527 41599
rect 10149 41565 10183 41599
rect 11621 41565 11655 41599
rect 11714 41565 11748 41599
rect 11989 41565 12023 41599
rect 12086 41565 12120 41599
rect 13461 41565 13495 41599
rect 15945 41565 15979 41599
rect 19395 41565 19429 41599
rect 19533 41565 19567 41599
rect 19808 41565 19842 41599
rect 19901 41565 19935 41599
rect 21189 41565 21223 41599
rect 24593 41565 24627 41599
rect 26985 41565 27019 41599
rect 27169 41565 27203 41599
rect 27445 41565 27479 41599
rect 27813 41565 27847 41599
rect 29762 41575 29796 41609
rect 29929 41565 29963 41599
rect 30389 41565 30423 41599
rect 30573 41565 30607 41599
rect 30757 41565 30791 41599
rect 31033 41565 31067 41599
rect 31125 41565 31159 41599
rect 31309 41565 31343 41599
rect 31585 41565 31619 41599
rect 31861 41565 31895 41599
rect 32229 41565 32263 41599
rect 32413 41565 32447 41599
rect 32505 41565 32539 41599
rect 32689 41565 32723 41599
rect 33057 41565 33091 41599
rect 33885 41565 33919 41599
rect 34069 41565 34103 41599
rect 34161 41565 34195 41599
rect 34253 41565 34287 41599
rect 34437 41565 34471 41599
rect 34713 41565 34747 41599
rect 34897 41565 34931 41599
rect 4629 41497 4663 41531
rect 4721 41497 4755 41531
rect 10416 41497 10450 41531
rect 11897 41497 11931 41531
rect 14105 41497 14139 41531
rect 16190 41497 16224 41531
rect 18705 41497 18739 41531
rect 19625 41497 19659 41531
rect 21465 41497 21499 41531
rect 23029 41497 23063 41531
rect 27077 41497 27111 41531
rect 27307 41497 27341 41531
rect 29848 41497 29882 41531
rect 30067 41497 30101 41531
rect 30665 41497 30699 41531
rect 31677 41497 31711 41531
rect 33425 41497 33459 41531
rect 33609 41497 33643 41531
rect 34805 41497 34839 41531
rect 35523 41497 35557 41531
rect 4169 41429 4203 41463
rect 6009 41429 6043 41463
rect 8953 41429 8987 41463
rect 9321 41429 9355 41463
rect 9413 41429 9447 41463
rect 13553 41429 13587 41463
rect 15393 41429 15427 41463
rect 18613 41429 18647 41463
rect 23229 41429 23263 41463
rect 23397 41429 23431 41463
rect 24869 41429 24903 41463
rect 31585 41429 31619 41463
rect 31953 41429 31987 41463
rect 33241 41429 33275 41463
rect 3065 41225 3099 41259
rect 9137 41225 9171 41259
rect 10517 41225 10551 41259
rect 11897 41225 11931 41259
rect 15209 41225 15243 41259
rect 15761 41225 15795 41259
rect 18797 41225 18831 41259
rect 21557 41225 21591 41259
rect 23581 41225 23615 41259
rect 28089 41225 28123 41259
rect 30205 41225 30239 41259
rect 30481 41225 30515 41259
rect 30573 41225 30607 41259
rect 34161 41225 34195 41259
rect 34529 41225 34563 41259
rect 4905 41157 4939 41191
rect 14381 41157 14415 41191
rect 14473 41157 14507 41191
rect 20545 41157 20579 41191
rect 24133 41157 24167 41191
rect 28641 41157 28675 41191
rect 28825 41157 28859 41191
rect 30941 41157 30975 41191
rect 34069 41157 34103 41191
rect 35633 41157 35667 41191
rect 28411 41123 28445 41157
rect 3980 41089 4014 41123
rect 4077 41089 4111 41123
rect 4169 41089 4203 41123
rect 4352 41089 4386 41123
rect 4445 41089 4479 41123
rect 4537 41089 4571 41123
rect 4685 41089 4719 41123
rect 4813 41089 4847 41123
rect 5002 41089 5036 41123
rect 5457 41089 5491 41123
rect 9689 41089 9723 41123
rect 10701 41089 10735 41123
rect 13461 41089 13495 41123
rect 14284 41089 14318 41123
rect 14656 41089 14690 41123
rect 14749 41089 14783 41123
rect 15025 41089 15059 41123
rect 18705 41089 18739 41123
rect 20269 41089 20303 41123
rect 21189 41089 21223 41123
rect 21465 41089 21499 41123
rect 21649 41089 21683 41123
rect 22017 41089 22051 41123
rect 22385 41089 22419 41123
rect 22845 41089 22879 41123
rect 23029 41089 23063 41123
rect 23213 41089 23247 41123
rect 23397 41089 23431 41123
rect 23758 41089 23792 41123
rect 23857 41089 23891 41123
rect 27905 41089 27939 41123
rect 28181 41089 28215 41123
rect 30205 41089 30239 41123
rect 30665 41089 30699 41123
rect 30757 41089 30791 41123
rect 31493 41089 31527 41123
rect 31677 41089 31711 41123
rect 32137 41089 32171 41123
rect 32312 41089 32346 41123
rect 32413 41089 32447 41123
rect 32597 41089 32631 41123
rect 33701 41089 33735 41123
rect 33885 41089 33919 41123
rect 34161 41089 34195 41123
rect 34345 41089 34379 41123
rect 34437 41089 34471 41123
rect 34621 41089 34655 41123
rect 3709 41021 3743 41055
rect 5273 41021 5307 41055
rect 5641 41021 5675 41055
rect 8125 41021 8159 41055
rect 11989 41021 12023 41055
rect 12173 41021 12207 41055
rect 13185 41021 13219 41055
rect 15853 41021 15887 41055
rect 16037 41021 16071 41055
rect 21833 41021 21867 41055
rect 22201 41021 22235 41055
rect 23305 41021 23339 41055
rect 24409 41021 24443 41055
rect 24685 41021 24719 41055
rect 26157 41021 26191 41055
rect 27537 41021 27571 41055
rect 29101 41021 29135 41055
rect 31125 41021 31159 41055
rect 31401 41021 31435 41055
rect 31585 41021 31619 41055
rect 32229 41021 32263 41055
rect 5181 40953 5215 40987
rect 11529 40953 11563 40987
rect 14105 40953 14139 40987
rect 15393 40953 15427 40987
rect 3801 40885 3835 40919
rect 7481 40885 7515 40919
rect 20913 40885 20947 40919
rect 22661 40885 22695 40919
rect 22937 40885 22971 40919
rect 26985 40885 27019 40919
rect 27721 40885 27755 40919
rect 28273 40885 28307 40919
rect 28457 40885 28491 40919
rect 30297 40885 30331 40919
rect 31217 40885 31251 40919
rect 32505 40885 32539 40919
rect 35541 40885 35575 40919
rect 4813 40681 4847 40715
rect 6377 40681 6411 40715
rect 25881 40681 25915 40715
rect 3341 40613 3375 40647
rect 12173 40613 12207 40647
rect 35817 40613 35851 40647
rect 1593 40545 1627 40579
rect 5365 40545 5399 40579
rect 6469 40545 6503 40579
rect 6745 40545 6779 40579
rect 8217 40545 8251 40579
rect 8677 40545 8711 40579
rect 10977 40545 11011 40579
rect 12817 40545 12851 40579
rect 16497 40545 16531 40579
rect 18245 40545 18279 40579
rect 26525 40545 26559 40579
rect 37381 40545 37415 40579
rect 4629 40477 4663 40511
rect 5733 40477 5767 40511
rect 8493 40477 8527 40511
rect 9505 40477 9539 40511
rect 11161 40477 11195 40511
rect 11345 40477 11379 40511
rect 11529 40477 11563 40511
rect 11622 40477 11656 40511
rect 11994 40477 12028 40511
rect 13737 40477 13771 40511
rect 18889 40477 18923 40511
rect 20177 40477 20211 40511
rect 23857 40477 23891 40511
rect 26065 40477 26099 40511
rect 26157 40477 26191 40511
rect 26249 40477 26283 40511
rect 26893 40477 26927 40511
rect 27261 40477 27295 40511
rect 27537 40477 27571 40511
rect 35265 40477 35299 40511
rect 35633 40477 35667 40511
rect 37657 40477 37691 40511
rect 1869 40409 1903 40443
rect 11805 40409 11839 40443
rect 11897 40409 11931 40443
rect 17969 40409 18003 40443
rect 18337 40409 18371 40443
rect 26367 40409 26401 40443
rect 35449 40409 35483 40443
rect 35541 40409 35575 40443
rect 4077 40341 4111 40375
rect 8309 40341 8343 40375
rect 8953 40341 8987 40375
rect 12265 40341 12299 40375
rect 13921 40341 13955 40375
rect 20821 40341 20855 40375
rect 24041 40341 24075 40375
rect 26709 40341 26743 40375
rect 27169 40341 27203 40375
rect 27445 40341 27479 40375
rect 35909 40341 35943 40375
rect 2881 40137 2915 40171
rect 8217 40137 8251 40171
rect 11989 40137 12023 40171
rect 13461 40137 13495 40171
rect 15301 40137 15335 40171
rect 16497 40137 16531 40171
rect 23213 40137 23247 40171
rect 27997 40137 28031 40171
rect 35265 40137 35299 40171
rect 35725 40137 35759 40171
rect 40601 40137 40635 40171
rect 3893 40069 3927 40103
rect 10793 40069 10827 40103
rect 13093 40069 13127 40103
rect 22385 40069 22419 40103
rect 23305 40069 23339 40103
rect 23857 40069 23891 40103
rect 24041 40069 24075 40103
rect 27629 40069 27663 40103
rect 3617 40001 3651 40035
rect 6377 40001 6411 40035
rect 8396 40001 8430 40035
rect 8493 40001 8527 40035
rect 8585 40001 8619 40035
rect 8713 40001 8747 40035
rect 8861 40001 8895 40035
rect 15853 40001 15887 40035
rect 15946 40001 15980 40035
rect 16129 40001 16163 40035
rect 16221 40001 16255 40035
rect 16318 40001 16352 40035
rect 17049 40001 17083 40035
rect 18337 40001 18371 40035
rect 18521 40001 18555 40035
rect 20545 40001 20579 40035
rect 24225 40001 24259 40035
rect 26801 40001 26835 40035
rect 27169 40001 27203 40035
rect 27353 40001 27387 40035
rect 27813 40001 27847 40035
rect 28089 40001 28123 40035
rect 33333 40001 33367 40035
rect 34161 40001 34195 40035
rect 34897 40001 34931 40035
rect 36277 40001 36311 40035
rect 3525 39933 3559 39967
rect 5365 39933 5399 39967
rect 5457 39933 5491 39967
rect 6653 39933 6687 39967
rect 8125 39933 8159 39967
rect 9321 39933 9355 39967
rect 11069 39933 11103 39967
rect 12541 39933 12575 39967
rect 12817 39933 12851 39967
rect 13001 39933 13035 39967
rect 13553 39933 13587 39967
rect 13829 39933 13863 39967
rect 18705 39933 18739 39967
rect 20269 39933 20303 39967
rect 20913 39933 20947 39967
rect 24409 39933 24443 39967
rect 26709 39933 26743 39967
rect 27261 39933 27295 39967
rect 27445 39933 27479 39967
rect 34253 39933 34287 39967
rect 34989 39933 35023 39967
rect 38853 39933 38887 39967
rect 39129 39933 39163 39967
rect 22109 39865 22143 39899
rect 6101 39797 6135 39831
rect 17601 39797 17635 39831
rect 18797 39797 18831 39831
rect 21557 39797 21591 39831
rect 23765 39797 23799 39831
rect 26433 39797 26467 39831
rect 26801 39797 26835 39831
rect 26985 39797 27019 39831
rect 4261 39593 4295 39627
rect 6929 39593 6963 39627
rect 9689 39593 9723 39627
rect 12357 39593 12391 39627
rect 16773 39593 16807 39627
rect 20545 39593 20579 39627
rect 26157 39593 26191 39627
rect 28273 39593 28307 39627
rect 30205 39525 30239 39559
rect 36185 39525 36219 39559
rect 10057 39457 10091 39491
rect 15393 39457 15427 39491
rect 24409 39457 24443 39491
rect 26525 39457 26559 39491
rect 26801 39457 26835 39491
rect 29653 39457 29687 39491
rect 32229 39457 32263 39491
rect 37749 39457 37783 39491
rect 41613 39457 41647 39491
rect 3065 39389 3099 39423
rect 5549 39389 5583 39423
rect 7573 39389 7607 39423
rect 7844 39389 7878 39423
rect 8216 39389 8250 39423
rect 8309 39389 8343 39423
rect 8953 39389 8987 39423
rect 9873 39389 9907 39423
rect 10977 39389 11011 39423
rect 12449 39389 12483 39423
rect 15117 39389 15151 39423
rect 17693 39389 17727 39423
rect 19625 39389 19659 39423
rect 22293 39389 22327 39423
rect 26433 39389 26467 39423
rect 29837 39389 29871 39423
rect 30113 39389 30147 39423
rect 30297 39389 30331 39423
rect 35633 39389 35667 39423
rect 36001 39389 36035 39423
rect 38025 39389 38059 39423
rect 39129 39389 39163 39423
rect 39405 39389 39439 39423
rect 39497 39389 39531 39423
rect 39865 39389 39899 39423
rect 42257 39389 42291 39423
rect 7941 39321 7975 39355
rect 8033 39321 8067 39355
rect 11244 39321 11278 39355
rect 12716 39321 12750 39355
rect 15638 39321 15672 39355
rect 22017 39321 22051 39355
rect 22477 39321 22511 39355
rect 24685 39321 24719 39355
rect 31953 39321 31987 39355
rect 35817 39321 35851 39355
rect 35909 39321 35943 39355
rect 39313 39321 39347 39355
rect 40141 39321 40175 39355
rect 2513 39253 2547 39287
rect 7665 39253 7699 39287
rect 9597 39253 9631 39287
rect 13829 39253 13863 39287
rect 15301 39253 15335 39287
rect 17141 39253 17175 39287
rect 20269 39253 20303 39287
rect 22753 39253 22787 39287
rect 26341 39253 26375 39287
rect 30021 39253 30055 39287
rect 30481 39253 30515 39287
rect 36277 39253 36311 39287
rect 39681 39253 39715 39287
rect 41705 39253 41739 39287
rect 2605 39049 2639 39083
rect 4169 39049 4203 39083
rect 8677 39049 8711 39083
rect 11529 39049 11563 39083
rect 12173 39049 12207 39083
rect 12909 39049 12943 39083
rect 13001 39049 13035 39083
rect 13461 39049 13495 39083
rect 14197 39049 14231 39083
rect 15577 39049 15611 39083
rect 15945 39049 15979 39083
rect 17141 39049 17175 39083
rect 20177 39049 20211 39083
rect 22477 39049 22511 39083
rect 24875 39049 24909 39083
rect 24961 39049 24995 39083
rect 26985 39049 27019 39083
rect 27879 39049 27913 39083
rect 28273 39049 28307 39083
rect 29561 39049 29595 39083
rect 31601 39049 31635 39083
rect 32413 39049 32447 39083
rect 34161 39049 34195 39083
rect 35449 39049 35483 39083
rect 36093 39049 36127 39083
rect 12265 38981 12299 39015
rect 19809 38981 19843 39015
rect 19901 38981 19935 39015
rect 28089 38981 28123 39015
rect 29929 38981 29963 39015
rect 30389 38981 30423 39015
rect 31401 38981 31435 39015
rect 33609 38981 33643 39015
rect 37289 38981 37323 39015
rect 2973 38913 3007 38947
rect 3433 38913 3467 38947
rect 4348 38913 4382 38947
rect 4445 38913 4479 38947
rect 4537 38913 4571 38947
rect 4720 38913 4754 38947
rect 4813 38913 4847 38947
rect 7205 38913 7239 38947
rect 7389 38913 7423 38947
rect 7573 38913 7607 38947
rect 8585 38913 8619 38947
rect 10057 38913 10091 38947
rect 11713 38913 11747 38947
rect 14013 38913 14047 38947
rect 14381 38913 14415 38947
rect 16037 38913 16071 38947
rect 17049 38913 17083 38947
rect 18061 38913 18095 38947
rect 18328 38913 18362 38947
rect 19533 38913 19567 38947
rect 19626 38913 19660 38947
rect 20039 38913 20073 38947
rect 20453 38913 20487 38947
rect 20637 38913 20671 38947
rect 20908 38913 20942 38947
rect 21005 38913 21039 38947
rect 21097 38913 21131 38947
rect 21280 38913 21314 38947
rect 21373 38913 21407 38947
rect 22569 38913 22603 38947
rect 22753 38913 22787 38947
rect 24041 38913 24075 38947
rect 24777 38913 24811 38947
rect 25053 38913 25087 38947
rect 27537 38913 27571 38947
rect 28365 38913 28399 38947
rect 29745 38913 29779 38947
rect 30205 38913 30239 38947
rect 30481 38913 30515 38947
rect 30665 38913 30699 38947
rect 32597 38913 32631 38947
rect 32873 38913 32907 38947
rect 32965 38913 32999 38947
rect 33149 38913 33183 38947
rect 33241 38913 33275 38947
rect 33333 38913 33367 38947
rect 34069 38913 34103 38947
rect 34437 38913 34471 38947
rect 34989 38913 35023 38947
rect 35725 38913 35759 38947
rect 36645 38913 36679 38947
rect 39957 38913 39991 38947
rect 3065 38845 3099 38879
rect 3157 38845 3191 38879
rect 3985 38845 4019 38879
rect 8861 38845 8895 38879
rect 9413 38845 9447 38879
rect 12357 38845 12391 38879
rect 12725 38845 12759 38879
rect 16129 38845 16163 38879
rect 17233 38845 17267 38879
rect 20269 38845 20303 38879
rect 21833 38845 21867 38879
rect 22937 38845 22971 38879
rect 23581 38845 23615 38879
rect 32505 38845 32539 38879
rect 32781 38845 32815 38879
rect 33977 38845 34011 38879
rect 34161 38845 34195 38879
rect 34897 38845 34931 38879
rect 35357 38845 35391 38879
rect 35449 38845 35483 38879
rect 39773 38845 39807 38879
rect 40233 38845 40267 38879
rect 11805 38777 11839 38811
rect 13369 38777 13403 38811
rect 19441 38777 19475 38811
rect 20729 38777 20763 38811
rect 33701 38777 33735 38811
rect 35633 38777 35667 38811
rect 39129 38777 39163 38811
rect 8217 38709 8251 38743
rect 16681 38709 16715 38743
rect 23029 38709 23063 38743
rect 24685 38709 24719 38743
rect 27721 38709 27755 38743
rect 27905 38709 27939 38743
rect 30021 38709 30055 38743
rect 30573 38709 30607 38743
rect 31585 38709 31619 38743
rect 31769 38709 31803 38743
rect 34069 38709 34103 38743
rect 34345 38709 34379 38743
rect 38577 38709 38611 38743
rect 41705 38709 41739 38743
rect 2973 38505 3007 38539
rect 5089 38505 5123 38539
rect 8769 38505 8803 38539
rect 17049 38505 17083 38539
rect 18613 38505 18647 38539
rect 24225 38505 24259 38539
rect 31217 38505 31251 38539
rect 33333 38505 33367 38539
rect 34069 38505 34103 38539
rect 35541 38505 35575 38539
rect 39129 38505 39163 38539
rect 40693 38505 40727 38539
rect 33057 38437 33091 38471
rect 39037 38437 39071 38471
rect 4997 38369 5031 38403
rect 7389 38369 7423 38403
rect 9505 38369 9539 38403
rect 15669 38369 15703 38403
rect 17417 38369 17451 38403
rect 18337 38369 18371 38403
rect 22477 38369 22511 38403
rect 22753 38369 22787 38403
rect 24961 38369 24995 38403
rect 32873 38369 32907 38403
rect 35081 38369 35115 38403
rect 40049 38369 40083 38403
rect 1593 38301 1627 38335
rect 6469 38301 6503 38335
rect 7113 38301 7147 38335
rect 9229 38301 9263 38335
rect 17233 38301 17267 38335
rect 18245 38301 18279 38335
rect 18797 38301 18831 38335
rect 19809 38301 19843 38335
rect 25513 38301 25547 38335
rect 29745 38301 29779 38335
rect 29837 38301 29871 38335
rect 30067 38301 30101 38335
rect 30205 38301 30239 38335
rect 30297 38301 30331 38335
rect 30849 38301 30883 38335
rect 31033 38301 31067 38335
rect 32597 38301 32631 38335
rect 32965 38301 32999 38335
rect 33425 38301 33459 38335
rect 33609 38301 33643 38335
rect 33885 38301 33919 38335
rect 34713 38301 34747 38335
rect 34897 38301 34931 38335
rect 35173 38301 35207 38335
rect 35357 38301 35391 38335
rect 35449 38301 35483 38335
rect 35633 38301 35667 38335
rect 36185 38301 36219 38335
rect 36645 38301 36679 38335
rect 36921 38301 36955 38335
rect 37037 38301 37071 38335
rect 37289 38301 37323 38335
rect 39313 38301 39347 38335
rect 39681 38301 39715 38335
rect 40785 38301 40819 38335
rect 42073 38301 42107 38335
rect 1860 38233 1894 38267
rect 6224 38233 6258 38267
rect 7634 38233 7668 38267
rect 9781 38233 9815 38267
rect 15936 38233 15970 38267
rect 25145 38233 25179 38267
rect 25973 38233 26007 38267
rect 29929 38233 29963 38267
rect 35265 38233 35299 38267
rect 36829 38233 36863 38267
rect 37565 38233 37599 38267
rect 39405 38233 39439 38267
rect 39497 38233 39531 38267
rect 41521 38233 41555 38267
rect 4353 38165 4387 38199
rect 7297 38165 7331 38199
rect 9413 38165 9447 38199
rect 11253 38165 11287 38199
rect 17785 38165 17819 38199
rect 18153 38165 18187 38199
rect 19257 38165 19291 38199
rect 24409 38165 24443 38199
rect 26249 38165 26283 38199
rect 29561 38165 29595 38199
rect 32689 38165 32723 38199
rect 36461 38165 36495 38199
rect 37197 38165 37231 38199
rect 41429 38165 41463 38199
rect 2145 37961 2179 37995
rect 4445 37961 4479 37995
rect 6745 37961 6779 37995
rect 8585 37961 8619 37995
rect 9045 37961 9079 37995
rect 9597 37961 9631 37995
rect 10057 37961 10091 37995
rect 15669 37961 15703 37995
rect 15945 37961 15979 37995
rect 17325 37961 17359 37995
rect 18797 37961 18831 37995
rect 21189 37961 21223 37995
rect 23213 37961 23247 37995
rect 29929 37961 29963 37995
rect 32774 37961 32808 37995
rect 39865 37961 39899 37995
rect 9965 37893 9999 37927
rect 12265 37893 12299 37927
rect 19717 37893 19751 37927
rect 28457 37893 28491 37927
rect 30205 37893 30239 37927
rect 39037 37893 39071 37927
rect 2329 37825 2363 37859
rect 2789 37825 2823 37859
rect 3065 37825 3099 37859
rect 3321 37825 3355 37859
rect 4896 37825 4930 37859
rect 7472 37825 7506 37859
rect 11989 37825 12023 37859
rect 13921 37825 13955 37859
rect 16129 37825 16163 37859
rect 17417 37825 17451 37859
rect 17684 37825 17718 37859
rect 23392 37825 23426 37859
rect 23489 37825 23523 37859
rect 23581 37825 23615 37859
rect 23764 37825 23798 37859
rect 23857 37825 23891 37859
rect 23949 37825 23983 37859
rect 24133 37825 24167 37859
rect 30389 37825 30423 37859
rect 30481 37825 30515 37859
rect 30665 37825 30699 37859
rect 32597 37825 32631 37859
rect 32689 37825 32723 37859
rect 32873 37825 32907 37859
rect 38485 37825 38519 37859
rect 38761 37825 38795 37859
rect 38853 37825 38887 37859
rect 39129 37825 39163 37859
rect 39221 37825 39255 37859
rect 40003 37825 40037 37859
rect 40141 37825 40175 37859
rect 40233 37825 40267 37859
rect 40417 37825 40451 37859
rect 41613 37825 41647 37859
rect 41889 37825 41923 37859
rect 41981 37825 42015 37859
rect 43913 37825 43947 37859
rect 4629 37757 4663 37791
rect 6561 37757 6595 37791
rect 6653 37757 6687 37791
rect 7205 37757 7239 37791
rect 9137 37757 9171 37791
rect 9229 37757 9263 37791
rect 10241 37757 10275 37791
rect 14197 37757 14231 37791
rect 16681 37757 16715 37791
rect 24317 37757 24351 37791
rect 25145 37757 25179 37791
rect 28181 37757 28215 37791
rect 37841 37757 37875 37791
rect 38577 37757 38611 37791
rect 42165 37757 42199 37791
rect 42441 37757 42475 37791
rect 43821 37757 43855 37791
rect 44465 37757 44499 37791
rect 2973 37689 3007 37723
rect 43177 37689 43211 37723
rect 6009 37621 6043 37655
rect 7113 37621 7147 37655
rect 8677 37621 8711 37655
rect 13737 37621 13771 37655
rect 25789 37621 25823 37655
rect 30021 37621 30055 37655
rect 30573 37621 30607 37655
rect 37289 37621 37323 37655
rect 38301 37621 38335 37655
rect 38761 37621 38795 37655
rect 39405 37621 39439 37655
rect 41705 37621 41739 37655
rect 43085 37621 43119 37655
rect 3893 37417 3927 37451
rect 5089 37417 5123 37451
rect 6929 37417 6963 37451
rect 7573 37417 7607 37451
rect 12449 37417 12483 37451
rect 17693 37417 17727 37451
rect 18705 37417 18739 37451
rect 28917 37417 28951 37451
rect 33241 37417 33275 37451
rect 38761 37417 38795 37451
rect 44189 37417 44223 37451
rect 2881 37281 2915 37315
rect 3065 37281 3099 37315
rect 4537 37281 4571 37315
rect 5825 37281 5859 37315
rect 5917 37281 5951 37315
rect 6745 37281 6779 37315
rect 18153 37281 18187 37315
rect 21465 37281 21499 37315
rect 25605 37281 25639 37315
rect 27077 37281 27111 37315
rect 32873 37281 32907 37315
rect 35541 37281 35575 37315
rect 35817 37281 35851 37315
rect 42717 37281 42751 37315
rect 1409 37213 1443 37247
rect 2145 37213 2179 37247
rect 4261 37213 4295 37247
rect 5273 37213 5307 37247
rect 7113 37213 7147 37247
rect 7757 37213 7791 37247
rect 12633 37213 12667 37247
rect 15025 37213 15059 37247
rect 17877 37213 17911 37247
rect 18245 37213 18279 37247
rect 19257 37213 19291 37247
rect 19533 37213 19567 37247
rect 23489 37213 23523 37247
rect 24409 37213 24443 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 29837 37213 29871 37247
rect 30021 37213 30055 37247
rect 32781 37213 32815 37247
rect 33057 37213 33091 37247
rect 38117 37213 38151 37247
rect 38485 37213 38519 37247
rect 39313 37213 39347 37247
rect 42441 37213 42475 37247
rect 5733 37145 5767 37179
rect 6193 37145 6227 37179
rect 19778 37145 19812 37179
rect 21710 37145 21744 37179
rect 27445 37145 27479 37179
rect 38301 37145 38335 37179
rect 38393 37145 38427 37179
rect 40601 37145 40635 37179
rect 1593 37077 1627 37111
rect 1961 37077 1995 37111
rect 2421 37077 2455 37111
rect 2789 37077 2823 37111
rect 4353 37077 4387 37111
rect 5365 37077 5399 37111
rect 14933 37077 14967 37111
rect 18337 37077 18371 37111
rect 19441 37077 19475 37111
rect 20913 37077 20947 37111
rect 22845 37077 22879 37111
rect 22937 37077 22971 37111
rect 25053 37077 25087 37111
rect 29929 37077 29963 37111
rect 37289 37077 37323 37111
rect 38669 37077 38703 37111
rect 41889 37077 41923 37111
rect 3341 36873 3375 36907
rect 12817 36873 12851 36907
rect 14105 36873 14139 36907
rect 17141 36873 17175 36907
rect 19533 36873 19567 36907
rect 20821 36873 20855 36907
rect 21281 36873 21315 36907
rect 23397 36873 23431 36907
rect 24593 36873 24627 36907
rect 26709 36873 26743 36907
rect 30849 36873 30883 36907
rect 31677 36873 31711 36907
rect 36001 36873 36035 36907
rect 37749 36873 37783 36907
rect 38301 36873 38335 36907
rect 44189 36873 44223 36907
rect 1777 36805 1811 36839
rect 6377 36805 6411 36839
rect 12449 36805 12483 36839
rect 12654 36805 12688 36839
rect 19993 36805 20027 36839
rect 27169 36805 27203 36839
rect 30481 36805 30515 36839
rect 31309 36805 31343 36839
rect 33149 36805 33183 36839
rect 34161 36805 34195 36839
rect 34253 36805 34287 36839
rect 35725 36805 35759 36839
rect 37289 36805 37323 36839
rect 39773 36805 39807 36839
rect 1501 36737 1535 36771
rect 10517 36737 10551 36771
rect 10701 36737 10735 36771
rect 10793 36737 10827 36771
rect 10885 36737 10919 36771
rect 12909 36737 12943 36771
rect 13093 36737 13127 36771
rect 13461 36737 13495 36771
rect 13645 36737 13679 36771
rect 13737 36737 13771 36771
rect 13829 36737 13863 36771
rect 14197 36737 14231 36771
rect 14381 36737 14415 36771
rect 17049 36737 17083 36771
rect 19901 36737 19935 36771
rect 20637 36737 20671 36771
rect 22017 36737 22051 36771
rect 22284 36737 22318 36771
rect 24772 36737 24806 36771
rect 24869 36737 24903 36771
rect 24961 36737 24995 36771
rect 25144 36737 25178 36771
rect 25237 36737 25271 36771
rect 25329 36737 25363 36771
rect 25513 36737 25547 36771
rect 26801 36737 26835 36771
rect 29193 36737 29227 36771
rect 29285 36737 29319 36771
rect 29377 36737 29411 36771
rect 29515 36737 29549 36771
rect 30665 36737 30699 36771
rect 30941 36737 30975 36771
rect 31033 36737 31067 36771
rect 31125 36737 31159 36771
rect 31401 36737 31435 36771
rect 31493 36737 31527 36771
rect 32597 36737 32631 36771
rect 33241 36737 33275 36771
rect 33977 36737 34011 36771
rect 34345 36737 34379 36771
rect 35449 36737 35483 36771
rect 35633 36737 35667 36771
rect 35817 36737 35851 36771
rect 36185 36737 36219 36771
rect 37565 36737 37599 36771
rect 37841 36737 37875 36771
rect 38025 36737 38059 36771
rect 40049 36737 40083 36771
rect 41245 36737 41279 36771
rect 41337 36737 41371 36771
rect 41613 36737 41647 36771
rect 41889 36737 41923 36771
rect 41981 36737 42015 36771
rect 42257 36737 42291 36771
rect 42441 36737 42475 36771
rect 3249 36669 3283 36703
rect 3893 36669 3927 36703
rect 14289 36669 14323 36703
rect 17325 36669 17359 36703
rect 20177 36669 20211 36703
rect 21373 36669 21407 36703
rect 21465 36669 21499 36703
rect 25697 36669 25731 36703
rect 29653 36669 29687 36703
rect 29745 36669 29779 36703
rect 30297 36669 30331 36703
rect 31677 36669 31711 36703
rect 32505 36669 32539 36703
rect 36461 36669 36495 36703
rect 37381 36669 37415 36703
rect 40969 36669 41003 36703
rect 41061 36669 41095 36703
rect 42717 36669 42751 36703
rect 13277 36601 13311 36635
rect 20913 36601 20947 36635
rect 31033 36601 31067 36635
rect 32965 36601 32999 36635
rect 36737 36601 36771 36635
rect 42165 36601 42199 36635
rect 7665 36533 7699 36567
rect 11161 36533 11195 36567
rect 12633 36533 12667 36567
rect 16681 36533 16715 36567
rect 28457 36533 28491 36567
rect 29009 36533 29043 36567
rect 34529 36533 34563 36567
rect 36553 36533 36587 36567
rect 37289 36533 37323 36567
rect 37933 36533 37967 36567
rect 40325 36533 40359 36567
rect 41521 36533 41555 36567
rect 41705 36533 41739 36567
rect 10517 36329 10551 36363
rect 12449 36329 12483 36363
rect 14197 36329 14231 36363
rect 16037 36329 16071 36363
rect 22293 36329 22327 36363
rect 23029 36329 23063 36363
rect 27708 36329 27742 36363
rect 30205 36329 30239 36363
rect 32505 36329 32539 36363
rect 40220 36329 40254 36363
rect 42809 36329 42843 36363
rect 13553 36261 13587 36295
rect 13829 36261 13863 36295
rect 22201 36261 22235 36295
rect 27261 36261 27295 36295
rect 29929 36261 29963 36295
rect 10701 36193 10735 36227
rect 10977 36193 11011 36227
rect 13645 36193 13679 36227
rect 15945 36193 15979 36227
rect 17509 36193 17543 36227
rect 17785 36193 17819 36227
rect 21649 36193 21683 36227
rect 22845 36193 22879 36227
rect 24961 36193 24995 36227
rect 27445 36193 27479 36227
rect 30757 36193 30791 36227
rect 31033 36193 31067 36227
rect 32597 36193 32631 36227
rect 33885 36193 33919 36227
rect 36185 36193 36219 36227
rect 36461 36193 36495 36227
rect 39221 36193 39255 36227
rect 39497 36193 39531 36227
rect 39957 36193 39991 36227
rect 42165 36193 42199 36227
rect 3801 36125 3835 36159
rect 5365 36125 5399 36159
rect 6285 36125 6319 36159
rect 9413 36125 9447 36159
rect 9597 36125 9631 36159
rect 9873 36125 9907 36159
rect 10425 36125 10459 36159
rect 10609 36125 10643 36159
rect 12633 36125 12667 36159
rect 12817 36125 12851 36159
rect 13369 36125 13403 36159
rect 13553 36125 13587 36159
rect 13921 36125 13955 36159
rect 18061 36125 18095 36159
rect 19257 36125 19291 36159
rect 19533 36125 19567 36159
rect 23213 36125 23247 36159
rect 24869 36125 24903 36159
rect 25789 36125 25823 36159
rect 26985 36125 27019 36159
rect 29561 36125 29595 36159
rect 29745 36125 29779 36159
rect 29837 36125 29871 36159
rect 30021 36125 30055 36159
rect 32781 36125 32815 36159
rect 32965 36125 32999 36159
rect 33083 36125 33117 36159
rect 33241 36125 33275 36159
rect 33333 36125 33367 36159
rect 6561 36057 6595 36091
rect 8953 36057 8987 36091
rect 9137 36057 9171 36091
rect 12725 36057 12759 36091
rect 15669 36057 15703 36091
rect 19778 36057 19812 36091
rect 21833 36057 21867 36091
rect 25237 36057 25271 36091
rect 32873 36057 32907 36091
rect 3893 35989 3927 36023
rect 5181 35989 5215 36023
rect 8033 35989 8067 36023
rect 9321 35989 9355 36023
rect 9505 35989 9539 36023
rect 9689 35989 9723 36023
rect 13645 35989 13679 36023
rect 17877 35989 17911 36023
rect 19441 35989 19475 36023
rect 20913 35989 20947 36023
rect 21741 35989 21775 36023
rect 24409 35989 24443 36023
rect 24777 35989 24811 36023
rect 29193 35989 29227 36023
rect 34713 35989 34747 36023
rect 37749 35989 37783 36023
rect 41705 35989 41739 36023
rect 4445 35785 4479 35819
rect 5457 35785 5491 35819
rect 5917 35785 5951 35819
rect 11253 35785 11287 35819
rect 13921 35785 13955 35819
rect 14197 35785 14231 35819
rect 20085 35785 20119 35819
rect 20453 35785 20487 35819
rect 20913 35785 20947 35819
rect 23857 35785 23891 35819
rect 25329 35785 25363 35819
rect 29929 35785 29963 35819
rect 31217 35785 31251 35819
rect 32689 35785 32723 35819
rect 33885 35785 33919 35819
rect 34345 35785 34379 35819
rect 34529 35785 34563 35819
rect 35725 35785 35759 35819
rect 37933 35785 37967 35819
rect 6469 35717 6503 35751
rect 6685 35717 6719 35751
rect 7941 35717 7975 35751
rect 14105 35717 14139 35751
rect 17693 35717 17727 35751
rect 20545 35717 20579 35751
rect 24194 35717 24228 35751
rect 32505 35717 32539 35751
rect 35449 35717 35483 35751
rect 3332 35649 3366 35683
rect 5089 35649 5123 35683
rect 5825 35649 5859 35683
rect 7113 35649 7147 35683
rect 7389 35649 7423 35683
rect 7573 35649 7607 35683
rect 8033 35649 8067 35683
rect 8953 35649 8987 35683
rect 11161 35649 11195 35683
rect 11345 35649 11379 35683
rect 11621 35649 11655 35683
rect 11713 35649 11747 35683
rect 13829 35649 13863 35683
rect 14749 35649 14783 35683
rect 16313 35649 16347 35683
rect 17417 35649 17451 35683
rect 21465 35649 21499 35683
rect 23673 35649 23707 35683
rect 27997 35649 28031 35683
rect 29469 35649 29503 35683
rect 30389 35649 30423 35683
rect 32413 35649 32447 35683
rect 32597 35649 32631 35683
rect 32873 35649 32907 35683
rect 33057 35649 33091 35683
rect 33517 35649 33551 35683
rect 33977 35649 34011 35683
rect 34161 35649 34195 35683
rect 35081 35649 35115 35683
rect 3065 35581 3099 35615
rect 6009 35581 6043 35615
rect 6929 35581 6963 35615
rect 7297 35581 7331 35615
rect 9229 35581 9263 35615
rect 20637 35581 20671 35615
rect 22385 35581 22419 35615
rect 23949 35581 23983 35615
rect 27721 35581 27755 35615
rect 29745 35581 29779 35615
rect 30297 35581 30331 35615
rect 33609 35581 33643 35615
rect 37381 35581 37415 35615
rect 41521 35581 41555 35615
rect 7757 35513 7791 35547
rect 14105 35513 14139 35547
rect 16497 35513 16531 35547
rect 29561 35513 29595 35547
rect 4537 35445 4571 35479
rect 6653 35445 6687 35479
rect 6837 35445 6871 35479
rect 10701 35445 10735 35479
rect 19165 35445 19199 35479
rect 21833 35445 21867 35479
rect 40969 35445 41003 35479
rect 3433 35241 3467 35275
rect 6837 35241 6871 35275
rect 9229 35241 9263 35275
rect 9413 35241 9447 35275
rect 17877 35241 17911 35275
rect 22017 35241 22051 35275
rect 24225 35241 24259 35275
rect 25893 35241 25927 35275
rect 30297 35241 30331 35275
rect 33793 35241 33827 35275
rect 3893 35173 3927 35207
rect 33241 35173 33275 35207
rect 4537 35105 4571 35139
rect 18337 35105 18371 35139
rect 18429 35105 18463 35139
rect 22477 35105 22511 35139
rect 22661 35105 22695 35139
rect 26157 35105 26191 35139
rect 28181 35105 28215 35139
rect 33701 35105 33735 35139
rect 40693 35105 40727 35139
rect 40969 35105 41003 35139
rect 42441 35105 42475 35139
rect 43085 35105 43119 35139
rect 1685 35037 1719 35071
rect 3617 35037 3651 35071
rect 4261 35037 4295 35071
rect 4721 35037 4755 35071
rect 7021 35037 7055 35071
rect 11713 35037 11747 35071
rect 18245 35037 18279 35071
rect 20453 35037 20487 35071
rect 23397 35037 23431 35071
rect 24041 35037 24075 35071
rect 29929 35037 29963 35071
rect 30113 35037 30147 35071
rect 33149 35037 33183 35071
rect 33333 35037 33367 35071
rect 33885 35037 33919 35071
rect 33977 35037 34011 35071
rect 37197 35037 37231 35071
rect 38669 35037 38703 35071
rect 40417 35037 40451 35071
rect 44833 35037 44867 35071
rect 1952 34969 1986 35003
rect 4997 34969 5031 35003
rect 9045 34969 9079 35003
rect 9261 34969 9295 35003
rect 22385 34969 22419 35003
rect 22845 34969 22879 35003
rect 27905 34969 27939 35003
rect 36921 34969 36955 35003
rect 3065 34901 3099 34935
rect 4353 34901 4387 34935
rect 6469 34901 6503 34935
rect 11805 34901 11839 34935
rect 19901 34901 19935 34935
rect 24409 34901 24443 34935
rect 26433 34901 26467 34935
rect 35449 34901 35483 34935
rect 38117 34901 38151 34935
rect 39865 34901 39899 34935
rect 42533 34901 42567 34935
rect 44649 34901 44683 34935
rect 2145 34697 2179 34731
rect 2697 34697 2731 34731
rect 3157 34697 3191 34731
rect 19901 34697 19935 34731
rect 20361 34697 20395 34731
rect 21649 34697 21683 34731
rect 23213 34697 23247 34731
rect 24317 34697 24351 34731
rect 24777 34697 24811 34731
rect 27813 34697 27847 34731
rect 33149 34697 33183 34731
rect 33701 34697 33735 34731
rect 36461 34697 36495 34731
rect 38209 34697 38243 34731
rect 41429 34697 41463 34731
rect 42717 34697 42751 34731
rect 22078 34629 22112 34663
rect 26433 34629 26467 34663
rect 36369 34629 36403 34663
rect 36737 34629 36771 34663
rect 43085 34629 43119 34663
rect 2329 34561 2363 34595
rect 3065 34561 3099 34595
rect 5365 34561 5399 34595
rect 7573 34561 7607 34595
rect 8585 34561 8619 34595
rect 10149 34561 10183 34595
rect 13093 34561 13127 34595
rect 13185 34561 13219 34595
rect 13553 34561 13587 34595
rect 13645 34561 13679 34595
rect 13829 34561 13863 34595
rect 13921 34561 13955 34595
rect 14105 34561 14139 34595
rect 17969 34561 18003 34595
rect 19809 34561 19843 34595
rect 20269 34561 20303 34595
rect 21465 34561 21499 34595
rect 23397 34561 23431 34595
rect 24685 34561 24719 34595
rect 26249 34561 26283 34595
rect 26525 34561 26559 34595
rect 26617 34561 26651 34595
rect 27169 34561 27203 34595
rect 32137 34561 32171 34595
rect 32321 34561 32355 34595
rect 33333 34561 33367 34595
rect 33517 34561 33551 34595
rect 33609 34561 33643 34595
rect 33793 34561 33827 34595
rect 35817 34561 35851 34595
rect 36645 34561 36679 34595
rect 36829 34561 36863 34595
rect 37013 34561 37047 34595
rect 38393 34561 38427 34595
rect 38485 34561 38519 34595
rect 38761 34561 38795 34595
rect 41613 34561 41647 34595
rect 41705 34561 41739 34595
rect 41981 34561 42015 34595
rect 42533 34561 42567 34595
rect 3341 34493 3375 34527
rect 8861 34493 8895 34527
rect 13461 34493 13495 34527
rect 17877 34493 17911 34527
rect 20453 34493 20487 34527
rect 21833 34493 21867 34527
rect 24869 34493 24903 34527
rect 32229 34493 32263 34527
rect 37473 34493 37507 34527
rect 38669 34493 38703 34527
rect 38853 34493 38887 34527
rect 39129 34493 39163 34527
rect 40601 34493 40635 34527
rect 41245 34493 41279 34527
rect 41889 34493 41923 34527
rect 42809 34493 42843 34527
rect 44833 34493 44867 34527
rect 13645 34425 13679 34459
rect 26801 34425 26835 34459
rect 4813 34357 4847 34391
rect 7389 34357 7423 34391
rect 8769 34357 8803 34391
rect 9505 34357 9539 34391
rect 9873 34357 9907 34391
rect 12909 34357 12943 34391
rect 14013 34357 14047 34391
rect 19625 34357 19659 34391
rect 23489 34357 23523 34391
rect 38117 34357 38151 34391
rect 40693 34357 40727 34391
rect 5181 34153 5215 34187
rect 8493 34153 8527 34187
rect 12633 34153 12667 34187
rect 13645 34153 13679 34187
rect 14657 34153 14691 34187
rect 14749 34153 14783 34187
rect 15761 34153 15795 34187
rect 17969 34153 18003 34187
rect 21005 34153 21039 34187
rect 33241 34153 33275 34187
rect 34069 34153 34103 34187
rect 37105 34153 37139 34187
rect 39405 34153 39439 34187
rect 42625 34153 42659 34187
rect 13369 34085 13403 34119
rect 14933 34085 14967 34119
rect 16313 34085 16347 34119
rect 18337 34085 18371 34119
rect 21373 34085 21407 34119
rect 8953 34017 8987 34051
rect 12449 34017 12483 34051
rect 14749 34017 14783 34051
rect 16957 34017 16991 34051
rect 17417 34017 17451 34051
rect 22109 34017 22143 34051
rect 22201 34017 22235 34051
rect 33057 34017 33091 34051
rect 37657 34017 37691 34051
rect 41981 34017 42015 34051
rect 42717 34017 42751 34051
rect 3249 33949 3283 33983
rect 3801 33949 3835 33983
rect 5733 33949 5767 33983
rect 7113 33949 7147 33983
rect 7380 33949 7414 33983
rect 10793 33949 10827 33983
rect 12725 33949 12759 33983
rect 12942 33949 12976 33983
rect 13461 33949 13495 33983
rect 13737 33949 13771 33983
rect 14565 33949 14599 33983
rect 15025 33949 15059 33983
rect 15209 33949 15243 33983
rect 15669 33949 15703 33983
rect 16037 33949 16071 33983
rect 16129 33949 16163 33983
rect 17049 33949 17083 33983
rect 17141 33949 17175 33983
rect 17325 33949 17359 33983
rect 18061 33949 18095 33983
rect 18337 33949 18371 33983
rect 19257 33949 19291 33983
rect 24593 33949 24627 33983
rect 29285 33949 29319 33983
rect 31217 33949 31251 33983
rect 32965 33949 32999 33983
rect 33333 33949 33367 33983
rect 33425 33949 33459 33983
rect 33609 33949 33643 33983
rect 33977 33949 34011 33983
rect 36001 33949 36035 33983
rect 36645 33949 36679 33983
rect 36829 33949 36863 33983
rect 36921 33949 36955 33983
rect 37197 33949 37231 33983
rect 41613 33949 41647 33983
rect 4046 33881 4080 33915
rect 9229 33881 9263 33915
rect 10885 33881 10919 33915
rect 11253 33881 11287 33915
rect 11437 33881 11471 33915
rect 15117 33881 15151 33915
rect 16405 33881 16439 33915
rect 16681 33881 16715 33915
rect 17509 33881 17543 33915
rect 17601 33881 17635 33915
rect 17785 33881 17819 33915
rect 19533 33881 19567 33915
rect 21189 33881 21223 33915
rect 35173 33881 35207 33915
rect 37933 33881 37967 33915
rect 39865 33881 39899 33915
rect 42165 33881 42199 33915
rect 42993 33881 43027 33915
rect 2697 33813 2731 33847
rect 6377 33813 6411 33847
rect 10701 33813 10735 33847
rect 11621 33813 11655 33847
rect 12173 33813 12207 33847
rect 12817 33813 12851 33847
rect 13001 33813 13035 33847
rect 16589 33813 16623 33847
rect 16773 33813 16807 33847
rect 18153 33813 18187 33847
rect 21649 33813 21683 33847
rect 22017 33813 22051 33847
rect 24777 33813 24811 33847
rect 27813 33813 27847 33847
rect 33057 33813 33091 33847
rect 33425 33813 33459 33847
rect 35449 33813 35483 33847
rect 36553 33813 36587 33847
rect 42257 33813 42291 33847
rect 44465 33813 44499 33847
rect 3341 33609 3375 33643
rect 3893 33609 3927 33643
rect 3985 33609 4019 33643
rect 4353 33609 4387 33643
rect 5089 33609 5123 33643
rect 5549 33609 5583 33643
rect 7573 33609 7607 33643
rect 8769 33609 8803 33643
rect 9137 33609 9171 33643
rect 9229 33609 9263 33643
rect 12173 33609 12207 33643
rect 14933 33609 14967 33643
rect 16681 33609 16715 33643
rect 17509 33609 17543 33643
rect 19901 33609 19935 33643
rect 24409 33609 24443 33643
rect 33793 33609 33827 33643
rect 36001 33609 36035 33643
rect 40325 33609 40359 33643
rect 42901 33609 42935 33643
rect 43453 33609 43487 33643
rect 3004 33541 3038 33575
rect 7941 33541 7975 33575
rect 10793 33541 10827 33575
rect 14105 33541 14139 33575
rect 14657 33541 14691 33575
rect 17325 33541 17359 33575
rect 24041 33541 24075 33575
rect 25881 33541 25915 33575
rect 3525 33473 3559 33507
rect 3709 33473 3743 33507
rect 5181 33473 5215 33507
rect 5825 33473 5859 33507
rect 7113 33473 7147 33507
rect 11069 33473 11103 33507
rect 11713 33473 11747 33507
rect 11851 33473 11885 33507
rect 12173 33473 12207 33507
rect 14013 33473 14047 33507
rect 14197 33473 14231 33507
rect 16405 33473 16439 33507
rect 16865 33473 16899 33507
rect 17693 33473 17727 33507
rect 17785 33473 17819 33507
rect 18061 33473 18095 33507
rect 18889 33473 18923 33507
rect 20177 33473 20211 33507
rect 21465 33473 21499 33507
rect 24225 33473 24259 33507
rect 26157 33473 26191 33507
rect 27629 33473 27663 33507
rect 27905 33473 27939 33507
rect 30021 33473 30055 33507
rect 33149 33473 33183 33507
rect 35541 33473 35575 33507
rect 35725 33473 35759 33507
rect 37289 33473 37323 33507
rect 39221 33473 39255 33507
rect 39497 33473 39531 33507
rect 39589 33473 39623 33507
rect 40233 33473 40267 33507
rect 40693 33473 40727 33507
rect 42073 33473 42107 33507
rect 42993 33473 43027 33507
rect 43637 33473 43671 33507
rect 3249 33405 3283 33439
rect 4445 33405 4479 33439
rect 4629 33405 4663 33439
rect 4997 33405 5031 33439
rect 6377 33405 6411 33439
rect 8033 33405 8067 33439
rect 8125 33405 8159 33439
rect 9413 33405 9447 33439
rect 10701 33405 10735 33439
rect 11161 33405 11195 33439
rect 15092 33405 15126 33439
rect 15209 33405 15243 33439
rect 15301 33405 15335 33439
rect 15577 33405 15611 33439
rect 17049 33405 17083 33439
rect 19257 33405 19291 33439
rect 28181 33405 28215 33439
rect 30297 33405 30331 33439
rect 31769 33405 31803 33439
rect 32689 33405 32723 33439
rect 35265 33405 35299 33439
rect 36461 33405 36495 33439
rect 37565 33405 37599 33439
rect 39313 33405 39347 33439
rect 40509 33405 40543 33439
rect 41245 33405 41279 33439
rect 42717 33405 42751 33439
rect 44373 33405 44407 33439
rect 7021 33337 7055 33371
rect 11345 33337 11379 33371
rect 14289 33337 14323 33371
rect 14841 33337 14875 33371
rect 17969 33337 18003 33371
rect 27813 33337 27847 33371
rect 33701 33337 33735 33371
rect 39773 33337 39807 33371
rect 43361 33337 43395 33371
rect 44097 33337 44131 33371
rect 1869 33269 1903 33303
rect 5641 33269 5675 33303
rect 7205 33269 7239 33303
rect 11989 33269 12023 33303
rect 14657 33269 14691 33303
rect 15853 33269 15887 33303
rect 16865 33269 16899 33303
rect 18797 33269 18831 33303
rect 20085 33269 20119 33303
rect 21281 33269 21315 33303
rect 29653 33269 29687 33303
rect 32137 33269 32171 33303
rect 37105 33269 37139 33303
rect 39037 33269 39071 33303
rect 39865 33269 39899 33303
rect 41521 33269 41555 33303
rect 43913 33269 43947 33303
rect 3617 33065 3651 33099
rect 5825 33065 5859 33099
rect 8125 33065 8159 33099
rect 11805 33065 11839 33099
rect 11989 33065 12023 33099
rect 14841 33065 14875 33099
rect 16773 33065 16807 33099
rect 17877 33065 17911 33099
rect 18429 33065 18463 33099
rect 24685 33065 24719 33099
rect 28181 33065 28215 33099
rect 30205 33065 30239 33099
rect 30573 33065 30607 33099
rect 31217 33065 31251 33099
rect 34345 33065 34379 33099
rect 35265 33065 35299 33099
rect 37105 33065 37139 33099
rect 41613 33065 41647 33099
rect 2053 32997 2087 33031
rect 13185 32997 13219 33031
rect 30113 32997 30147 33031
rect 31033 32997 31067 33031
rect 33057 32997 33091 33031
rect 37565 32997 37599 33031
rect 39681 32997 39715 33031
rect 2513 32929 2547 32963
rect 2697 32929 2731 32963
rect 3065 32929 3099 32963
rect 6745 32929 6779 32963
rect 9505 32929 9539 32963
rect 11161 32929 11195 32963
rect 11713 32929 11747 32963
rect 15117 32929 15151 32963
rect 15301 32929 15335 32963
rect 20729 32929 20763 32963
rect 25237 32929 25271 32963
rect 26341 32929 26375 32963
rect 28825 32929 28859 32963
rect 29653 32929 29687 32963
rect 30297 32929 30331 32963
rect 31861 32929 31895 32963
rect 32505 32929 32539 32963
rect 33145 32929 33179 32963
rect 38669 32929 38703 32963
rect 40141 32929 40175 32963
rect 1961 32861 1995 32895
rect 2421 32861 2455 32895
rect 3249 32861 3283 32895
rect 4445 32861 4479 32895
rect 6101 32861 6135 32895
rect 8953 32861 8987 32895
rect 10793 32861 10827 32895
rect 10977 32861 11011 32895
rect 11253 32861 11287 32895
rect 11437 32861 11471 32895
rect 11621 32861 11655 32895
rect 12909 32861 12943 32895
rect 13001 32861 13035 32895
rect 13277 32861 13311 32895
rect 15025 32861 15059 32895
rect 15209 32861 15243 32895
rect 15485 32861 15519 32895
rect 17325 32861 17359 32895
rect 17601 32861 17635 32895
rect 17693 32861 17727 32895
rect 18705 32861 18739 32895
rect 23857 32861 23891 32895
rect 25053 32861 25087 32895
rect 25145 32861 25179 32895
rect 26065 32861 26099 32895
rect 29745 32861 29779 32895
rect 30205 32861 30239 32895
rect 30941 32861 30975 32895
rect 31125 32861 31159 32895
rect 31401 32861 31435 32895
rect 31493 32861 31527 32895
rect 31585 32861 31619 32895
rect 32597 32861 32631 32895
rect 32781 32861 32815 32895
rect 32965 32861 32999 32895
rect 33241 32861 33275 32895
rect 33517 32861 33551 32895
rect 33793 32861 33827 32895
rect 34161 32861 34195 32895
rect 37013 32861 37047 32895
rect 37289 32861 37323 32895
rect 37381 32861 37415 32895
rect 37657 32861 37691 32895
rect 39497 32861 39531 32895
rect 39865 32861 39899 32895
rect 41797 32861 41831 32895
rect 4712 32793 4746 32827
rect 7012 32793 7046 32827
rect 17509 32793 17543 32827
rect 21005 32793 21039 32827
rect 24225 32793 24259 32827
rect 26617 32793 26651 32827
rect 28549 32793 28583 32827
rect 31723 32793 31757 32827
rect 33977 32793 34011 32827
rect 34069 32793 34103 32827
rect 36737 32793 36771 32827
rect 1777 32725 1811 32759
rect 3157 32725 3191 32759
rect 5917 32725 5951 32759
rect 11437 32725 11471 32759
rect 12725 32725 12759 32759
rect 18245 32725 18279 32759
rect 22477 32725 22511 32759
rect 26249 32725 26283 32759
rect 28089 32725 28123 32759
rect 28641 32725 28675 32759
rect 32137 32725 32171 32759
rect 38025 32725 38059 32759
rect 41889 32725 41923 32759
rect 2881 32521 2915 32555
rect 3801 32521 3835 32555
rect 6745 32521 6779 32555
rect 6837 32521 6871 32555
rect 7205 32521 7239 32555
rect 7849 32521 7883 32555
rect 15669 32521 15703 32555
rect 16405 32521 16439 32555
rect 21373 32521 21407 32555
rect 22845 32521 22879 32555
rect 26985 32521 27019 32555
rect 27353 32521 27387 32555
rect 29745 32521 29779 32555
rect 30941 32521 30975 32555
rect 32137 32521 32171 32555
rect 33241 32521 33275 32555
rect 40325 32521 40359 32555
rect 1768 32453 1802 32487
rect 3893 32453 3927 32487
rect 5641 32453 5675 32487
rect 13553 32453 13587 32487
rect 16773 32453 16807 32487
rect 17509 32453 17543 32487
rect 23213 32453 23247 32487
rect 31585 32453 31619 32487
rect 31769 32453 31803 32487
rect 31953 32453 31987 32487
rect 40693 32453 40727 32487
rect 3157 32385 3191 32419
rect 6193 32385 6227 32419
rect 7389 32385 7423 32419
rect 10241 32385 10275 32419
rect 10333 32385 10367 32419
rect 10701 32385 10735 32419
rect 10793 32385 10827 32419
rect 10977 32385 11011 32419
rect 12173 32385 12207 32419
rect 12449 32385 12483 32419
rect 12541 32385 12575 32419
rect 12725 32385 12759 32419
rect 13415 32385 13449 32419
rect 13645 32385 13679 32419
rect 13773 32385 13807 32419
rect 13921 32385 13955 32419
rect 15853 32385 15887 32419
rect 15945 32385 15979 32419
rect 16129 32385 16163 32419
rect 16313 32385 16347 32419
rect 16497 32385 16531 32419
rect 16957 32385 16991 32419
rect 17049 32385 17083 32419
rect 17325 32385 17359 32419
rect 17785 32385 17819 32419
rect 18153 32385 18187 32419
rect 18705 32385 18739 32419
rect 21281 32385 21315 32419
rect 22661 32385 22695 32419
rect 29285 32385 29319 32419
rect 29561 32385 29595 32419
rect 30849 32385 30883 32419
rect 32321 32385 32355 32419
rect 32505 32385 32539 32419
rect 32873 32385 32907 32419
rect 40141 32385 40175 32419
rect 44005 32385 44039 32419
rect 1501 32317 1535 32351
rect 6929 32317 6963 32351
rect 7941 32317 7975 32351
rect 8033 32317 8067 32351
rect 10609 32317 10643 32351
rect 12265 32317 12299 32351
rect 16037 32317 16071 32351
rect 17877 32317 17911 32351
rect 18245 32317 18279 32351
rect 21097 32317 21131 32351
rect 22937 32317 22971 32351
rect 25973 32317 26007 32351
rect 27445 32317 27479 32351
rect 27629 32317 27663 32351
rect 29377 32317 29411 32351
rect 32965 32317 32999 32351
rect 40417 32317 40451 32351
rect 6377 32249 6411 32283
rect 7481 32249 7515 32283
rect 10793 32249 10827 32283
rect 16773 32249 16807 32283
rect 18061 32249 18095 32283
rect 6009 32181 6043 32215
rect 10057 32181 10091 32215
rect 12725 32181 12759 32215
rect 13277 32181 13311 32215
rect 17141 32181 17175 32215
rect 17693 32181 17727 32215
rect 18613 32181 18647 32215
rect 20545 32181 20579 32215
rect 24685 32181 24719 32215
rect 26525 32181 26559 32215
rect 42165 32181 42199 32215
rect 43821 32181 43855 32215
rect 10333 31977 10367 32011
rect 10793 31977 10827 32011
rect 14197 31977 14231 32011
rect 14289 31977 14323 32011
rect 17325 31977 17359 32011
rect 20637 31977 20671 32011
rect 23489 31977 23523 32011
rect 28733 31977 28767 32011
rect 30113 31977 30147 32011
rect 32413 31977 32447 32011
rect 40877 31977 40911 32011
rect 7021 31909 7055 31943
rect 9321 31909 9355 31943
rect 9873 31909 9907 31943
rect 9965 31909 9999 31943
rect 22661 31909 22695 31943
rect 24777 31909 24811 31943
rect 26893 31909 26927 31943
rect 35817 31909 35851 31943
rect 36093 31909 36127 31943
rect 38485 31909 38519 31943
rect 42717 31909 42751 31943
rect 2881 31841 2915 31875
rect 3065 31841 3099 31875
rect 5457 31841 5491 31875
rect 6929 31841 6963 31875
rect 7573 31841 7607 31875
rect 9137 31841 9171 31875
rect 10425 31841 10459 31875
rect 13001 31841 13035 31875
rect 13369 31841 13403 31875
rect 14289 31841 14323 31875
rect 17785 31841 17819 31875
rect 21097 31841 21131 31875
rect 21189 31841 21223 31875
rect 23121 31841 23155 31875
rect 23213 31841 23247 31875
rect 24133 31841 24167 31875
rect 25421 31841 25455 31875
rect 26985 31841 27019 31875
rect 27261 31841 27295 31875
rect 29837 31841 29871 31875
rect 36553 31841 36587 31875
rect 36645 31841 36679 31875
rect 38945 31841 38979 31875
rect 39037 31841 39071 31875
rect 41429 31841 41463 31875
rect 43085 31841 43119 31875
rect 5181 31773 5215 31807
rect 7757 31773 7791 31807
rect 7849 31773 7883 31807
rect 9229 31773 9263 31807
rect 9597 31773 9631 31807
rect 9781 31773 9815 31807
rect 10057 31773 10091 31807
rect 10609 31773 10643 31807
rect 12909 31773 12943 31807
rect 13277 31773 13311 31807
rect 13921 31773 13955 31807
rect 14105 31773 14139 31807
rect 14473 31773 14507 31807
rect 17693 31773 17727 31807
rect 20361 31773 20395 31807
rect 21005 31773 21039 31807
rect 22201 31773 22235 31807
rect 22385 31773 22419 31807
rect 23949 31773 23983 31807
rect 24501 31773 24535 31807
rect 25237 31773 25271 31807
rect 26249 31773 26283 31807
rect 26525 31773 26559 31807
rect 26709 31773 26743 31807
rect 28825 31773 28859 31807
rect 29193 31773 29227 31807
rect 29745 31773 29779 31807
rect 32321 31773 32355 31807
rect 32505 31773 32539 31807
rect 35265 31773 35299 31807
rect 36001 31773 36035 31807
rect 38393 31773 38427 31807
rect 41245 31773 41279 31807
rect 41337 31773 41371 31807
rect 42533 31773 42567 31807
rect 42809 31773 42843 31807
rect 9321 31705 9355 31739
rect 10333 31705 10367 31739
rect 13829 31705 13863 31739
rect 23857 31705 23891 31739
rect 25145 31705 25179 31739
rect 25605 31705 25639 31739
rect 2421 31637 2455 31671
rect 2789 31637 2823 31671
rect 9505 31637 9539 31671
rect 10241 31637 10275 31671
rect 13553 31637 13587 31671
rect 20177 31637 20211 31671
rect 22017 31637 22051 31671
rect 22569 31637 22603 31671
rect 23029 31637 23063 31671
rect 24685 31637 24719 31671
rect 26341 31637 26375 31671
rect 34713 31637 34747 31671
rect 36461 31637 36495 31671
rect 38209 31637 38243 31671
rect 38853 31637 38887 31671
rect 44557 31637 44591 31671
rect 9229 31433 9263 31467
rect 9965 31433 9999 31467
rect 10517 31433 10551 31467
rect 18245 31433 18279 31467
rect 21281 31433 21315 31467
rect 21557 31433 21591 31467
rect 23673 31433 23707 31467
rect 24133 31433 24167 31467
rect 25973 31433 26007 31467
rect 27169 31433 27203 31467
rect 27537 31433 27571 31467
rect 29837 31433 29871 31467
rect 32321 31433 32355 31467
rect 32873 31433 32907 31467
rect 34069 31433 34103 31467
rect 39497 31433 39531 31467
rect 42625 31433 42659 31467
rect 43085 31433 43119 31467
rect 8861 31365 8895 31399
rect 9597 31365 9631 31399
rect 10057 31365 10091 31399
rect 10701 31365 10735 31399
rect 12449 31365 12483 31399
rect 15117 31365 15151 31399
rect 15209 31365 15243 31399
rect 15669 31365 15703 31399
rect 19809 31365 19843 31399
rect 22109 31365 22143 31399
rect 24768 31365 24802 31399
rect 33793 31365 33827 31399
rect 34437 31365 34471 31399
rect 38025 31365 38059 31399
rect 2145 31297 2179 31331
rect 7941 31297 7975 31331
rect 8401 31297 8435 31331
rect 8585 31297 8619 31331
rect 8677 31297 8711 31331
rect 8953 31297 8987 31331
rect 9045 31297 9079 31331
rect 9505 31297 9539 31331
rect 9781 31297 9815 31331
rect 10333 31297 10367 31331
rect 10609 31297 10643 31331
rect 10793 31297 10827 31331
rect 12173 31297 12207 31331
rect 12321 31297 12355 31331
rect 12541 31297 12575 31331
rect 12638 31297 12672 31331
rect 14749 31297 14783 31331
rect 14841 31297 14875 31331
rect 14934 31297 14968 31331
rect 15347 31297 15381 31331
rect 15761 31297 15795 31331
rect 18337 31297 18371 31331
rect 21649 31297 21683 31331
rect 24041 31297 24075 31331
rect 26341 31297 26375 31331
rect 29653 31297 29687 31331
rect 29837 31297 29871 31331
rect 32505 31297 32539 31331
rect 32689 31297 32723 31331
rect 32781 31297 32815 31331
rect 32965 31297 32999 31331
rect 33517 31297 33551 31331
rect 33701 31297 33735 31331
rect 33885 31297 33919 31331
rect 37749 31297 37783 31331
rect 42993 31297 43027 31331
rect 43637 31297 43671 31331
rect 43913 31297 43947 31331
rect 2513 31229 2547 31263
rect 2789 31229 2823 31263
rect 7849 31229 7883 31263
rect 10149 31229 10183 31263
rect 19533 31229 19567 31263
rect 21833 31229 21867 31263
rect 23581 31229 23615 31263
rect 24225 31229 24259 31263
rect 24501 31229 24535 31263
rect 26433 31229 26467 31263
rect 26525 31229 26559 31263
rect 27629 31229 27663 31263
rect 27721 31229 27755 31263
rect 34161 31229 34195 31263
rect 43177 31229 43211 31263
rect 25881 31161 25915 31195
rect 35909 31161 35943 31195
rect 43729 31161 43763 31195
rect 43821 31161 43855 31195
rect 1961 31093 1995 31127
rect 4261 31093 4295 31127
rect 8309 31093 8343 31127
rect 8401 31093 8435 31127
rect 10333 31093 10367 31127
rect 12817 31093 12851 31127
rect 13461 31093 13495 31127
rect 15485 31093 15519 31127
rect 43453 31093 43487 31127
rect 3341 30889 3375 30923
rect 9413 30889 9447 30923
rect 12633 30889 12667 30923
rect 13369 30889 13403 30923
rect 14243 30889 14277 30923
rect 14381 30889 14415 30923
rect 18429 30889 18463 30923
rect 22293 30889 22327 30923
rect 26801 30889 26835 30923
rect 30021 30889 30055 30923
rect 33517 30889 33551 30923
rect 33885 30889 33919 30923
rect 3249 30821 3283 30855
rect 3801 30821 3835 30855
rect 13829 30821 13863 30855
rect 16037 30821 16071 30855
rect 26065 30821 26099 30855
rect 1501 30753 1535 30787
rect 1777 30753 1811 30787
rect 4445 30753 4479 30787
rect 10057 30753 10091 30787
rect 12081 30753 12115 30787
rect 12817 30753 12851 30787
rect 13185 30753 13219 30787
rect 14473 30753 14507 30787
rect 14565 30753 14599 30787
rect 16681 30753 16715 30787
rect 16957 30753 16991 30787
rect 22845 30753 22879 30787
rect 26157 30753 26191 30787
rect 27813 30753 27847 30787
rect 29837 30753 29871 30787
rect 33333 30753 33367 30787
rect 35909 30753 35943 30787
rect 37657 30753 37691 30787
rect 40325 30753 40359 30787
rect 42809 30753 42843 30787
rect 43269 30753 43303 30787
rect 3525 30685 3559 30719
rect 4629 30685 4663 30719
rect 5181 30685 5215 30719
rect 8959 30685 8993 30719
rect 9137 30685 9171 30719
rect 9597 30685 9631 30719
rect 9689 30685 9723 30719
rect 10149 30685 10183 30719
rect 10241 30685 10275 30719
rect 10333 30685 10367 30719
rect 10885 30685 10919 30719
rect 11299 30685 11333 30719
rect 11437 30685 11471 30719
rect 11657 30685 11691 30719
rect 11805 30685 11839 30719
rect 12173 30684 12207 30718
rect 12449 30685 12483 30719
rect 12541 30685 12575 30719
rect 12909 30685 12943 30719
rect 13369 30685 13403 30719
rect 13553 30685 13587 30719
rect 13645 30685 13679 30719
rect 15853 30685 15887 30719
rect 16313 30685 16347 30719
rect 16589 30685 16623 30719
rect 18889 30685 18923 30719
rect 21005 30685 21039 30719
rect 24685 30685 24719 30719
rect 24952 30685 24986 30719
rect 27169 30685 27203 30719
rect 29745 30685 29779 30719
rect 33241 30685 33275 30719
rect 33977 30685 34011 30719
rect 35633 30685 35667 30719
rect 40233 30685 40267 30719
rect 43177 30685 43211 30719
rect 4261 30617 4295 30651
rect 4721 30617 4755 30651
rect 9965 30617 9999 30651
rect 10977 30617 11011 30651
rect 11529 30617 11563 30651
rect 13277 30617 13311 30651
rect 14105 30617 14139 30651
rect 23090 30617 23124 30651
rect 4169 30549 4203 30583
rect 4997 30549 5031 30583
rect 9045 30549 9079 30583
rect 11161 30549 11195 30583
rect 11897 30549 11931 30583
rect 16129 30549 16163 30583
rect 16497 30549 16531 30583
rect 19073 30549 19107 30583
rect 24225 30549 24259 30583
rect 27353 30549 27387 30583
rect 28457 30549 28491 30583
rect 40601 30549 40635 30583
rect 5917 30345 5951 30379
rect 16129 30345 16163 30379
rect 23673 30345 23707 30379
rect 32321 30345 32355 30379
rect 33701 30345 33735 30379
rect 40693 30345 40727 30379
rect 4445 30277 4479 30311
rect 6561 30277 6595 30311
rect 6929 30277 6963 30311
rect 12357 30277 12391 30311
rect 16297 30277 16331 30311
rect 16497 30277 16531 30311
rect 16773 30277 16807 30311
rect 16957 30277 16991 30311
rect 19533 30277 19567 30311
rect 22201 30277 22235 30311
rect 27261 30277 27295 30311
rect 32505 30277 32539 30311
rect 33517 30277 33551 30311
rect 38025 30277 38059 30311
rect 39681 30277 39715 30311
rect 43637 30277 43671 30311
rect 4169 30209 4203 30243
rect 6745 30209 6779 30243
rect 6837 30209 6871 30243
rect 7021 30209 7055 30243
rect 12633 30209 12667 30243
rect 16681 30209 16715 30243
rect 24225 30209 24259 30243
rect 26617 30209 26651 30243
rect 29469 30209 29503 30243
rect 29745 30209 29779 30243
rect 32229 30209 32263 30243
rect 32689 30209 32723 30243
rect 33001 30209 33035 30243
rect 33149 30209 33183 30243
rect 33333 30209 33367 30243
rect 33609 30209 33643 30243
rect 33977 30209 34011 30243
rect 37289 30209 37323 30243
rect 37933 30209 37967 30243
rect 38577 30209 38611 30243
rect 39313 30209 39347 30243
rect 39497 30209 39531 30243
rect 39589 30209 39623 30243
rect 39865 30209 39899 30243
rect 39957 30209 39991 30243
rect 40969 30209 41003 30243
rect 43361 30209 43395 30243
rect 12541 30141 12575 30175
rect 19257 30141 19291 30175
rect 21005 30141 21039 30175
rect 22845 30141 22879 30175
rect 26985 30141 27019 30175
rect 28733 30141 28767 30175
rect 33701 30141 33735 30175
rect 38117 30141 38151 30175
rect 39221 30141 39255 30175
rect 40693 30141 40727 30175
rect 43453 30141 43487 30175
rect 12817 30073 12851 30107
rect 16681 30073 16715 30107
rect 29561 30073 29595 30107
rect 32781 30073 32815 30107
rect 32873 30073 32907 30107
rect 37565 30073 37599 30107
rect 6377 30005 6411 30039
rect 12633 30005 12667 30039
rect 16313 30005 16347 30039
rect 26801 30005 26835 30039
rect 29929 30005 29963 30039
rect 33885 30005 33919 30039
rect 37473 30005 37507 30039
rect 39313 30005 39347 30039
rect 39681 30005 39715 30039
rect 40877 30005 40911 30039
rect 43177 30005 43211 30039
rect 43361 30005 43395 30039
rect 5181 29801 5215 29835
rect 5365 29801 5399 29835
rect 11253 29801 11287 29835
rect 14197 29801 14231 29835
rect 19717 29801 19751 29835
rect 27077 29801 27111 29835
rect 27169 29801 27203 29835
rect 28917 29801 28951 29835
rect 29377 29801 29411 29835
rect 30205 29801 30239 29835
rect 32413 29801 32447 29835
rect 32965 29801 32999 29835
rect 33517 29801 33551 29835
rect 40141 29801 40175 29835
rect 40509 29801 40543 29835
rect 42993 29801 43027 29835
rect 43637 29801 43671 29835
rect 31769 29733 31803 29767
rect 41797 29733 41831 29767
rect 6377 29665 6411 29699
rect 20361 29665 20395 29699
rect 27721 29665 27755 29699
rect 29009 29665 29043 29699
rect 29837 29665 29871 29699
rect 30573 29665 30607 29699
rect 35357 29665 35391 29699
rect 39497 29665 39531 29699
rect 40417 29665 40451 29699
rect 40969 29665 41003 29699
rect 41153 29665 41187 29699
rect 41429 29665 41463 29699
rect 41521 29665 41555 29699
rect 43821 29665 43855 29699
rect 5917 29597 5951 29631
rect 6009 29597 6043 29631
rect 6101 29597 6135 29631
rect 6285 29597 6319 29631
rect 10057 29597 10091 29631
rect 11161 29597 11195 29631
rect 14289 29597 14323 29631
rect 15301 29597 15335 29631
rect 15485 29597 15519 29631
rect 15761 29597 15795 29631
rect 20085 29597 20119 29631
rect 22293 29597 22327 29631
rect 22385 29597 22419 29631
rect 22937 29597 22971 29631
rect 24961 29597 24995 29631
rect 26065 29597 26099 29631
rect 26433 29597 26467 29631
rect 27537 29597 27571 29631
rect 29193 29597 29227 29631
rect 29745 29597 29779 29631
rect 30389 29597 30423 29631
rect 30481 29597 30515 29631
rect 30665 29597 30699 29631
rect 31769 29597 31803 29631
rect 31953 29597 31987 29631
rect 32137 29597 32171 29631
rect 32229 29597 32263 29631
rect 32781 29597 32815 29631
rect 33609 29597 33643 29631
rect 33793 29597 33827 29631
rect 35173 29597 35207 29631
rect 39221 29597 39255 29631
rect 39405 29597 39439 29631
rect 40509 29597 40543 29631
rect 40785 29597 40819 29631
rect 41061 29597 41095 29631
rect 41337 29597 41371 29631
rect 41613 29597 41647 29631
rect 41797 29597 41831 29631
rect 41981 29597 42015 29631
rect 42073 29597 42107 29631
rect 42717 29597 42751 29631
rect 42809 29597 42843 29631
rect 43545 29597 43579 29631
rect 5349 29529 5383 29563
rect 5549 29529 5583 29563
rect 5641 29529 5675 29563
rect 6653 29529 6687 29563
rect 15669 29529 15703 29563
rect 24409 29529 24443 29563
rect 27629 29529 27663 29563
rect 28917 29529 28951 29563
rect 32597 29529 32631 29563
rect 33149 29529 33183 29563
rect 33333 29529 33367 29563
rect 35081 29529 35115 29563
rect 35633 29529 35667 29563
rect 38945 29529 38979 29563
rect 42993 29529 43027 29563
rect 8125 29461 8159 29495
rect 10149 29461 10183 29495
rect 15393 29461 15427 29495
rect 20177 29461 20211 29495
rect 22109 29461 22143 29495
rect 25513 29461 25547 29495
rect 30113 29461 30147 29495
rect 33793 29461 33827 29495
rect 37105 29461 37139 29495
rect 37473 29461 37507 29495
rect 39037 29461 39071 29495
rect 40601 29461 40635 29495
rect 43821 29461 43855 29495
rect 6377 29257 6411 29291
rect 11345 29257 11379 29291
rect 12817 29257 12851 29291
rect 14565 29257 14599 29291
rect 15511 29257 15545 29291
rect 16037 29257 16071 29291
rect 16497 29257 16531 29291
rect 18429 29257 18463 29291
rect 23213 29257 23247 29291
rect 24869 29257 24903 29291
rect 32229 29257 32263 29291
rect 33425 29257 33459 29291
rect 35449 29257 35483 29291
rect 39037 29257 39071 29291
rect 39313 29257 39347 29291
rect 39865 29257 39899 29291
rect 40778 29257 40812 29291
rect 41061 29257 41095 29291
rect 10977 29189 11011 29223
rect 11069 29189 11103 29223
rect 11805 29189 11839 29223
rect 12449 29189 12483 29223
rect 14933 29189 14967 29223
rect 15301 29189 15335 29223
rect 16957 29189 16991 29223
rect 22089 29189 22123 29223
rect 24961 29189 24995 29223
rect 27261 29189 27295 29223
rect 32781 29189 32815 29223
rect 32965 29189 32999 29223
rect 35081 29189 35115 29223
rect 35173 29189 35207 29223
rect 35541 29189 35575 29223
rect 37565 29189 37599 29223
rect 40693 29189 40727 29223
rect 41429 29189 41463 29223
rect 5733 29121 5767 29155
rect 5917 29121 5951 29155
rect 6377 29121 6411 29155
rect 6561 29121 6595 29155
rect 10701 29121 10735 29155
rect 10794 29121 10828 29155
rect 11207 29121 11241 29155
rect 11713 29121 11747 29155
rect 12173 29121 12207 29155
rect 12266 29121 12300 29155
rect 12541 29121 12575 29155
rect 12679 29121 12713 29155
rect 14744 29121 14778 29155
rect 14841 29121 14875 29155
rect 15061 29121 15095 29155
rect 15209 29121 15243 29155
rect 15761 29121 15795 29155
rect 16037 29121 16071 29155
rect 16221 29121 16255 29155
rect 16313 29121 16347 29155
rect 18705 29121 18739 29155
rect 18889 29121 18923 29155
rect 18981 29121 19015 29155
rect 20637 29121 20671 29155
rect 23489 29121 23523 29155
rect 23756 29121 23790 29155
rect 29929 29121 29963 29155
rect 30389 29121 30423 29155
rect 30573 29121 30607 29155
rect 32321 29121 32355 29155
rect 33241 29121 33275 29155
rect 33425 29121 33459 29155
rect 34897 29121 34931 29155
rect 35265 29121 35299 29155
rect 36185 29121 36219 29155
rect 39129 29121 39163 29155
rect 39497 29121 39531 29155
rect 39773 29121 39807 29155
rect 40049 29121 40083 29155
rect 40601 29121 40635 29155
rect 40877 29121 40911 29155
rect 41153 29121 41187 29155
rect 41705 29121 41739 29155
rect 42073 29121 42107 29155
rect 42257 29121 42291 29155
rect 42809 29121 42843 29155
rect 42993 29121 43027 29155
rect 43361 29121 43395 29155
rect 43729 29121 43763 29155
rect 44649 29121 44683 29155
rect 16681 29053 16715 29087
rect 21833 29053 21867 29087
rect 26985 29053 27019 29087
rect 30021 29053 30055 29087
rect 30481 29053 30515 29087
rect 37289 29053 37323 29087
rect 40141 29053 40175 29087
rect 40233 29053 40267 29087
rect 40325 29053 40359 29087
rect 41245 29053 41279 29087
rect 41613 29053 41647 29087
rect 42533 29053 42567 29087
rect 43269 29053 43303 29087
rect 43821 29053 43855 29087
rect 43913 29053 43947 29087
rect 44005 29053 44039 29087
rect 44557 29053 44591 29087
rect 5825 28985 5859 29019
rect 15853 28985 15887 29019
rect 19165 28985 19199 29019
rect 26249 28985 26283 29019
rect 28733 28985 28767 29019
rect 30297 28985 30331 29019
rect 42625 28985 42659 29019
rect 44281 28985 44315 29019
rect 15485 28917 15519 28951
rect 15669 28917 15703 28951
rect 18521 28917 18555 28951
rect 20453 28917 20487 28951
rect 33149 28917 33183 28951
rect 39589 28917 39623 28951
rect 44189 28917 44223 28951
rect 6561 28713 6595 28747
rect 8493 28713 8527 28747
rect 9137 28713 9171 28747
rect 10517 28713 10551 28747
rect 11253 28713 11287 28747
rect 12909 28713 12943 28747
rect 13737 28713 13771 28747
rect 15301 28713 15335 28747
rect 18153 28713 18187 28747
rect 21373 28713 21407 28747
rect 22477 28713 22511 28747
rect 26341 28713 26375 28747
rect 26709 28713 26743 28747
rect 35081 28713 35115 28747
rect 43361 28713 43395 28747
rect 18337 28645 18371 28679
rect 24225 28645 24259 28679
rect 39405 28645 39439 28679
rect 44189 28645 44223 28679
rect 5273 28577 5307 28611
rect 8217 28577 8251 28611
rect 10057 28577 10091 28611
rect 13461 28577 13495 28611
rect 15761 28577 15795 28611
rect 18429 28577 18463 28611
rect 21281 28577 21315 28611
rect 22017 28577 22051 28611
rect 23121 28577 23155 28611
rect 23581 28577 23615 28611
rect 27353 28577 27387 28611
rect 32597 28577 32631 28611
rect 33333 28577 33367 28611
rect 34069 28577 34103 28611
rect 35265 28577 35299 28611
rect 38761 28577 38795 28611
rect 40509 28577 40543 28611
rect 5457 28509 5491 28543
rect 6101 28509 6135 28543
rect 6193 28509 6227 28543
rect 6561 28509 6595 28543
rect 6745 28509 6779 28543
rect 7941 28509 7975 28543
rect 8033 28509 8067 28543
rect 9413 28509 9447 28543
rect 10149 28509 10183 28543
rect 11161 28509 11195 28543
rect 13093 28509 13127 28543
rect 13185 28509 13219 28543
rect 13829 28509 13863 28543
rect 15669 28509 15703 28543
rect 17417 28509 17451 28543
rect 17601 28509 17635 28543
rect 17693 28509 17727 28543
rect 17877 28509 17911 28543
rect 18981 28509 19015 28543
rect 19257 28509 19291 28543
rect 21741 28509 21775 28543
rect 22845 28509 22879 28543
rect 23765 28509 23799 28543
rect 24961 28509 24995 28543
rect 27077 28509 27111 28543
rect 32689 28509 32723 28543
rect 33609 28509 33643 28543
rect 33793 28509 33827 28543
rect 34161 28509 34195 28543
rect 34345 28509 34379 28543
rect 35357 28509 35391 28543
rect 36001 28509 36035 28543
rect 36185 28509 36219 28543
rect 38945 28509 38979 28543
rect 39405 28509 39439 28543
rect 39865 28509 39899 28543
rect 40049 28509 40083 28543
rect 40417 28509 40451 28543
rect 40877 28509 40911 28543
rect 42073 28509 42107 28543
rect 43913 28509 43947 28543
rect 44189 28509 44223 28543
rect 5733 28441 5767 28475
rect 5917 28441 5951 28475
rect 8217 28441 8251 28475
rect 8677 28441 8711 28475
rect 8953 28441 8987 28475
rect 9169 28441 9203 28475
rect 9505 28441 9539 28475
rect 13553 28441 13587 28475
rect 17969 28441 18003 28475
rect 19533 28441 19567 28475
rect 21833 28441 21867 28475
rect 22937 28441 22971 28475
rect 23857 28441 23891 28475
rect 25228 28441 25262 28475
rect 27169 28441 27203 28475
rect 32321 28441 32355 28475
rect 33425 28441 33459 28475
rect 33701 28441 33735 28475
rect 33911 28441 33945 28475
rect 36093 28441 36127 28475
rect 40693 28441 40727 28475
rect 5641 28373 5675 28407
rect 6377 28373 6411 28407
rect 8309 28373 8343 28407
rect 8477 28373 8511 28407
rect 9321 28373 9355 28407
rect 17601 28373 17635 28407
rect 17877 28373 17911 28407
rect 18169 28373 18203 28407
rect 30849 28373 30883 28407
rect 34161 28373 34195 28407
rect 44005 28373 44039 28407
rect 3801 28169 3835 28203
rect 7665 28169 7699 28203
rect 14473 28169 14507 28203
rect 14636 28169 14670 28203
rect 21833 28169 21867 28203
rect 23673 28169 23707 28203
rect 25421 28169 25455 28203
rect 25697 28169 25731 28203
rect 38945 28169 38979 28203
rect 39773 28169 39807 28203
rect 44281 28169 44315 28203
rect 5641 28101 5675 28135
rect 6009 28101 6043 28135
rect 12909 28101 12943 28135
rect 14815 28101 14849 28135
rect 24961 28101 24995 28135
rect 34805 28101 34839 28135
rect 35725 28101 35759 28135
rect 1409 28033 1443 28067
rect 5549 28033 5583 28067
rect 5825 28033 5859 28067
rect 6377 28033 6411 28067
rect 6561 28033 6595 28067
rect 6653 28033 6687 28067
rect 6745 28033 6779 28067
rect 12541 28033 12575 28067
rect 12633 28033 12667 28067
rect 12817 28033 12851 28067
rect 13185 28033 13219 28067
rect 13645 28033 13679 28067
rect 14197 28033 14231 28067
rect 15209 28033 15243 28067
rect 18245 28033 18279 28067
rect 19993 28033 20027 28067
rect 20260 28033 20294 28067
rect 23857 28033 23891 28067
rect 25605 28033 25639 28067
rect 26341 28033 26375 28067
rect 34989 28033 35023 28067
rect 35081 28033 35115 28067
rect 35265 28033 35299 28067
rect 35357 28033 35391 28067
rect 35633 28033 35667 28067
rect 35817 28033 35851 28067
rect 35909 28033 35943 28067
rect 38853 28033 38887 28067
rect 39037 28033 39071 28067
rect 39497 28033 39531 28067
rect 42441 28033 42475 28067
rect 42625 28033 42659 28067
rect 42993 28033 43027 28067
rect 43453 28033 43487 28067
rect 43729 28033 43763 28067
rect 43913 28033 43947 28067
rect 44005 28033 44039 28067
rect 44097 28033 44131 28067
rect 44373 28033 44407 28067
rect 5273 27965 5307 27999
rect 9137 27965 9171 27999
rect 9413 27965 9447 27999
rect 9597 27965 9631 27999
rect 11069 27965 11103 27999
rect 11345 27965 11379 27999
rect 12909 27965 12943 27999
rect 14381 27965 14415 27999
rect 14933 27965 14967 27999
rect 15117 27965 15151 27999
rect 17877 27965 17911 27999
rect 19717 27965 19751 27999
rect 22385 27965 22419 27999
rect 24685 27965 24719 27999
rect 24869 27965 24903 27999
rect 36737 27965 36771 27999
rect 42901 27965 42935 27999
rect 12449 27897 12483 27931
rect 13093 27897 13127 27931
rect 21373 27897 21407 27931
rect 25329 27897 25363 27931
rect 43361 27897 43395 27931
rect 1593 27829 1627 27863
rect 7021 27829 7055 27863
rect 12817 27829 12851 27863
rect 13553 27829 13587 27863
rect 14013 27829 14047 27863
rect 14657 27829 14691 27863
rect 15025 27829 15059 27863
rect 34805 27829 34839 27863
rect 35265 27829 35299 27863
rect 36001 27829 36035 27863
rect 36185 27829 36219 27863
rect 43545 27829 43579 27863
rect 44097 27829 44131 27863
rect 4813 27625 4847 27659
rect 5457 27625 5491 27659
rect 5825 27625 5859 27659
rect 9045 27625 9079 27659
rect 12344 27625 12378 27659
rect 13829 27625 13863 27659
rect 16037 27625 16071 27659
rect 26617 27625 26651 27659
rect 26966 27625 27000 27659
rect 36737 27625 36771 27659
rect 38221 27625 38255 27659
rect 39405 27625 39439 27659
rect 5273 27557 5307 27591
rect 10241 27557 10275 27591
rect 22017 27557 22051 27591
rect 23489 27557 23523 27591
rect 34437 27557 34471 27591
rect 34713 27557 34747 27591
rect 39313 27557 39347 27591
rect 12081 27489 12115 27523
rect 14289 27489 14323 27523
rect 22109 27489 22143 27523
rect 24961 27489 24995 27523
rect 26709 27489 26743 27523
rect 35081 27489 35115 27523
rect 38485 27489 38519 27523
rect 4629 27421 4663 27455
rect 5733 27421 5767 27455
rect 7021 27421 7055 27455
rect 9229 27421 9263 27455
rect 9413 27421 9447 27455
rect 10057 27421 10091 27455
rect 19901 27421 19935 27455
rect 21833 27421 21867 27455
rect 24041 27421 24075 27455
rect 24777 27421 24811 27455
rect 26433 27421 26467 27455
rect 34345 27421 34379 27455
rect 34529 27421 34563 27455
rect 35265 27421 35299 27455
rect 35633 27421 35667 27455
rect 36001 27421 36035 27455
rect 36369 27421 36403 27455
rect 39865 27421 39899 27455
rect 40325 27421 40359 27455
rect 40509 27421 40543 27455
rect 5641 27353 5675 27387
rect 14565 27353 14599 27387
rect 20177 27353 20211 27387
rect 22354 27353 22388 27387
rect 23673 27353 23707 27387
rect 38945 27353 38979 27387
rect 5441 27285 5475 27319
rect 8309 27285 8343 27319
rect 24409 27285 24443 27319
rect 24869 27285 24903 27319
rect 28457 27285 28491 27319
rect 8401 27081 8435 27115
rect 8953 27081 8987 27115
rect 13461 27081 13495 27115
rect 14933 27081 14967 27115
rect 22385 27081 22419 27115
rect 22753 27081 22787 27115
rect 25789 27081 25823 27115
rect 26985 27081 27019 27115
rect 27353 27081 27387 27115
rect 29009 27081 29043 27115
rect 35265 27081 35299 27115
rect 35541 27081 35575 27115
rect 6653 27013 6687 27047
rect 14749 27013 14783 27047
rect 36027 27013 36061 27047
rect 42625 27013 42659 27047
rect 43729 27013 43763 27047
rect 6377 26945 6411 26979
rect 8585 26945 8619 26979
rect 8861 26945 8895 26979
rect 9045 26945 9079 26979
rect 14841 26945 14875 26979
rect 15025 26945 15059 26979
rect 18153 26945 18187 26979
rect 20545 26945 20579 26979
rect 24133 26945 24167 26979
rect 24409 26945 24443 26979
rect 24665 26945 24699 26979
rect 28641 26945 28675 26979
rect 29377 26945 29411 26979
rect 30573 26945 30607 26979
rect 34621 26945 34655 26979
rect 35725 26945 35759 26979
rect 35817 26945 35851 26979
rect 35909 26945 35943 26979
rect 36185 26945 36219 26979
rect 36277 26945 36311 26979
rect 36461 26945 36495 26979
rect 42441 26945 42475 26979
rect 42717 26945 42751 26979
rect 42809 26945 42843 26979
rect 43453 26945 43487 26979
rect 43913 26945 43947 26979
rect 8769 26877 8803 26911
rect 12081 26877 12115 26911
rect 20729 26877 20763 26911
rect 22845 26877 22879 26911
rect 23029 26877 23063 26911
rect 27445 26877 27479 26911
rect 27537 26877 27571 26911
rect 28733 26877 28767 26911
rect 29653 26877 29687 26911
rect 30205 26877 30239 26911
rect 34345 26877 34379 26911
rect 36369 26877 36403 26911
rect 43545 26877 43579 26911
rect 8125 26809 8159 26843
rect 24317 26809 24351 26843
rect 30665 26809 30699 26843
rect 44097 26809 44131 26843
rect 11529 26741 11563 26775
rect 17969 26741 18003 26775
rect 42993 26741 43027 26775
rect 43085 26741 43119 26775
rect 11529 26537 11563 26571
rect 16313 26537 16347 26571
rect 18521 26537 18555 26571
rect 28825 26537 28859 26571
rect 29561 26537 29595 26571
rect 30021 26537 30055 26571
rect 35081 26537 35115 26571
rect 35725 26537 35759 26571
rect 41521 26537 41555 26571
rect 44741 26537 44775 26571
rect 22937 26469 22971 26503
rect 24225 26469 24259 26503
rect 33425 26469 33459 26503
rect 42165 26469 42199 26503
rect 10977 26401 11011 26435
rect 12173 26401 12207 26435
rect 16773 26401 16807 26435
rect 20545 26401 20579 26435
rect 21373 26401 21407 26435
rect 21557 26401 21591 26435
rect 23581 26401 23615 26435
rect 24685 26401 24719 26435
rect 29653 26401 29687 26435
rect 30573 26401 30607 26435
rect 32321 26401 32355 26435
rect 32965 26401 32999 26435
rect 33149 26401 33183 26435
rect 33793 26401 33827 26435
rect 33977 26401 34011 26435
rect 34437 26401 34471 26435
rect 39221 26401 39255 26435
rect 40141 26401 40175 26435
rect 41061 26401 41095 26435
rect 41153 26401 41187 26435
rect 42533 26401 42567 26435
rect 42993 26401 43027 26435
rect 10701 26333 10735 26367
rect 11989 26333 12023 26367
rect 15761 26333 15795 26367
rect 16405 26333 16439 26367
rect 20453 26333 20487 26367
rect 24041 26333 24075 26367
rect 24409 26333 24443 26367
rect 29009 26333 29043 26367
rect 29101 26333 29135 26367
rect 29193 26333 29227 26367
rect 29285 26333 29319 26367
rect 29837 26333 29871 26367
rect 33701 26333 33735 26367
rect 34069 26333 34103 26367
rect 34529 26333 34563 26367
rect 34713 26333 34747 26367
rect 34897 26333 34931 26367
rect 35541 26333 35575 26367
rect 37473 26333 37507 26367
rect 39313 26333 39347 26367
rect 39865 26333 39899 26367
rect 40049 26333 40083 26367
rect 40233 26333 40267 26367
rect 40417 26333 40451 26367
rect 40693 26333 40727 26367
rect 40877 26333 40911 26367
rect 41245 26333 41279 26367
rect 41429 26333 41463 26367
rect 41705 26333 41739 26367
rect 41889 26333 41923 26367
rect 42073 26333 42107 26367
rect 42349 26333 42383 26367
rect 42625 26333 42659 26367
rect 42717 26333 42751 26367
rect 42901 26333 42935 26367
rect 10793 26265 10827 26299
rect 11897 26265 11931 26299
rect 15485 26265 15519 26299
rect 17049 26265 17083 26299
rect 20361 26265 20395 26299
rect 20821 26265 20855 26299
rect 21802 26265 21836 26299
rect 29561 26265 29595 26299
rect 30849 26265 30883 26299
rect 35357 26265 35391 26299
rect 37749 26265 37783 26299
rect 39497 26265 39531 26299
rect 39681 26265 39715 26299
rect 40601 26265 40635 26299
rect 41797 26265 41831 26299
rect 43269 26265 43303 26299
rect 10333 26197 10367 26231
rect 19993 26197 20027 26231
rect 23029 26197 23063 26231
rect 26157 26197 26191 26231
rect 32413 26197 32447 26231
rect 33609 26197 33643 26231
rect 33977 26197 34011 26231
rect 34161 26197 34195 26231
rect 17233 25993 17267 26027
rect 17601 25993 17635 26027
rect 17969 25993 18003 26027
rect 19717 25993 19751 26027
rect 21189 25993 21223 26027
rect 21649 25993 21683 26027
rect 21833 25993 21867 26027
rect 22201 25993 22235 26027
rect 24225 25993 24259 26027
rect 24593 25993 24627 26027
rect 26801 25993 26835 26027
rect 29653 25993 29687 26027
rect 31309 25993 31343 26027
rect 32505 25993 32539 26027
rect 37841 25993 37875 26027
rect 40233 25993 40267 26027
rect 40969 25993 41003 26027
rect 42441 25993 42475 26027
rect 43269 25993 43303 26027
rect 20076 25925 20110 25959
rect 27261 25925 27295 25959
rect 31861 25925 31895 25959
rect 31953 25925 31987 25959
rect 39865 25925 39899 25959
rect 41153 25925 41187 25959
rect 41337 25925 41371 25959
rect 13010 25857 13044 25891
rect 13277 25857 13311 25891
rect 13737 25857 13771 25891
rect 16313 25857 16347 25891
rect 17417 25857 17451 25891
rect 18061 25857 18095 25891
rect 19257 25857 19291 25891
rect 19533 25857 19567 25891
rect 21465 25857 21499 25891
rect 23581 25857 23615 25891
rect 26617 25857 26651 25891
rect 29469 25857 29503 25891
rect 31585 25857 31619 25891
rect 32229 25857 32263 25891
rect 32321 25857 32355 25891
rect 32597 25857 32631 25891
rect 32965 25857 32999 25891
rect 33701 25857 33735 25891
rect 33977 25857 34011 25891
rect 39313 25857 39347 25891
rect 39405 25857 39439 25891
rect 39589 25857 39623 25891
rect 39681 25857 39715 25891
rect 39957 25857 39991 25891
rect 40049 25857 40083 25891
rect 42625 25857 42659 25891
rect 42717 25857 42751 25891
rect 42901 25857 42935 25891
rect 42993 25857 43027 25891
rect 43821 25857 43855 25891
rect 7481 25789 7515 25823
rect 7757 25789 7791 25823
rect 9413 25789 9447 25823
rect 9689 25789 9723 25823
rect 11161 25789 11195 25823
rect 13829 25789 13863 25823
rect 13921 25789 13955 25823
rect 16037 25789 16071 25823
rect 18245 25789 18279 25823
rect 19809 25789 19843 25823
rect 22293 25789 22327 25823
rect 22477 25789 22511 25823
rect 22845 25789 22879 25823
rect 23489 25789 23523 25823
rect 24685 25789 24719 25823
rect 24777 25789 24811 25823
rect 26985 25789 27019 25823
rect 29193 25789 29227 25823
rect 31493 25789 31527 25823
rect 34069 25789 34103 25823
rect 38393 25789 38427 25823
rect 44557 25789 44591 25823
rect 9229 25653 9263 25687
rect 11897 25653 11931 25687
rect 13369 25653 13403 25687
rect 15393 25653 15427 25687
rect 16129 25653 16163 25687
rect 19441 25653 19475 25687
rect 23765 25653 23799 25687
rect 28733 25653 28767 25687
rect 29285 25653 29319 25687
rect 38669 25653 38703 25687
rect 39497 25653 39531 25687
rect 44005 25653 44039 25687
rect 8217 25449 8251 25483
rect 9873 25449 9907 25483
rect 11897 25449 11931 25483
rect 12817 25449 12851 25483
rect 15564 25449 15598 25483
rect 17049 25449 17083 25483
rect 19073 25449 19107 25483
rect 20913 25449 20947 25483
rect 26709 25449 26743 25483
rect 29561 25449 29595 25483
rect 31769 25449 31803 25483
rect 32873 25449 32907 25483
rect 37841 25449 37875 25483
rect 43361 25449 43395 25483
rect 11713 25381 11747 25415
rect 31677 25381 31711 25415
rect 33149 25381 33183 25415
rect 34253 25381 34287 25415
rect 42257 25381 42291 25415
rect 9597 25313 9631 25347
rect 10333 25313 10367 25347
rect 12449 25313 12483 25347
rect 14749 25313 14783 25347
rect 15301 25313 15335 25347
rect 17325 25313 17359 25347
rect 23857 25313 23891 25347
rect 24133 25313 24167 25347
rect 27261 25313 27295 25347
rect 29101 25313 29135 25347
rect 29377 25313 29411 25347
rect 33241 25313 33275 25347
rect 36277 25313 36311 25347
rect 36553 25313 36587 25347
rect 38209 25313 38243 25347
rect 43913 25313 43947 25347
rect 8401 25245 8435 25279
rect 9321 25245 9355 25279
rect 10057 25245 10091 25279
rect 12633 25245 12667 25279
rect 13829 25245 13863 25279
rect 14565 25245 14599 25279
rect 19533 25245 19567 25279
rect 19789 25245 19823 25279
rect 29009 25245 29043 25279
rect 29745 25245 29779 25279
rect 31493 25245 31527 25279
rect 31677 25245 31711 25279
rect 31953 25245 31987 25279
rect 32045 25245 32079 25279
rect 32689 25245 32723 25279
rect 33057 25245 33091 25279
rect 33333 25245 33367 25279
rect 33517 25245 33551 25279
rect 33701 25245 33735 25279
rect 34069 25245 34103 25279
rect 38117 25245 38151 25279
rect 41981 25245 42015 25279
rect 42073 25245 42107 25279
rect 42257 25245 42291 25279
rect 42901 25245 42935 25279
rect 43177 25245 43211 25279
rect 44557 25245 44591 25279
rect 44649 25245 44683 25279
rect 44833 25245 44867 25279
rect 10600 25177 10634 25211
rect 14473 25177 14507 25211
rect 17601 25177 17635 25211
rect 27077 25177 27111 25211
rect 29929 25177 29963 25211
rect 32505 25177 32539 25211
rect 33885 25177 33919 25211
rect 33977 25177 34011 25211
rect 8953 25109 8987 25143
rect 9413 25109 9447 25143
rect 13645 25109 13679 25143
rect 14105 25109 14139 25143
rect 22385 25109 22419 25143
rect 27169 25109 27203 25143
rect 32413 25109 32447 25143
rect 34805 25109 34839 25143
rect 42349 25109 42383 25143
rect 44741 25109 44775 25143
rect 10885 24905 10919 24939
rect 11529 24905 11563 24939
rect 14749 24905 14783 24939
rect 16221 24905 16255 24939
rect 16773 24905 16807 24939
rect 17141 24905 17175 24939
rect 17693 24905 17727 24939
rect 18337 24905 18371 24939
rect 19901 24905 19935 24939
rect 20269 24905 20303 24939
rect 23029 24905 23063 24939
rect 23397 24905 23431 24939
rect 24869 24905 24903 24939
rect 27261 24905 27295 24939
rect 29009 24905 29043 24939
rect 30389 24905 30423 24939
rect 33609 24905 33643 24939
rect 34437 24905 34471 24939
rect 42993 24905 43027 24939
rect 25237 24837 25271 24871
rect 32413 24837 32447 24871
rect 32597 24837 32631 24871
rect 38853 24837 38887 24871
rect 42625 24837 42659 24871
rect 42825 24837 42859 24871
rect 11069 24769 11103 24803
rect 12081 24769 12115 24803
rect 13001 24769 13035 24803
rect 14841 24769 14875 24803
rect 15108 24769 15142 24803
rect 17877 24769 17911 24803
rect 22569 24769 22603 24803
rect 22937 24769 22971 24803
rect 24685 24769 24719 24803
rect 28733 24769 28767 24803
rect 29193 24769 29227 24803
rect 29837 24769 29871 24803
rect 30573 24769 30607 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32781 24769 32815 24803
rect 32873 24769 32907 24803
rect 33057 24769 33091 24803
rect 33333 24769 33367 24803
rect 33425 24769 33459 24803
rect 34989 24769 35023 24803
rect 38117 24769 38151 24803
rect 38209 24769 38243 24803
rect 38393 24769 38427 24803
rect 38669 24769 38703 24803
rect 39037 24769 39071 24803
rect 39129 24769 39163 24803
rect 39313 24769 39347 24803
rect 40509 24769 40543 24803
rect 40601 24769 40635 24803
rect 40785 24769 40819 24803
rect 41705 24769 41739 24803
rect 41889 24769 41923 24803
rect 43085 24769 43119 24803
rect 13277 24701 13311 24735
rect 17233 24701 17267 24735
rect 17417 24701 17451 24735
rect 18429 24701 18463 24735
rect 18613 24701 18647 24735
rect 20361 24701 20395 24735
rect 20545 24701 20579 24735
rect 21925 24701 21959 24735
rect 22845 24701 22879 24735
rect 24961 24701 24995 24735
rect 29469 24701 29503 24735
rect 29745 24701 29779 24735
rect 30205 24701 30239 24735
rect 33241 24701 33275 24735
rect 33609 24701 33643 24735
rect 38577 24701 38611 24735
rect 17969 24633 18003 24667
rect 32137 24633 32171 24667
rect 39221 24633 39255 24667
rect 26709 24565 26743 24599
rect 29377 24565 29411 24599
rect 37933 24565 37967 24599
rect 40785 24565 40819 24599
rect 41705 24565 41739 24599
rect 42809 24565 42843 24599
rect 44557 24565 44591 24599
rect 15025 24361 15059 24395
rect 19257 24361 19291 24395
rect 24869 24361 24903 24395
rect 29285 24361 29319 24395
rect 29745 24361 29779 24395
rect 37644 24361 37678 24395
rect 39129 24361 39163 24395
rect 40049 24361 40083 24395
rect 42901 24361 42935 24395
rect 11621 24293 11655 24327
rect 40969 24293 41003 24327
rect 10057 24225 10091 24259
rect 12357 24225 12391 24259
rect 14381 24225 14415 24259
rect 15761 24225 15795 24259
rect 18429 24225 18463 24259
rect 19073 24225 19107 24259
rect 25421 24225 25455 24259
rect 35541 24225 35575 24259
rect 37381 24225 37415 24259
rect 41061 24225 41095 24259
rect 42809 24225 42843 24259
rect 44373 24225 44407 24259
rect 44649 24225 44683 24259
rect 10425 24157 10459 24191
rect 10885 24157 10919 24191
rect 11805 24157 11839 24191
rect 12081 24157 12115 24191
rect 14105 24157 14139 24191
rect 14841 24157 14875 24191
rect 15485 24157 15519 24191
rect 15577 24157 15611 24191
rect 18061 24157 18095 24191
rect 19809 24157 19843 24191
rect 26249 24157 26283 24191
rect 28089 24157 28123 24191
rect 28181 24157 28215 24191
rect 28365 24157 28399 24191
rect 29193 24157 29227 24191
rect 29653 24157 29687 24191
rect 29837 24157 29871 24191
rect 32689 24157 32723 24191
rect 33057 24157 33091 24191
rect 39405 24157 39439 24191
rect 39589 24157 39623 24191
rect 40417 24157 40451 24191
rect 9873 24089 9907 24123
rect 17794 24089 17828 24123
rect 25237 24089 25271 24123
rect 27905 24089 27939 24123
rect 32873 24089 32907 24123
rect 32965 24089 32999 24123
rect 35817 24089 35851 24123
rect 40233 24089 40267 24123
rect 41337 24089 41371 24123
rect 9413 24021 9447 24055
rect 9781 24021 9815 24055
rect 10241 24021 10275 24055
rect 10609 24021 10643 24055
rect 11897 24021 11931 24055
rect 12449 24021 12483 24055
rect 12541 24021 12575 24055
rect 12909 24021 12943 24055
rect 15117 24021 15151 24055
rect 16681 24021 16715 24055
rect 25329 24021 25363 24055
rect 25697 24021 25731 24055
rect 27721 24021 27755 24055
rect 28273 24021 28307 24055
rect 33241 24021 33275 24055
rect 37289 24021 37323 24055
rect 39497 24021 39531 24055
rect 39865 24021 39899 24055
rect 40033 24021 40067 24055
rect 10609 23817 10643 23851
rect 10977 23817 11011 23851
rect 12265 23817 12299 23851
rect 12633 23817 12667 23851
rect 13093 23817 13127 23851
rect 16865 23817 16899 23851
rect 17601 23817 17635 23851
rect 18429 23817 18463 23851
rect 35449 23817 35483 23851
rect 38209 23817 38243 23851
rect 40509 23817 40543 23851
rect 41337 23817 41371 23851
rect 42165 23817 42199 23851
rect 42809 23817 42843 23851
rect 12725 23749 12759 23783
rect 24041 23749 24075 23783
rect 25789 23749 25823 23783
rect 26525 23749 26559 23783
rect 32321 23749 32355 23783
rect 32873 23749 32907 23783
rect 33701 23749 33735 23783
rect 35265 23749 35299 23783
rect 37289 23749 37323 23783
rect 39037 23749 39071 23783
rect 10517 23681 10551 23715
rect 11069 23681 11103 23715
rect 12173 23681 12207 23715
rect 17417 23681 17451 23715
rect 17785 23681 17819 23715
rect 19717 23681 19751 23715
rect 19809 23681 19843 23715
rect 20076 23681 20110 23715
rect 22744 23681 22778 23715
rect 26985 23681 27019 23715
rect 32137 23681 32171 23715
rect 32413 23681 32447 23715
rect 32505 23681 32539 23715
rect 33609 23681 33643 23715
rect 35173 23681 35207 23715
rect 35357 23681 35391 23715
rect 35633 23681 35667 23715
rect 35725 23681 35759 23715
rect 35817 23681 35851 23715
rect 36001 23681 36035 23715
rect 36093 23681 36127 23715
rect 36277 23681 36311 23715
rect 38117 23681 38151 23715
rect 38761 23681 38795 23715
rect 41061 23681 41095 23715
rect 41245 23681 41279 23715
rect 42073 23681 42107 23715
rect 42257 23681 42291 23715
rect 44557 23681 44591 23715
rect 44833 23681 44867 23715
rect 11253 23613 11287 23647
rect 11529 23613 11563 23647
rect 12817 23613 12851 23647
rect 13645 23613 13679 23647
rect 22477 23613 22511 23647
rect 27261 23613 27295 23647
rect 28733 23613 28767 23647
rect 29377 23613 29411 23647
rect 33425 23613 33459 23647
rect 36553 23613 36587 23647
rect 37841 23613 37875 23647
rect 41889 23613 41923 23647
rect 44281 23613 44315 23647
rect 21189 23545 21223 23579
rect 32689 23545 32723 23579
rect 40877 23545 40911 23579
rect 9045 23477 9079 23511
rect 23857 23477 23891 23511
rect 26249 23477 26283 23511
rect 28825 23477 28859 23511
rect 36461 23477 36495 23511
rect 44649 23477 44683 23511
rect 11069 23273 11103 23307
rect 11345 23273 11379 23307
rect 14473 23273 14507 23307
rect 17417 23273 17451 23307
rect 19625 23273 19659 23307
rect 22385 23273 22419 23307
rect 27537 23273 27571 23307
rect 29745 23273 29779 23307
rect 31401 23273 31435 23307
rect 32689 23273 32723 23307
rect 36461 23273 36495 23307
rect 39221 23273 39255 23307
rect 41981 23273 42015 23307
rect 43269 23273 43303 23307
rect 29377 23205 29411 23239
rect 29929 23205 29963 23239
rect 31953 23205 31987 23239
rect 9321 23137 9355 23171
rect 9597 23137 9631 23171
rect 14657 23137 14691 23171
rect 16773 23137 16807 23171
rect 20453 23137 20487 23171
rect 23029 23137 23063 23171
rect 24961 23137 24995 23171
rect 28181 23137 28215 23171
rect 30941 23137 30975 23171
rect 34161 23137 34195 23171
rect 40233 23137 40267 23171
rect 9137 23069 9171 23103
rect 12725 23069 12759 23103
rect 13001 23069 13035 23103
rect 17509 23069 17543 23103
rect 19441 23069 19475 23103
rect 20269 23069 20303 23103
rect 20729 23069 20763 23103
rect 21005 23069 21039 23103
rect 22937 23069 22971 23103
rect 24685 23069 24719 23103
rect 27721 23069 27755 23103
rect 27813 23069 27847 23103
rect 29101 23069 29135 23103
rect 30113 23069 30147 23103
rect 30297 23069 30331 23103
rect 30573 23069 30607 23103
rect 31033 23069 31067 23103
rect 32597 23069 32631 23103
rect 34437 23069 34471 23103
rect 36369 23069 36403 23103
rect 36553 23069 36587 23103
rect 43177 23069 43211 23103
rect 12480 23001 12514 23035
rect 14197 23001 14231 23035
rect 14933 23001 14967 23035
rect 17049 23001 17083 23035
rect 17776 23001 17810 23035
rect 21250 23001 21284 23035
rect 22845 23001 22879 23035
rect 25237 23001 25271 23035
rect 27905 23001 27939 23035
rect 28043 23001 28077 23035
rect 29193 23001 29227 23035
rect 29377 23001 29411 23035
rect 29561 23001 29595 23035
rect 37933 23001 37967 23035
rect 40509 23001 40543 23035
rect 8953 22933 8987 22967
rect 12817 22933 12851 22967
rect 16405 22933 16439 22967
rect 16957 22933 16991 22967
rect 18889 22933 18923 22967
rect 19901 22933 19935 22967
rect 20361 22933 20395 22967
rect 20913 22933 20947 22967
rect 22477 22933 22511 22967
rect 24869 22933 24903 22967
rect 26709 22933 26743 22967
rect 29761 22933 29795 22967
rect 30757 22933 30791 22967
rect 9781 22729 9815 22763
rect 12909 22729 12943 22763
rect 15025 22729 15059 22763
rect 15669 22729 15703 22763
rect 17877 22729 17911 22763
rect 18521 22729 18555 22763
rect 21833 22729 21867 22763
rect 22201 22729 22235 22763
rect 22845 22729 22879 22763
rect 25145 22729 25179 22763
rect 25513 22729 25547 22763
rect 29469 22729 29503 22763
rect 29837 22729 29871 22763
rect 30573 22729 30607 22763
rect 33885 22729 33919 22763
rect 11796 22661 11830 22695
rect 14381 22661 14415 22695
rect 15761 22661 15795 22695
rect 18613 22661 18647 22695
rect 20545 22661 20579 22695
rect 24685 22661 24719 22695
rect 25053 22661 25087 22695
rect 35357 22661 35391 22695
rect 35771 22661 35805 22695
rect 35909 22661 35943 22695
rect 36001 22661 36035 22695
rect 8033 22593 8067 22627
rect 11529 22593 11563 22627
rect 14473 22593 14507 22627
rect 15209 22593 15243 22627
rect 18061 22593 18095 22627
rect 19533 22593 19567 22627
rect 22661 22593 22695 22627
rect 24409 22593 24443 22627
rect 28641 22593 28675 22627
rect 28825 22593 28859 22627
rect 29101 22593 29135 22627
rect 29377 22593 29411 22627
rect 29653 22593 29687 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 33977 22593 34011 22627
rect 35173 22593 35207 22627
rect 36093 22593 36127 22627
rect 40141 22593 40175 22627
rect 41705 22593 41739 22627
rect 8309 22525 8343 22559
rect 15853 22525 15887 22559
rect 17233 22525 17267 22559
rect 18705 22525 18739 22559
rect 22293 22525 22327 22559
rect 22477 22525 22511 22559
rect 23121 22525 23155 22559
rect 23765 22525 23799 22559
rect 25605 22525 25639 22559
rect 25697 22525 25731 22559
rect 32137 22525 32171 22559
rect 32413 22525 32447 22559
rect 35633 22525 35667 22559
rect 36369 22525 36403 22559
rect 37013 22525 37047 22559
rect 40049 22525 40083 22559
rect 40509 22525 40543 22559
rect 15301 22457 15335 22491
rect 18981 22457 19015 22491
rect 35541 22457 35575 22491
rect 41061 22457 41095 22491
rect 16681 22389 16715 22423
rect 18153 22389 18187 22423
rect 20269 22389 20303 22423
rect 24317 22389 24351 22423
rect 29285 22389 29319 22423
rect 34069 22389 34103 22423
rect 36277 22389 36311 22423
rect 17601 22185 17635 22219
rect 18153 22185 18187 22219
rect 20637 22185 20671 22219
rect 29101 22185 29135 22219
rect 36264 22185 36298 22219
rect 37749 22185 37783 22219
rect 30113 22117 30147 22151
rect 34253 22117 34287 22151
rect 19257 22049 19291 22083
rect 21373 22049 21407 22083
rect 24869 22049 24903 22083
rect 25053 22049 25087 22083
rect 25881 22049 25915 22083
rect 29653 22049 29687 22083
rect 36001 22049 36035 22083
rect 37841 22049 37875 22083
rect 39589 22049 39623 22083
rect 40417 22049 40451 22083
rect 13553 21981 13587 22015
rect 15301 21981 15335 22015
rect 16957 21981 16991 22015
rect 18705 21981 18739 22015
rect 23765 21981 23799 22015
rect 29101 21981 29135 22015
rect 29745 21981 29779 22015
rect 33885 21981 33919 22015
rect 34345 21981 34379 22015
rect 34529 21981 34563 22015
rect 34713 21981 34747 22015
rect 34897 21981 34931 22015
rect 35173 21981 35207 22015
rect 35357 21981 35391 22015
rect 35449 21981 35483 22015
rect 35541 21981 35575 22015
rect 15568 21913 15602 21947
rect 19502 21913 19536 21947
rect 26157 21913 26191 21947
rect 28825 21913 28859 21947
rect 29009 21913 29043 21947
rect 34069 21913 34103 21947
rect 34805 21913 34839 21947
rect 38117 21913 38151 21947
rect 13369 21845 13403 21879
rect 16681 21845 16715 21879
rect 20729 21845 20763 21879
rect 23581 21845 23615 21879
rect 24409 21845 24443 21879
rect 24777 21845 24811 21879
rect 27629 21845 27663 21879
rect 34529 21845 34563 21879
rect 35817 21845 35851 21879
rect 39865 21845 39899 21879
rect 14565 21641 14599 21675
rect 14657 21641 14691 21675
rect 15761 21641 15795 21675
rect 17049 21641 17083 21675
rect 19073 21641 19107 21675
rect 19533 21641 19567 21675
rect 23213 21641 23247 21675
rect 25145 21641 25179 21675
rect 26157 21641 26191 21675
rect 26985 21641 27019 21675
rect 29745 21641 29779 21675
rect 35357 21641 35391 21675
rect 36093 21641 36127 21675
rect 36369 21641 36403 21675
rect 38209 21641 38243 21675
rect 13093 21573 13127 21607
rect 15025 21573 15059 21607
rect 27353 21573 27387 21607
rect 35909 21573 35943 21607
rect 15945 21505 15979 21539
rect 18889 21505 18923 21539
rect 21373 21505 21407 21539
rect 21833 21505 21867 21539
rect 22089 21505 22123 21539
rect 26341 21505 26375 21539
rect 28089 21505 28123 21539
rect 28365 21505 28399 21539
rect 28917 21505 28951 21539
rect 29561 21505 29595 21539
rect 29837 21505 29871 21539
rect 35265 21505 35299 21539
rect 35449 21505 35483 21539
rect 35725 21505 35759 21539
rect 36001 21505 36035 21539
rect 36185 21505 36219 21539
rect 36277 21505 36311 21539
rect 36461 21505 36495 21539
rect 39313 21505 39347 21539
rect 12817 21437 12851 21471
rect 15117 21437 15151 21471
rect 15209 21437 15243 21471
rect 17141 21437 17175 21471
rect 17325 21437 17359 21471
rect 18613 21437 18647 21471
rect 19625 21437 19659 21471
rect 19809 21437 19843 21471
rect 23397 21437 23431 21471
rect 23673 21437 23707 21471
rect 25237 21437 25271 21471
rect 25881 21437 25915 21471
rect 27445 21437 27479 21471
rect 27537 21437 27571 21471
rect 28181 21437 28215 21471
rect 29009 21437 29043 21471
rect 29377 21437 29411 21471
rect 35541 21437 35575 21471
rect 38853 21437 38887 21471
rect 39405 21437 39439 21471
rect 19165 21369 19199 21403
rect 21557 21369 21591 21403
rect 29285 21369 29319 21403
rect 38945 21369 38979 21403
rect 16681 21301 16715 21335
rect 18061 21301 18095 21335
rect 28089 21301 28123 21335
rect 28549 21301 28583 21335
rect 11253 21097 11287 21131
rect 13737 21097 13771 21131
rect 18705 21097 18739 21131
rect 22385 21097 22419 21131
rect 32321 21097 32355 21131
rect 39313 21097 39347 21131
rect 9505 20961 9539 20995
rect 23305 20961 23339 20995
rect 23581 20961 23615 20995
rect 32045 20961 32079 20995
rect 39129 20961 39163 20995
rect 11989 20893 12023 20927
rect 14105 20893 14139 20927
rect 17325 20893 17359 20927
rect 20729 20893 20763 20927
rect 21005 20893 21039 20927
rect 24409 20893 24443 20927
rect 31953 20893 31987 20927
rect 35541 20893 35575 20927
rect 35725 20893 35759 20927
rect 38945 20893 38979 20927
rect 39221 20893 39255 20927
rect 39405 20893 39439 20927
rect 9781 20825 9815 20859
rect 12265 20825 12299 20859
rect 17592 20825 17626 20859
rect 21250 20825 21284 20859
rect 23857 20825 23891 20859
rect 24685 20825 24719 20859
rect 35633 20825 35667 20859
rect 14749 20757 14783 20791
rect 20913 20757 20947 20791
rect 22753 20757 22787 20791
rect 23765 20757 23799 20791
rect 24225 20757 24259 20791
rect 26157 20757 26191 20791
rect 38761 20757 38795 20791
rect 10057 20553 10091 20587
rect 10517 20553 10551 20587
rect 10885 20553 10919 20587
rect 14381 20553 14415 20587
rect 15669 20553 15703 20587
rect 16037 20553 16071 20587
rect 17785 20553 17819 20587
rect 18429 20553 18463 20587
rect 20913 20553 20947 20587
rect 21373 20553 21407 20587
rect 21833 20553 21867 20587
rect 22201 20553 22235 20587
rect 24041 20553 24075 20587
rect 24317 20553 24351 20587
rect 31953 20553 31987 20587
rect 32781 20553 32815 20587
rect 39957 20553 39991 20587
rect 12173 20485 12207 20519
rect 10241 20417 10275 20451
rect 11897 20417 11931 20451
rect 15577 20417 15611 20451
rect 17969 20417 18003 20451
rect 18521 20417 18555 20451
rect 19165 20417 19199 20451
rect 19809 20417 19843 20451
rect 21281 20417 21315 20451
rect 22661 20417 22695 20451
rect 23305 20417 23339 20451
rect 23397 20417 23431 20451
rect 24133 20417 24167 20451
rect 31217 20417 31251 20451
rect 31401 20417 31435 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 32137 20417 32171 20451
rect 32413 20417 32447 20451
rect 32505 20417 32539 20451
rect 36001 20417 36035 20451
rect 36185 20417 36219 20451
rect 37933 20417 37967 20451
rect 38209 20417 38243 20451
rect 10977 20349 11011 20383
rect 11161 20349 11195 20383
rect 14473 20349 14507 20383
rect 14657 20349 14691 20383
rect 16129 20349 16163 20383
rect 16221 20349 16255 20383
rect 18613 20349 18647 20383
rect 21465 20349 21499 20383
rect 22293 20349 22327 20383
rect 22477 20349 22511 20383
rect 31493 20349 31527 20383
rect 32321 20349 32355 20383
rect 32597 20349 32631 20383
rect 38485 20349 38519 20383
rect 12081 20281 12115 20315
rect 14013 20281 14047 20315
rect 18061 20281 18095 20315
rect 38117 20281 38151 20315
rect 13645 20213 13679 20247
rect 15393 20213 15427 20247
rect 31217 20213 31251 20247
rect 36001 20213 36035 20247
rect 28825 20009 28859 20043
rect 29285 20009 29319 20043
rect 32229 20009 32263 20043
rect 32689 20009 32723 20043
rect 34713 20009 34747 20043
rect 35909 20009 35943 20043
rect 38853 20009 38887 20043
rect 13553 19941 13587 19975
rect 15117 19941 15151 19975
rect 19257 19941 19291 19975
rect 35265 19941 35299 19975
rect 15209 19873 15243 19907
rect 16957 19873 16991 19907
rect 19901 19873 19935 19907
rect 29009 19873 29043 19907
rect 29653 19873 29687 19907
rect 31677 19873 31711 19907
rect 31769 19873 31803 19907
rect 35081 19873 35115 19907
rect 35173 19873 35207 19907
rect 35633 19873 35667 19907
rect 37197 19873 37231 19907
rect 10149 19805 10183 19839
rect 12173 19805 12207 19839
rect 14565 19805 14599 19839
rect 17141 19805 17175 19839
rect 17693 19805 17727 19839
rect 18889 19805 18923 19839
rect 19625 19805 19659 19839
rect 22109 19805 22143 19839
rect 22477 19805 22511 19839
rect 26433 19805 26467 19839
rect 29101 19805 29135 19839
rect 29745 19805 29779 19839
rect 31033 19805 31067 19839
rect 31217 19805 31251 19839
rect 31401 19805 31435 19839
rect 31493 19805 31527 19839
rect 31861 19805 31895 19839
rect 32045 19805 32079 19839
rect 32321 19805 32355 19839
rect 32505 19805 32539 19839
rect 33701 19805 33735 19839
rect 33977 19805 34011 19839
rect 34161 19805 34195 19839
rect 34989 19805 35023 19839
rect 35449 19805 35483 19839
rect 35541 19805 35575 19839
rect 35725 19805 35759 19839
rect 36001 19805 36035 19839
rect 36185 19805 36219 19839
rect 37289 19805 37323 19839
rect 39037 19805 39071 19839
rect 10416 19737 10450 19771
rect 12418 19737 12452 19771
rect 15485 19737 15519 19771
rect 24041 19737 24075 19771
rect 28825 19737 28859 19771
rect 39221 19737 39255 19771
rect 11529 19669 11563 19703
rect 18705 19669 18739 19703
rect 19717 19669 19751 19703
rect 21557 19669 21591 19703
rect 26617 19669 26651 19703
rect 30113 19669 30147 19703
rect 31217 19669 31251 19703
rect 33793 19669 33827 19703
rect 36829 19669 36863 19703
rect 36921 19669 36955 19703
rect 10701 19465 10735 19499
rect 11529 19465 11563 19499
rect 11897 19465 11931 19499
rect 12357 19465 12391 19499
rect 12633 19465 12667 19499
rect 13001 19465 13035 19499
rect 14841 19465 14875 19499
rect 14933 19465 14967 19499
rect 15393 19465 15427 19499
rect 17049 19465 17083 19499
rect 17417 19465 17451 19499
rect 19717 19465 19751 19499
rect 20913 19465 20947 19499
rect 28733 19465 28767 19499
rect 29377 19465 29411 19499
rect 31125 19465 31159 19499
rect 31401 19465 31435 19499
rect 31953 19465 31987 19499
rect 34805 19465 34839 19499
rect 34897 19465 34931 19499
rect 35541 19465 35575 19499
rect 13093 19397 13127 19431
rect 18604 19397 18638 19431
rect 21649 19397 21683 19431
rect 22078 19397 22112 19431
rect 26433 19397 26467 19431
rect 27261 19397 27295 19431
rect 36369 19397 36403 19431
rect 37657 19397 37691 19431
rect 10885 19329 10919 19363
rect 12541 19329 12575 19363
rect 13461 19329 13495 19363
rect 13728 19329 13762 19363
rect 15301 19329 15335 19363
rect 16313 19329 16347 19363
rect 16957 19329 16991 19363
rect 17509 19329 17543 19363
rect 20729 19329 20763 19363
rect 21833 19329 21867 19363
rect 23581 19329 23615 19363
rect 23857 19329 23891 19363
rect 26341 19329 26375 19363
rect 26985 19329 27019 19363
rect 28917 19329 28951 19363
rect 29101 19329 29135 19363
rect 29193 19329 29227 19363
rect 29653 19329 29687 19363
rect 30297 19329 30331 19363
rect 30573 19329 30607 19363
rect 30665 19329 30699 19363
rect 30849 19329 30883 19363
rect 31033 19329 31067 19363
rect 31217 19329 31251 19363
rect 31493 19329 31527 19363
rect 31585 19329 31619 19363
rect 31769 19329 31803 19363
rect 33885 19329 33919 19363
rect 34437 19329 34471 19363
rect 35081 19329 35115 19363
rect 35173 19329 35207 19363
rect 35449 19329 35483 19363
rect 35725 19329 35759 19363
rect 35909 19329 35943 19363
rect 36277 19329 36311 19363
rect 36461 19329 36495 19363
rect 36579 19329 36613 19363
rect 36737 19329 36771 19363
rect 36829 19329 36863 19363
rect 37013 19329 37047 19363
rect 37289 19329 37323 19363
rect 37473 19329 37507 19363
rect 11989 19261 12023 19295
rect 12173 19261 12207 19295
rect 13185 19261 13219 19295
rect 15485 19261 15519 19295
rect 16773 19261 16807 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 21097 19261 21131 19295
rect 24133 19261 24167 19295
rect 26249 19261 26283 19295
rect 29745 19261 29779 19295
rect 30113 19261 30147 19295
rect 32137 19261 32171 19295
rect 34345 19261 34379 19295
rect 23765 19193 23799 19227
rect 26801 19193 26835 19227
rect 29009 19193 29043 19227
rect 30021 19193 30055 19227
rect 36921 19193 36955 19227
rect 16129 19125 16163 19159
rect 23213 19125 23247 19159
rect 25605 19125 25639 19159
rect 30481 19125 30515 19159
rect 30757 19125 30791 19159
rect 35357 19125 35391 19159
rect 36093 19125 36127 19159
rect 12449 18921 12483 18955
rect 14105 18921 14139 18955
rect 17049 18921 17083 18955
rect 19257 18921 19291 18955
rect 22017 18921 22051 18955
rect 23489 18921 23523 18955
rect 24409 18921 24443 18955
rect 33425 18921 33459 18955
rect 35725 18921 35759 18955
rect 36093 18921 36127 18955
rect 9321 18853 9355 18887
rect 10057 18853 10091 18887
rect 21925 18853 21959 18887
rect 28181 18853 28215 18887
rect 33149 18853 33183 18887
rect 11805 18785 11839 18819
rect 15209 18785 15243 18819
rect 15669 18785 15703 18819
rect 20545 18785 20579 18819
rect 22661 18785 22695 18819
rect 24041 18785 24075 18819
rect 24869 18785 24903 18819
rect 24961 18785 24995 18819
rect 26709 18785 26743 18819
rect 28641 18785 28675 18819
rect 29377 18785 29411 18819
rect 30665 18785 30699 18819
rect 34713 18785 34747 18819
rect 37841 18785 37875 18819
rect 1409 18717 1443 18751
rect 14289 18717 14323 18751
rect 14657 18717 14691 18751
rect 15936 18717 15970 18751
rect 19073 18717 19107 18751
rect 19809 18717 19843 18751
rect 23213 18717 23247 18751
rect 23857 18717 23891 18751
rect 26525 18717 26559 18751
rect 27813 18717 27847 18751
rect 27997 18717 28031 18751
rect 28549 18717 28583 18751
rect 29653 18717 29687 18751
rect 31862 18695 31896 18729
rect 31953 18717 31987 18751
rect 32321 18717 32355 18751
rect 32781 18717 32815 18751
rect 33057 18717 33091 18751
rect 33241 18717 33275 18751
rect 33517 18717 33551 18751
rect 33885 18717 33919 18751
rect 34345 18717 34379 18751
rect 34897 18717 34931 18751
rect 35081 18717 35115 18751
rect 35173 18717 35207 18751
rect 35265 18717 35299 18751
rect 35541 18717 35575 18751
rect 35633 18717 35667 18751
rect 35817 18717 35851 18751
rect 9689 18649 9723 18683
rect 9781 18649 9815 18683
rect 18828 18649 18862 18683
rect 20790 18649 20824 18683
rect 26617 18649 26651 18683
rect 32045 18649 32079 18683
rect 32183 18649 32217 18683
rect 32965 18649 32999 18683
rect 33977 18649 34011 18683
rect 34069 18649 34103 18683
rect 34207 18649 34241 18683
rect 35449 18649 35483 18683
rect 37565 18649 37599 18683
rect 38301 18649 38335 18683
rect 1593 18581 1627 18615
rect 9229 18581 9263 18615
rect 10241 18581 10275 18615
rect 17693 18581 17727 18615
rect 22385 18581 22419 18615
rect 22477 18581 22511 18615
rect 23397 18581 23431 18615
rect 23949 18581 23983 18615
rect 24777 18581 24811 18615
rect 26157 18581 26191 18615
rect 31677 18581 31711 18615
rect 32597 18581 32631 18615
rect 33701 18581 33735 18615
rect 35357 18581 35391 18615
rect 38209 18581 38243 18615
rect 18337 18377 18371 18411
rect 19809 18377 19843 18411
rect 20637 18377 20671 18411
rect 20729 18377 20763 18411
rect 21097 18377 21131 18411
rect 23765 18377 23799 18411
rect 25605 18377 25639 18411
rect 28641 18377 28675 18411
rect 32781 18377 32815 18411
rect 34253 18377 34287 18411
rect 36001 18377 36035 18411
rect 39313 18377 39347 18411
rect 15117 18309 15151 18343
rect 9873 18241 9907 18275
rect 10793 18241 10827 18275
rect 19257 18241 19291 18275
rect 19533 18241 19567 18275
rect 19625 18241 19659 18275
rect 20453 18241 20487 18275
rect 22109 18241 22143 18275
rect 22385 18241 22419 18275
rect 22641 18241 22675 18275
rect 23857 18241 23891 18275
rect 26157 18241 26191 18275
rect 28825 18241 28859 18275
rect 29101 18241 29135 18275
rect 36093 18241 36127 18275
rect 11713 18173 11747 18207
rect 18705 18173 18739 18207
rect 18797 18173 18831 18207
rect 18981 18173 19015 18207
rect 21189 18173 21223 18207
rect 21373 18173 21407 18207
rect 24133 18173 24167 18207
rect 29009 18173 29043 18207
rect 32137 18173 32171 18207
rect 33609 18173 33643 18207
rect 37565 18173 37599 18207
rect 37841 18173 37875 18207
rect 15393 18105 15427 18139
rect 22293 18105 22327 18139
rect 10057 18037 10091 18071
rect 10977 18037 11011 18071
rect 12357 18037 12391 18071
rect 15577 18037 15611 18071
rect 19349 18037 19383 18071
rect 26341 18037 26375 18071
rect 11529 17833 11563 17867
rect 22201 17833 22235 17867
rect 27721 17833 27755 17867
rect 30941 17833 30975 17867
rect 32781 17833 32815 17867
rect 6929 17765 6963 17799
rect 16313 17765 16347 17799
rect 9781 17697 9815 17731
rect 11621 17697 11655 17731
rect 11897 17697 11931 17731
rect 22753 17697 22787 17731
rect 25973 17697 26007 17731
rect 26249 17697 26283 17731
rect 32413 17697 32447 17731
rect 32689 17697 32723 17731
rect 34253 17697 34287 17731
rect 34529 17697 34563 17731
rect 16129 17629 16163 17663
rect 22569 17629 22603 17663
rect 28917 17629 28951 17663
rect 6653 17561 6687 17595
rect 10057 17561 10091 17595
rect 35817 17561 35851 17595
rect 7113 17493 7147 17527
rect 13369 17493 13403 17527
rect 22661 17493 22695 17527
rect 28365 17493 28399 17527
rect 37105 17493 37139 17527
rect 13277 17289 13311 17323
rect 15761 17289 15795 17323
rect 19809 17289 19843 17323
rect 19993 17289 20027 17323
rect 20453 17289 20487 17323
rect 22477 17289 22511 17323
rect 28733 17289 28767 17323
rect 38117 17289 38151 17323
rect 11805 17221 11839 17255
rect 19257 17221 19291 17255
rect 29653 17221 29687 17255
rect 7481 17153 7515 17187
rect 11529 17153 11563 17187
rect 15117 17153 15151 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 15853 17153 15887 17187
rect 16037 17153 16071 17187
rect 18981 17153 19015 17187
rect 19349 17153 19383 17187
rect 19812 17153 19846 17187
rect 20177 17153 20211 17187
rect 38025 17153 38059 17187
rect 16865 17085 16899 17119
rect 17049 17085 17083 17119
rect 17785 17085 17819 17119
rect 17902 17085 17936 17119
rect 18061 17085 18095 17119
rect 19257 17085 19291 17119
rect 20453 17085 20487 17119
rect 21833 17085 21867 17119
rect 26985 17085 27019 17119
rect 27261 17085 27295 17119
rect 29377 17085 29411 17119
rect 34989 17085 35023 17119
rect 17509 17017 17543 17051
rect 35357 17017 35391 17051
rect 7297 16949 7331 16983
rect 16037 16949 16071 16983
rect 18705 16949 18739 16983
rect 19073 16949 19107 16983
rect 19441 16949 19475 16983
rect 20269 16949 20303 16983
rect 31125 16949 31159 16983
rect 35449 16949 35483 16983
rect 15945 16745 15979 16779
rect 17417 16745 17451 16779
rect 17693 16745 17727 16779
rect 18797 16745 18831 16779
rect 27892 16745 27926 16779
rect 35252 16745 35286 16779
rect 37092 16745 37126 16779
rect 32689 16677 32723 16711
rect 7021 16609 7055 16643
rect 7297 16609 7331 16643
rect 8769 16609 8803 16643
rect 9137 16609 9171 16643
rect 14289 16609 14323 16643
rect 14749 16609 14783 16643
rect 15025 16609 15059 16643
rect 15301 16609 15335 16643
rect 16037 16609 16071 16643
rect 17325 16609 17359 16643
rect 17509 16609 17543 16643
rect 18245 16609 18279 16643
rect 23765 16609 23799 16643
rect 27629 16609 27663 16643
rect 29561 16609 29595 16643
rect 32873 16609 32907 16643
rect 34989 16609 35023 16643
rect 36829 16609 36863 16643
rect 38577 16609 38611 16643
rect 39221 16609 39255 16643
rect 14105 16541 14139 16575
rect 15142 16541 15176 16575
rect 16221 16541 16255 16575
rect 16497 16541 16531 16575
rect 17601 16541 17635 16575
rect 18521 16541 18555 16575
rect 18797 16541 18831 16575
rect 23673 16541 23707 16575
rect 23857 16541 23891 16575
rect 24869 16541 24903 16575
rect 24961 16541 24995 16575
rect 25053 16541 25087 16575
rect 25237 16541 25271 16575
rect 31309 16541 31343 16575
rect 33149 16541 33183 16575
rect 44557 16541 44591 16575
rect 24593 16473 24627 16507
rect 32413 16473 32447 16507
rect 9781 16405 9815 16439
rect 16405 16405 16439 16439
rect 18061 16405 18095 16439
rect 18153 16405 18187 16439
rect 18613 16405 18647 16439
rect 29377 16405 29411 16439
rect 32965 16405 32999 16439
rect 36737 16405 36771 16439
rect 38669 16405 38703 16439
rect 44741 16405 44775 16439
rect 13461 16201 13495 16235
rect 14841 16201 14875 16235
rect 15485 16201 15519 16235
rect 17417 16201 17451 16235
rect 19717 16201 19751 16235
rect 22937 16201 22971 16235
rect 24317 16201 24351 16235
rect 25145 16201 25179 16235
rect 36001 16201 36035 16235
rect 38025 16201 38059 16235
rect 9505 16133 9539 16167
rect 14749 16133 14783 16167
rect 21925 16133 21959 16167
rect 23857 16133 23891 16167
rect 27905 16133 27939 16167
rect 32597 16133 32631 16167
rect 34161 16133 34195 16167
rect 8125 16065 8159 16099
rect 15025 16065 15059 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 16037 16065 16071 16099
rect 16957 16065 16991 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 19441 16065 19475 16099
rect 22109 16065 22143 16099
rect 22293 16065 22327 16099
rect 22385 16065 22419 16099
rect 22753 16065 22787 16099
rect 23121 16065 23155 16099
rect 23213 16065 23247 16099
rect 23397 16065 23431 16099
rect 23489 16065 23523 16099
rect 24685 16065 24719 16099
rect 25329 16065 25363 16099
rect 27629 16065 27663 16099
rect 30573 16065 30607 16099
rect 30757 16065 30791 16099
rect 31401 16065 31435 16099
rect 31670 16065 31704 16099
rect 32321 16065 32355 16099
rect 36185 16065 36219 16099
rect 37289 16065 37323 16099
rect 38485 16065 38519 16099
rect 7205 15997 7239 16031
rect 7665 15997 7699 16031
rect 9229 15997 9263 16031
rect 11253 15997 11287 16031
rect 15301 15997 15335 16031
rect 19717 15997 19751 16031
rect 22477 15997 22511 16031
rect 24777 15997 24811 16031
rect 24869 15997 24903 16031
rect 25421 15997 25455 16031
rect 25513 15997 25547 16031
rect 25605 15997 25639 16031
rect 31493 15997 31527 16031
rect 42993 15997 43027 16031
rect 43545 15997 43579 16031
rect 7481 15929 7515 15963
rect 17601 15929 17635 15963
rect 43821 15929 43855 15963
rect 8309 15861 8343 15895
rect 15209 15861 15243 15895
rect 17233 15861 17267 15895
rect 19533 15861 19567 15895
rect 22569 15861 22603 15895
rect 22661 15861 22695 15895
rect 24133 15861 24167 15895
rect 29377 15861 29411 15895
rect 30757 15861 30791 15895
rect 31677 15861 31711 15895
rect 31861 15861 31895 15895
rect 34069 15861 34103 15895
rect 35633 15861 35667 15895
rect 37933 15861 37967 15895
rect 38393 15861 38427 15895
rect 42441 15861 42475 15895
rect 44005 15861 44039 15895
rect 10701 15657 10735 15691
rect 14565 15657 14599 15691
rect 20545 15657 20579 15691
rect 21005 15657 21039 15691
rect 21281 15657 21315 15691
rect 24225 15657 24259 15691
rect 24409 15657 24443 15691
rect 25329 15657 25363 15691
rect 27169 15657 27203 15691
rect 29975 15657 30009 15691
rect 41613 15657 41647 15691
rect 43637 15657 43671 15691
rect 12633 15589 12667 15623
rect 14197 15589 14231 15623
rect 19625 15589 19659 15623
rect 22017 15589 22051 15623
rect 25973 15589 26007 15623
rect 30113 15589 30147 15623
rect 35817 15589 35851 15623
rect 9229 15521 9263 15555
rect 12081 15521 12115 15555
rect 13277 15521 13311 15555
rect 13369 15521 13403 15555
rect 13645 15521 13679 15555
rect 14381 15521 14415 15555
rect 15301 15521 15335 15555
rect 15577 15521 15611 15555
rect 21649 15521 21683 15555
rect 21741 15521 21775 15555
rect 23949 15521 23983 15555
rect 24961 15521 24995 15555
rect 26525 15521 26559 15555
rect 27261 15521 27295 15555
rect 30205 15521 30239 15555
rect 31585 15521 31619 15555
rect 34713 15521 34747 15555
rect 36001 15521 36035 15555
rect 37473 15521 37507 15555
rect 39129 15521 39163 15555
rect 39865 15521 39899 15555
rect 41889 15521 41923 15555
rect 42165 15521 42199 15555
rect 8953 15453 8987 15487
rect 12219 15453 12253 15487
rect 12357 15453 12391 15487
rect 13093 15453 13127 15487
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 13829 15453 13863 15487
rect 14105 15453 14139 15487
rect 14473 15453 14507 15487
rect 14657 15453 14691 15487
rect 15209 15453 15243 15487
rect 15393 15453 15427 15487
rect 15485 15453 15519 15487
rect 15669 15453 15703 15487
rect 16684 15431 16718 15465
rect 16884 15453 16918 15487
rect 19901 15453 19935 15487
rect 20453 15453 20487 15487
rect 20729 15453 20763 15487
rect 21005 15453 21039 15487
rect 21189 15453 21223 15487
rect 21465 15453 21499 15487
rect 21557 15453 21591 15487
rect 21925 15453 21959 15487
rect 22201 15453 22235 15487
rect 22569 15453 22603 15487
rect 22845 15453 22879 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 23213 15453 23247 15487
rect 23305 15453 23339 15487
rect 23489 15453 23523 15487
rect 23765 15453 23799 15487
rect 23857 15453 23891 15487
rect 24041 15453 24075 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 26985 15453 27019 15487
rect 29837 15453 29871 15487
rect 31033 15453 31067 15487
rect 31309 15453 31343 15487
rect 31493 15453 31527 15487
rect 31769 15453 31803 15487
rect 32045 15453 32079 15487
rect 32229 15453 32263 15487
rect 37749 15453 37783 15487
rect 39497 15453 39531 15487
rect 11437 15385 11471 15419
rect 14381 15385 14415 15419
rect 16967 15385 17001 15419
rect 20913 15385 20947 15419
rect 22293 15385 22327 15419
rect 22385 15385 22419 15419
rect 23397 15385 23431 15419
rect 24777 15385 24811 15419
rect 26801 15385 26835 15419
rect 35449 15385 35483 15419
rect 38644 15385 38678 15419
rect 40141 15385 40175 15419
rect 16773 15317 16807 15351
rect 19809 15317 19843 15351
rect 19993 15317 20027 15351
rect 20177 15317 20211 15351
rect 22661 15317 22695 15351
rect 24869 15317 24903 15351
rect 26341 15317 26375 15351
rect 26433 15317 26467 15351
rect 30481 15317 30515 15351
rect 30849 15317 30883 15351
rect 35357 15317 35391 15351
rect 35909 15317 35943 15351
rect 38485 15317 38519 15351
rect 38761 15317 38795 15351
rect 38853 15317 38887 15351
rect 39681 15317 39715 15351
rect 12173 15113 12207 15147
rect 12725 15113 12759 15147
rect 14565 15113 14599 15147
rect 16957 15113 16991 15147
rect 17969 15113 18003 15147
rect 20545 15113 20579 15147
rect 20913 15113 20947 15147
rect 22661 15113 22695 15147
rect 25605 15113 25639 15147
rect 26985 15113 27019 15147
rect 37289 15113 37323 15147
rect 44281 15113 44315 15147
rect 16865 15045 16899 15079
rect 19809 15045 19843 15079
rect 23305 15045 23339 15079
rect 29469 15045 29503 15079
rect 8401 14977 8435 15011
rect 10149 14977 10183 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12357 14977 12391 15011
rect 12541 14977 12575 15011
rect 13001 14977 13035 15011
rect 13179 14977 13213 15011
rect 13921 14977 13955 15011
rect 14105 14977 14139 15011
rect 14381 14977 14415 15011
rect 16773 14977 16807 15011
rect 17233 14977 17267 15011
rect 17601 14977 17635 15011
rect 19625 14977 19659 15011
rect 20177 14977 20211 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 20821 14977 20855 15011
rect 21005 14977 21039 15011
rect 22845 14977 22879 15011
rect 23121 14977 23155 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 25973 14977 26007 15011
rect 26065 14977 26099 15011
rect 27353 14977 27387 15011
rect 29377 14977 29411 15011
rect 29561 14977 29595 15011
rect 29653 14977 29687 15011
rect 29837 14977 29871 15011
rect 30113 14977 30147 15011
rect 30389 14977 30423 15011
rect 30481 14977 30515 15011
rect 30665 14977 30699 15011
rect 30757 14977 30791 15011
rect 31125 14977 31159 15011
rect 31309 14977 31343 15011
rect 31401 14977 31435 15011
rect 31585 14977 31619 15011
rect 31677 14977 31711 15011
rect 35173 14977 35207 15011
rect 35449 14977 35483 15011
rect 44097 14977 44131 15011
rect 10793 14909 10827 14943
rect 17509 14909 17543 14943
rect 17693 14909 17727 14943
rect 17785 14909 17819 14943
rect 19349 14909 19383 14943
rect 19441 14909 19475 14943
rect 19901 14909 19935 14943
rect 20361 14909 20395 14943
rect 21925 14909 21959 14943
rect 26157 14909 26191 14943
rect 27445 14909 27479 14943
rect 27537 14909 27571 14943
rect 33425 14909 33459 14943
rect 34897 14909 34931 14943
rect 35725 14909 35759 14943
rect 37841 14909 37875 14943
rect 13185 14841 13219 14875
rect 14197 14841 14231 14875
rect 14289 14841 14323 14875
rect 20729 14841 20763 14875
rect 10241 14773 10275 14807
rect 17141 14773 17175 14807
rect 17233 14773 17267 14807
rect 19993 14773 20027 14807
rect 22569 14773 22603 14807
rect 23029 14773 23063 14807
rect 30297 14773 30331 14807
rect 30941 14773 30975 14807
rect 35265 14773 35299 14807
rect 36277 14773 36311 14807
rect 8769 14569 8803 14603
rect 11989 14569 12023 14603
rect 12173 14569 12207 14603
rect 14841 14569 14875 14603
rect 15485 14569 15519 14603
rect 15853 14569 15887 14603
rect 16865 14569 16899 14603
rect 17417 14569 17451 14603
rect 17877 14569 17911 14603
rect 19349 14569 19383 14603
rect 20637 14569 20671 14603
rect 25145 14569 25179 14603
rect 26157 14569 26191 14603
rect 27077 14569 27111 14603
rect 29561 14569 29595 14603
rect 31953 14569 31987 14603
rect 36461 14569 36495 14603
rect 14933 14501 14967 14535
rect 17233 14501 17267 14535
rect 17785 14501 17819 14535
rect 7021 14433 7055 14467
rect 8953 14433 8987 14467
rect 9229 14433 9263 14467
rect 11437 14433 11471 14467
rect 14565 14433 14599 14467
rect 15301 14433 15335 14467
rect 15761 14433 15795 14467
rect 16497 14433 16531 14467
rect 16681 14433 16715 14467
rect 17601 14433 17635 14467
rect 17969 14433 18003 14467
rect 20177 14433 20211 14467
rect 20361 14433 20395 14467
rect 20545 14433 20579 14467
rect 20637 14433 20671 14467
rect 25789 14433 25823 14467
rect 26709 14433 26743 14467
rect 30113 14433 30147 14467
rect 34713 14433 34747 14467
rect 34989 14433 35023 14467
rect 12081 14365 12115 14399
rect 12265 14365 12299 14399
rect 14657 14365 14691 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 15853 14365 15887 14399
rect 16405 14365 16439 14399
rect 16865 14365 16899 14399
rect 17049 14365 17083 14399
rect 17325 14365 17359 14399
rect 17693 14365 17727 14399
rect 17877 14365 17911 14399
rect 18613 14365 18647 14399
rect 18889 14365 18923 14399
rect 19257 14365 19291 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 20085 14365 20119 14399
rect 20453 14365 20487 14399
rect 26985 14365 27019 14399
rect 27169 14365 27203 14399
rect 30205 14365 30239 14399
rect 30849 14365 30883 14399
rect 32137 14365 32171 14399
rect 32229 14365 32263 14399
rect 7297 14297 7331 14331
rect 16681 14297 16715 14331
rect 20821 14297 20855 14331
rect 25513 14297 25547 14331
rect 31953 14297 31987 14331
rect 10701 14229 10735 14263
rect 11529 14229 11563 14263
rect 11621 14229 11655 14263
rect 14197 14229 14231 14263
rect 18245 14229 18279 14263
rect 18705 14229 18739 14263
rect 19073 14229 19107 14263
rect 19625 14229 19659 14263
rect 25605 14229 25639 14263
rect 26525 14229 26559 14263
rect 26617 14229 26651 14263
rect 32413 14229 32447 14263
rect 7389 14025 7423 14059
rect 12357 14025 12391 14059
rect 14473 14025 14507 14059
rect 14749 14025 14783 14059
rect 16221 14025 16255 14059
rect 17693 14025 17727 14059
rect 19073 14025 19107 14059
rect 24317 14025 24351 14059
rect 24593 14025 24627 14059
rect 25053 14025 25087 14059
rect 25145 14025 25179 14059
rect 31953 14025 31987 14059
rect 12863 13957 12897 13991
rect 18705 13957 18739 13991
rect 18905 13957 18939 13991
rect 31493 13957 31527 13991
rect 33149 13957 33183 13991
rect 36461 13957 36495 13991
rect 39865 13957 39899 13991
rect 7205 13889 7239 13923
rect 12541 13889 12575 13923
rect 12633 13889 12667 13923
rect 12725 13889 12759 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 14841 13889 14875 13923
rect 15577 13889 15611 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 17417 13889 17451 13923
rect 24317 13889 24351 13923
rect 24501 13889 24535 13923
rect 24869 13889 24903 13923
rect 25237 13889 25271 13923
rect 28917 13889 28951 13923
rect 31769 13889 31803 13923
rect 32873 13889 32907 13923
rect 36737 13889 36771 13923
rect 37841 13889 37875 13923
rect 13001 13821 13035 13855
rect 14013 13821 14047 13855
rect 16681 13821 16715 13855
rect 17325 13821 17359 13855
rect 17693 13821 17727 13855
rect 24777 13821 24811 13855
rect 28733 13821 28767 13855
rect 29101 13821 29135 13855
rect 31677 13821 31711 13855
rect 34989 13821 35023 13855
rect 41153 13753 41187 13787
rect 17509 13685 17543 13719
rect 18889 13685 18923 13719
rect 31493 13685 31527 13719
rect 34621 13685 34655 13719
rect 38104 13685 38138 13719
rect 39589 13685 39623 13719
rect 7113 13481 7147 13515
rect 11897 13481 11931 13515
rect 12817 13481 12851 13515
rect 26617 13481 26651 13515
rect 36921 13481 36955 13515
rect 6929 13413 6963 13447
rect 10701 13413 10735 13447
rect 22017 13413 22051 13447
rect 24133 13413 24167 13447
rect 25329 13413 25363 13447
rect 26065 13413 26099 13447
rect 26433 13413 26467 13447
rect 27261 13413 27295 13447
rect 31585 13413 31619 13447
rect 31677 13413 31711 13447
rect 32229 13413 32263 13447
rect 42349 13413 42383 13447
rect 6653 13345 6687 13379
rect 8953 13345 8987 13379
rect 12909 13334 12943 13368
rect 21925 13345 21959 13379
rect 22661 13345 22695 13379
rect 25053 13345 25087 13379
rect 26157 13345 26191 13379
rect 26709 13345 26743 13379
rect 26893 13345 26927 13379
rect 27077 13345 27111 13379
rect 27721 13345 27755 13379
rect 27813 13345 27847 13379
rect 28641 13345 28675 13379
rect 32413 13345 32447 13379
rect 36277 13345 36311 13379
rect 36645 13345 36679 13379
rect 37657 13345 37691 13379
rect 39865 13345 39899 13379
rect 44097 13345 44131 13379
rect 11437 13277 11471 13311
rect 11529 13277 11563 13311
rect 11713 13277 11747 13311
rect 12633 13277 12667 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 22109 13277 22143 13311
rect 22200 13255 22234 13289
rect 22385 13277 22419 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25881 13277 25915 13311
rect 25973 13277 26007 13311
rect 26801 13277 26835 13311
rect 27169 13277 27203 13311
rect 28549 13277 28583 13311
rect 29285 13277 29319 13311
rect 31493 13277 31527 13311
rect 31769 13277 31803 13311
rect 35633 13277 35667 13311
rect 36553 13277 36587 13311
rect 36737 13277 36771 13311
rect 37013 13277 37047 13311
rect 37289 13277 37323 13311
rect 37473 13277 37507 13311
rect 40601 13277 40635 13311
rect 41153 13277 41187 13311
rect 9229 13209 9263 13243
rect 26893 13209 26927 13243
rect 29101 13209 29135 13243
rect 31953 13209 31987 13243
rect 34805 13209 34839 13243
rect 43821 13209 43855 13243
rect 13093 13141 13127 13175
rect 24501 13141 24535 13175
rect 27629 13141 27663 13175
rect 28089 13141 28123 13175
rect 28457 13141 28491 13175
rect 28917 13141 28951 13175
rect 31309 13141 31343 13175
rect 34897 13141 34931 13175
rect 40509 13141 40543 13175
rect 7941 12937 7975 12971
rect 11529 12937 11563 12971
rect 11713 12937 11747 12971
rect 12265 12937 12299 12971
rect 13191 12937 13225 12971
rect 14749 12937 14783 12971
rect 16221 12937 16255 12971
rect 17509 12937 17543 12971
rect 19625 12937 19659 12971
rect 19901 12937 19935 12971
rect 21097 12937 21131 12971
rect 22753 12937 22787 12971
rect 23213 12937 23247 12971
rect 25329 12937 25363 12971
rect 25789 12937 25823 12971
rect 29469 12937 29503 12971
rect 38945 12937 38979 12971
rect 43545 12937 43579 12971
rect 6837 12869 6871 12903
rect 9689 12869 9723 12903
rect 17785 12869 17819 12903
rect 18337 12869 18371 12903
rect 19809 12869 19843 12903
rect 23581 12869 23615 12903
rect 25697 12869 25731 12903
rect 27721 12869 27755 12903
rect 40417 12869 40451 12903
rect 44373 12869 44407 12903
rect 7757 12801 7791 12835
rect 11161 12801 11195 12835
rect 11345 12801 11379 12835
rect 11710 12801 11744 12835
rect 12173 12801 12207 12835
rect 12541 12801 12575 12835
rect 12633 12801 12667 12835
rect 12725 12801 12759 12835
rect 13093 12801 13127 12835
rect 13277 12801 13311 12835
rect 13369 12801 13403 12835
rect 14657 12801 14691 12835
rect 14841 12801 14875 12835
rect 15117 12801 15151 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 15853 12801 15887 12835
rect 16037 12801 16071 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 17647 12801 17681 12835
rect 17877 12801 17911 12835
rect 18060 12801 18094 12835
rect 18153 12801 18187 12835
rect 18429 12801 18463 12835
rect 19533 12801 19567 12835
rect 20269 12801 20303 12835
rect 20545 12801 20579 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 20913 12801 20947 12835
rect 22293 12801 22327 12835
rect 23121 12801 23155 12835
rect 23857 12801 23891 12835
rect 23949 12801 23983 12835
rect 24041 12801 24075 12835
rect 24225 12801 24259 12835
rect 24317 12801 24351 12835
rect 27445 12801 27479 12835
rect 29653 12801 29687 12835
rect 31033 12801 31067 12835
rect 31217 12801 31251 12835
rect 31309 12801 31343 12835
rect 31493 12801 31527 12835
rect 32229 12801 32263 12835
rect 32413 12801 32447 12835
rect 32689 12801 32723 12835
rect 32781 12801 32815 12835
rect 32873 12801 32907 12835
rect 43361 12801 43395 12835
rect 7297 12733 7331 12767
rect 12449 12733 12483 12767
rect 14933 12733 14967 12767
rect 15301 12733 15335 12767
rect 20085 12733 20119 12767
rect 20177 12733 20211 12767
rect 20361 12733 20395 12767
rect 23397 12733 23431 12767
rect 25881 12733 25915 12767
rect 27721 12733 27755 12767
rect 29837 12733 29871 12767
rect 31769 12733 31803 12767
rect 40693 12733 40727 12767
rect 43913 12733 43947 12767
rect 7113 12665 7147 12699
rect 11345 12665 11379 12699
rect 12081 12665 12115 12699
rect 19809 12665 19843 12699
rect 24501 12665 24535 12699
rect 30849 12665 30883 12699
rect 31677 12665 31711 12699
rect 44097 12665 44131 12699
rect 9597 12597 9631 12631
rect 17049 12597 17083 12631
rect 22477 12597 22511 12631
rect 27537 12597 27571 12631
rect 11897 12393 11931 12427
rect 13645 12393 13679 12427
rect 15117 12393 15151 12427
rect 15393 12393 15427 12427
rect 17417 12393 17451 12427
rect 20821 12393 20855 12427
rect 21189 12393 21223 12427
rect 22477 12393 22511 12427
rect 28457 12393 28491 12427
rect 30113 12393 30147 12427
rect 30757 12393 30791 12427
rect 36093 12393 36127 12427
rect 12449 12325 12483 12359
rect 14381 12325 14415 12359
rect 17233 12325 17267 12359
rect 17509 12325 17543 12359
rect 21649 12325 21683 12359
rect 22661 12325 22695 12359
rect 34805 12325 34839 12359
rect 12265 12257 12299 12291
rect 15761 12257 15795 12291
rect 17417 12257 17451 12291
rect 20453 12257 20487 12291
rect 21373 12257 21407 12291
rect 23121 12257 23155 12291
rect 23305 12257 23339 12291
rect 35173 12257 35207 12291
rect 37841 12257 37875 12291
rect 11805 12189 11839 12223
rect 12081 12189 12115 12223
rect 12357 12189 12391 12223
rect 12633 12189 12667 12223
rect 12909 12189 12943 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14197 12189 14231 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 14933 12189 14967 12223
rect 15209 12189 15243 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 15853 12189 15887 12223
rect 15945 12189 15979 12223
rect 16049 12167 16083 12201
rect 17601 12189 17635 12223
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 20361 12189 20395 12223
rect 20545 12189 20579 12223
rect 20637 12189 20671 12223
rect 21465 12189 21499 12223
rect 22385 12189 22419 12223
rect 22569 12189 22603 12223
rect 28365 12189 28399 12223
rect 28549 12189 28583 12223
rect 29745 12189 29779 12223
rect 30297 12189 30331 12223
rect 30389 12189 30423 12223
rect 30481 12189 30515 12223
rect 30573 12189 30607 12223
rect 30909 12189 30943 12223
rect 31033 12189 31067 12223
rect 31125 12189 31159 12223
rect 31309 12189 31343 12223
rect 31399 12167 31433 12201
rect 31677 12189 31711 12223
rect 31861 12189 31895 12223
rect 31953 12189 31987 12223
rect 32045 12189 32079 12223
rect 32229 12189 32263 12223
rect 11529 12121 11563 12155
rect 11713 12121 11747 12155
rect 19809 12121 19843 12155
rect 21189 12121 21223 12155
rect 29929 12121 29963 12155
rect 37565 12121 37599 12155
rect 11805 12053 11839 12087
rect 12817 12053 12851 12087
rect 16221 12053 16255 12087
rect 19533 12053 19567 12087
rect 23029 12053 23063 12087
rect 29561 12053 29595 12087
rect 31493 12053 31527 12087
rect 34713 12053 34747 12087
rect 11529 11849 11563 11883
rect 12541 11849 12575 11883
rect 13822 11849 13856 11883
rect 14841 11849 14875 11883
rect 15117 11849 15151 11883
rect 19901 11849 19935 11883
rect 20453 11849 20487 11883
rect 24777 11849 24811 11883
rect 25237 11849 25271 11883
rect 27077 11849 27111 11883
rect 29929 11849 29963 11883
rect 31125 11849 31159 11883
rect 19625 11781 19659 11815
rect 20637 11781 20671 11815
rect 27537 11781 27571 11815
rect 28365 11781 28399 11815
rect 30297 11781 30331 11815
rect 35173 11781 35207 11815
rect 11713 11713 11747 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 13645 11713 13679 11747
rect 13737 11713 13771 11747
rect 13921 11713 13955 11747
rect 14473 11713 14507 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 18245 11713 18279 11747
rect 18429 11713 18463 11747
rect 18524 11719 18558 11753
rect 18706 11713 18740 11747
rect 18981 11713 19015 11747
rect 19257 11713 19291 11747
rect 19349 11713 19383 11747
rect 19533 11713 19567 11747
rect 19717 11713 19751 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 20545 11713 20579 11747
rect 20729 11713 20763 11747
rect 25145 11713 25179 11747
rect 25973 11713 26007 11747
rect 27445 11713 27479 11747
rect 28641 11713 28675 11747
rect 29009 11713 29043 11747
rect 29193 11713 29227 11747
rect 30113 11713 30147 11747
rect 30481 11713 30515 11747
rect 30573 11713 30607 11747
rect 30665 11713 30699 11747
rect 31309 11713 31343 11747
rect 31493 11713 31527 11747
rect 31585 11713 31619 11747
rect 32229 11713 32263 11747
rect 32505 11713 32539 11747
rect 37841 11713 37875 11747
rect 11805 11645 11839 11679
rect 11897 11645 11931 11679
rect 11989 11645 12023 11679
rect 14565 11645 14599 11679
rect 18889 11645 18923 11679
rect 19165 11645 19199 11679
rect 25421 11645 25455 11679
rect 26065 11645 26099 11679
rect 26157 11645 26191 11679
rect 27629 11645 27663 11679
rect 28365 11645 28399 11679
rect 29101 11645 29135 11679
rect 18797 11577 18831 11611
rect 25605 11577 25639 11611
rect 34989 11577 35023 11611
rect 14657 11509 14691 11543
rect 18061 11509 18095 11543
rect 28549 11509 28583 11543
rect 32413 11509 32447 11543
rect 37289 11509 37323 11543
rect 18981 11305 19015 11339
rect 19257 11305 19291 11339
rect 22201 11305 22235 11339
rect 24869 11305 24903 11339
rect 26985 11305 27019 11339
rect 28641 11305 28675 11339
rect 29009 11305 29043 11339
rect 17785 11237 17819 11271
rect 22661 11237 22695 11271
rect 35633 11237 35667 11271
rect 38117 11237 38151 11271
rect 14565 11169 14599 11203
rect 15025 11169 15059 11203
rect 16129 11169 16163 11203
rect 16589 11169 16623 11203
rect 16982 11169 17016 11203
rect 17141 11169 17175 11203
rect 18245 11169 18279 11203
rect 18521 11169 18555 11203
rect 19717 11169 19751 11203
rect 27445 11169 27479 11203
rect 27537 11169 27571 11203
rect 29101 11169 29135 11203
rect 31769 11169 31803 11203
rect 31861 11169 31895 11203
rect 38209 11169 38243 11203
rect 38761 11169 38795 11203
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 14841 11101 14875 11135
rect 15209 11101 15243 11135
rect 15393 11101 15427 11135
rect 15485 11101 15519 11135
rect 15945 11101 15979 11135
rect 16865 11101 16899 11135
rect 17877 11101 17911 11135
rect 18337 11101 18371 11135
rect 18889 11101 18923 11135
rect 19073 11101 19107 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 19625 11101 19659 11135
rect 22385 11101 22419 11135
rect 22477 11101 22511 11135
rect 22753 11101 22787 11135
rect 25145 11101 25179 11135
rect 25237 11101 25271 11135
rect 25329 11101 25363 11135
rect 25513 11101 25547 11135
rect 28365 11101 28399 11135
rect 28825 11101 28859 11135
rect 30941 11101 30975 11135
rect 31125 11101 31159 11135
rect 31309 11101 31343 11135
rect 31401 11101 31435 11135
rect 31678 11101 31712 11135
rect 31953 11101 31987 11135
rect 32137 11101 32171 11135
rect 32229 11101 32263 11135
rect 32321 11101 32355 11135
rect 34713 11101 34747 11135
rect 36369 11101 36403 11135
rect 38945 11101 38979 11135
rect 27353 11033 27387 11067
rect 28273 11033 28307 11067
rect 31033 11033 31067 11067
rect 35357 11033 35391 11067
rect 35909 11033 35943 11067
rect 36645 11033 36679 11067
rect 17969 10965 18003 10999
rect 18061 10965 18095 10999
rect 30757 10965 30791 10999
rect 31493 10965 31527 10999
rect 35449 10965 35483 10999
rect 39129 10965 39163 10999
rect 16957 10761 16991 10795
rect 19073 10761 19107 10795
rect 22569 10761 22603 10795
rect 22661 10761 22695 10795
rect 23581 10761 23615 10795
rect 25605 10761 25639 10795
rect 28917 10761 28951 10795
rect 31033 10761 31067 10795
rect 32505 10761 32539 10795
rect 33609 10761 33643 10795
rect 37013 10761 37047 10795
rect 22201 10693 22235 10727
rect 23213 10693 23247 10727
rect 23857 10693 23891 10727
rect 26985 10693 27019 10727
rect 35081 10693 35115 10727
rect 39865 10693 39899 10727
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 12449 10625 12483 10659
rect 12541 10625 12575 10659
rect 12909 10625 12943 10659
rect 13369 10625 13403 10659
rect 13553 10625 13587 10659
rect 13737 10625 13771 10659
rect 16221 10625 16255 10659
rect 16405 10625 16439 10659
rect 16497 10625 16531 10659
rect 17141 10625 17175 10659
rect 17417 10625 17451 10659
rect 19349 10625 19383 10659
rect 19625 10625 19659 10659
rect 22937 10625 22971 10659
rect 23397 10625 23431 10659
rect 23673 10625 23707 10659
rect 23945 10647 23979 10681
rect 25973 10625 26007 10659
rect 27169 10625 27203 10659
rect 27261 10625 27295 10659
rect 27430 10625 27464 10659
rect 27527 10625 27561 10659
rect 28365 10625 28399 10659
rect 28825 10625 28859 10659
rect 29469 10625 29503 10659
rect 29561 10625 29595 10659
rect 29745 10625 29779 10659
rect 30021 10625 30055 10659
rect 30205 10625 30239 10659
rect 31033 10625 31067 10659
rect 31217 10625 31251 10659
rect 31493 10625 31527 10659
rect 32137 10625 32171 10659
rect 32229 10625 32263 10659
rect 36921 10625 36955 10659
rect 37105 10625 37139 10659
rect 40141 10625 40175 10659
rect 11713 10557 11747 10591
rect 12633 10557 12667 10591
rect 12725 10557 12759 10591
rect 13829 10557 13863 10591
rect 14013 10557 14047 10591
rect 22017 10557 22051 10591
rect 22109 10557 22143 10591
rect 22661 10557 22695 10591
rect 26065 10557 26099 10591
rect 26249 10557 26283 10591
rect 28549 10557 28583 10591
rect 29193 10557 29227 10591
rect 31953 10557 31987 10591
rect 35357 10557 35391 10591
rect 37289 10557 37323 10591
rect 37841 10557 37875 10591
rect 40509 10557 40543 10591
rect 17233 10489 17267 10523
rect 17325 10489 17359 10523
rect 23673 10489 23707 10523
rect 29561 10489 29595 10523
rect 12265 10421 12299 10455
rect 13369 10421 13403 10455
rect 13921 10421 13955 10455
rect 16221 10421 16255 10455
rect 19717 10421 19751 10455
rect 22845 10421 22879 10455
rect 28181 10421 28215 10455
rect 28733 10421 28767 10455
rect 29377 10421 29411 10455
rect 29929 10421 29963 10455
rect 31677 10421 31711 10455
rect 32229 10421 32263 10455
rect 38393 10421 38427 10455
rect 41153 10421 41187 10455
rect 11069 10217 11103 10251
rect 13553 10217 13587 10251
rect 13921 10217 13955 10251
rect 14933 10217 14967 10251
rect 16497 10217 16531 10251
rect 25697 10217 25731 10251
rect 28641 10217 28675 10251
rect 29009 10217 29043 10251
rect 29193 10217 29227 10251
rect 31125 10217 31159 10251
rect 31585 10217 31619 10251
rect 36737 10217 36771 10251
rect 39589 10217 39623 10251
rect 14565 10149 14599 10183
rect 24501 10149 24535 10183
rect 11713 10081 11747 10115
rect 12265 10081 12299 10115
rect 12725 10081 12759 10115
rect 14473 10081 14507 10115
rect 20085 10081 20119 10115
rect 20545 10081 20579 10115
rect 21005 10081 21039 10115
rect 25053 10081 25087 10115
rect 26341 10081 26375 10115
rect 26500 10081 26534 10115
rect 26617 10081 26651 10115
rect 26893 10081 26927 10115
rect 27537 10081 27571 10115
rect 37289 10081 37323 10115
rect 39221 10081 39255 10115
rect 41337 10081 41371 10115
rect 41613 10081 41647 10115
rect 43453 10081 43487 10115
rect 11872 10013 11906 10047
rect 11989 10013 12023 10047
rect 12909 10013 12943 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 14749 10013 14783 10047
rect 16221 10013 16255 10047
rect 16497 10013 16531 10047
rect 16589 10013 16623 10047
rect 16773 10013 16807 10047
rect 19257 10013 19291 10047
rect 19441 10013 19475 10047
rect 19533 10013 19567 10047
rect 19625 10013 19659 10047
rect 19999 10013 20033 10047
rect 20177 10013 20211 10047
rect 20269 10013 20303 10047
rect 20453 10015 20487 10049
rect 20637 10013 20671 10047
rect 20821 10013 20855 10047
rect 24961 10013 24995 10047
rect 27353 10013 27387 10047
rect 28825 10013 28859 10047
rect 29009 10013 29043 10047
rect 29285 10013 29319 10047
rect 30941 10013 30975 10047
rect 31125 10013 31159 10047
rect 31493 10013 31527 10047
rect 31668 10013 31702 10047
rect 31769 10013 31803 10047
rect 31953 10013 31987 10047
rect 34161 10013 34195 10047
rect 34437 10013 34471 10047
rect 39313 10013 39347 10047
rect 22569 9945 22603 9979
rect 35449 9945 35483 9979
rect 37565 9945 37599 9979
rect 43177 9945 43211 9979
rect 16313 9877 16347 9911
rect 16681 9877 16715 9911
rect 19901 9877 19935 9911
rect 22293 9877 22327 9911
rect 24869 9877 24903 9911
rect 31769 9877 31803 9911
rect 33977 9877 34011 9911
rect 34253 9877 34287 9911
rect 39037 9877 39071 9911
rect 39865 9877 39899 9911
rect 41705 9877 41739 9911
rect 16037 9673 16071 9707
rect 22661 9673 22695 9707
rect 23857 9673 23891 9707
rect 26157 9673 26191 9707
rect 30941 9673 30975 9707
rect 39681 9673 39715 9707
rect 41613 9673 41647 9707
rect 12265 9605 12299 9639
rect 12541 9605 12575 9639
rect 18981 9605 19015 9639
rect 19441 9605 19475 9639
rect 22937 9605 22971 9639
rect 37473 9605 37507 9639
rect 39129 9605 39163 9639
rect 41873 9605 41907 9639
rect 42073 9605 42107 9639
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 12669 9537 12703 9571
rect 13093 9537 13127 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 14289 9537 14323 9571
rect 14565 9537 14599 9571
rect 14841 9537 14875 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 18705 9537 18739 9571
rect 18797 9537 18831 9571
rect 19165 9537 19199 9571
rect 19809 9537 19843 9571
rect 20361 9537 20395 9571
rect 22477 9537 22511 9571
rect 22753 9537 22787 9571
rect 22845 9537 22879 9571
rect 23029 9537 23063 9571
rect 23489 9537 23523 9571
rect 23673 9537 23707 9571
rect 24041 9537 24075 9571
rect 26065 9537 26099 9571
rect 27353 9537 27387 9571
rect 30113 9537 30147 9571
rect 30389 9537 30423 9571
rect 31309 9537 31343 9571
rect 31677 9537 31711 9571
rect 31953 9537 31987 9571
rect 34897 9537 34931 9571
rect 35909 9537 35943 9571
rect 36829 9537 36863 9571
rect 36921 9537 36955 9571
rect 37105 9537 37139 9571
rect 38945 9537 38979 9571
rect 41429 9537 41463 9571
rect 42625 9537 42659 9571
rect 42809 9537 42843 9571
rect 12541 9469 12575 9503
rect 14473 9469 14507 9503
rect 19441 9469 19475 9503
rect 19533 9469 19567 9503
rect 19625 9469 19659 9503
rect 20085 9469 20119 9503
rect 24317 9469 24351 9503
rect 26341 9469 26375 9503
rect 27445 9469 27479 9503
rect 27537 9469 27571 9503
rect 29653 9469 29687 9503
rect 31217 9469 31251 9503
rect 34621 9469 34655 9503
rect 36001 9469 36035 9503
rect 36277 9469 36311 9503
rect 38117 9469 38151 9503
rect 38485 9469 38519 9503
rect 38577 9469 38611 9503
rect 38669 9469 38703 9503
rect 40233 9469 40267 9503
rect 18981 9401 19015 9435
rect 26985 9401 27019 9435
rect 30297 9401 30331 9435
rect 37105 9401 37139 9435
rect 41705 9401 41739 9435
rect 11253 9333 11287 9367
rect 14105 9333 14139 9367
rect 14657 9333 14691 9367
rect 16773 9333 16807 9367
rect 19257 9333 19291 9367
rect 19993 9333 20027 9367
rect 20177 9333 20211 9367
rect 20545 9333 20579 9367
rect 22477 9333 22511 9367
rect 25697 9333 25731 9367
rect 31125 9333 31159 9367
rect 31401 9333 31435 9367
rect 31769 9333 31803 9367
rect 33149 9333 33183 9367
rect 38853 9333 38887 9367
rect 39313 9333 39347 9367
rect 41889 9333 41923 9367
rect 42441 9333 42475 9367
rect 1593 9129 1627 9163
rect 13461 9129 13495 9163
rect 13829 9129 13863 9163
rect 14933 9129 14967 9163
rect 15117 9129 15151 9163
rect 18061 9129 18095 9163
rect 19993 9129 20027 9163
rect 25881 9129 25915 9163
rect 27353 9129 27387 9163
rect 28089 9129 28123 9163
rect 28733 9129 28767 9163
rect 28917 9129 28951 9163
rect 30297 9129 30331 9163
rect 30521 9129 30555 9163
rect 31861 9129 31895 9163
rect 32229 9129 32263 9163
rect 37381 9129 37415 9163
rect 37565 9129 37599 9163
rect 40049 9129 40083 9163
rect 41889 9129 41923 9163
rect 15485 9061 15519 9095
rect 16957 9061 16991 9095
rect 17509 9061 17543 9095
rect 22385 9061 22419 9095
rect 26341 9061 26375 9095
rect 30849 9061 30883 9095
rect 39865 9061 39899 9095
rect 11989 8993 12023 9027
rect 14105 8993 14139 9027
rect 20157 8993 20191 9027
rect 23949 8993 23983 9027
rect 25145 8993 25179 9027
rect 25329 8993 25363 9027
rect 26985 8993 27019 9027
rect 28273 8993 28307 9027
rect 30205 8993 30239 9027
rect 33517 8993 33551 9027
rect 1409 8925 1443 8959
rect 12357 8925 12391 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 13737 8925 13771 8959
rect 13921 8925 13955 8959
rect 14197 8925 14231 8959
rect 14473 8925 14507 8959
rect 15301 8925 15335 8959
rect 15485 8925 15519 8959
rect 16589 8925 16623 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17384 8925 17418 8959
rect 17601 8925 17635 8959
rect 17877 8925 17911 8959
rect 19717 8925 19751 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 22569 8925 22603 8959
rect 22937 8925 22971 8959
rect 23029 8925 23063 8959
rect 23213 8925 23247 8959
rect 25053 8925 25087 8959
rect 26709 8925 26743 8959
rect 27537 8925 27571 8959
rect 28089 8925 28123 8959
rect 28365 8925 28399 8959
rect 28457 8925 28491 8959
rect 29561 8925 29595 8959
rect 29745 8925 29779 8959
rect 29837 8925 29871 8959
rect 29975 8925 30009 8959
rect 30757 8925 30791 8959
rect 30941 8925 30975 8959
rect 31217 8925 31251 8959
rect 31861 8925 31895 8959
rect 32045 8925 32079 8959
rect 32137 8925 32171 8959
rect 32321 8925 32355 8959
rect 38117 8925 38151 8959
rect 38301 8925 38335 8959
rect 41797 8925 41831 8959
rect 41981 8925 42015 8959
rect 42441 8925 42475 8959
rect 42625 8925 42659 8959
rect 42809 8925 42843 8959
rect 11713 8857 11747 8891
rect 14565 8857 14599 8891
rect 16681 8857 16715 8891
rect 19809 8857 19843 8891
rect 19993 8857 20027 8891
rect 20085 8857 20119 8891
rect 22661 8857 22695 8891
rect 22753 8857 22787 8891
rect 23121 8857 23155 8891
rect 23765 8857 23799 8891
rect 25605 8857 25639 8891
rect 26801 8857 26835 8891
rect 28901 8857 28935 8891
rect 29101 8857 29135 8891
rect 30449 8857 30483 8891
rect 30665 8857 30699 8891
rect 31401 8857 31435 8891
rect 37749 8857 37783 8891
rect 40233 8857 40267 8891
rect 42533 8857 42567 8891
rect 12449 8789 12483 8823
rect 14942 8789 14976 8823
rect 17325 8789 17359 8823
rect 17693 8789 17727 8823
rect 23397 8789 23431 8823
rect 23857 8789 23891 8823
rect 24685 8789 24719 8823
rect 31585 8789 31619 8823
rect 31677 8789 31711 8823
rect 34161 8789 34195 8823
rect 37539 8789 37573 8823
rect 38301 8789 38335 8823
rect 40023 8789 40057 8823
rect 42993 8789 43027 8823
rect 15577 8585 15611 8619
rect 17233 8585 17267 8619
rect 17601 8585 17635 8619
rect 21833 8585 21867 8619
rect 24409 8585 24443 8619
rect 24869 8585 24903 8619
rect 25237 8585 25271 8619
rect 25697 8585 25731 8619
rect 26985 8585 27019 8619
rect 27445 8585 27479 8619
rect 28273 8585 28307 8619
rect 31953 8585 31987 8619
rect 42257 8585 42291 8619
rect 43177 8585 43211 8619
rect 11897 8517 11931 8551
rect 28549 8517 28583 8551
rect 31309 8517 31343 8551
rect 34253 8517 34287 8551
rect 36001 8517 36035 8551
rect 41061 8517 41095 8551
rect 41889 8517 41923 8551
rect 42089 8517 42123 8551
rect 12081 8449 12115 8483
rect 14013 8449 14047 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 17049 8449 17083 8483
rect 17325 8449 17359 8483
rect 22017 8449 22051 8483
rect 22109 8449 22143 8483
rect 24777 8449 24811 8483
rect 25605 8449 25639 8483
rect 27353 8449 27387 8483
rect 28181 8449 28215 8483
rect 28365 8449 28399 8483
rect 28641 8449 28675 8483
rect 28917 8449 28951 8483
rect 29193 8449 29227 8483
rect 29469 8449 29503 8483
rect 29653 8449 29687 8483
rect 30020 8449 30054 8483
rect 30113 8449 30147 8483
rect 30205 8449 30239 8483
rect 30389 8449 30423 8483
rect 30665 8449 30699 8483
rect 30849 8449 30883 8483
rect 30941 8449 30975 8483
rect 31125 8449 31159 8483
rect 31585 8449 31619 8483
rect 31739 8449 31773 8483
rect 33425 8449 33459 8483
rect 40325 8449 40359 8483
rect 40509 8449 40543 8483
rect 40601 8449 40635 8483
rect 16957 8381 16991 8415
rect 17417 8381 17451 8415
rect 21833 8381 21867 8415
rect 25053 8381 25087 8415
rect 25789 8381 25823 8415
rect 27537 8381 27571 8415
rect 27997 8381 28031 8415
rect 30757 8381 30791 8415
rect 33793 8381 33827 8415
rect 41613 8381 41647 8415
rect 42993 8381 43027 8415
rect 43729 8381 43763 8415
rect 11713 8313 11747 8347
rect 14289 8313 14323 8347
rect 28733 8313 28767 8347
rect 29745 8313 29779 8347
rect 33977 8313 34011 8347
rect 12265 8245 12299 8279
rect 30481 8245 30515 8279
rect 31493 8245 31527 8279
rect 33609 8245 33643 8279
rect 35909 8245 35943 8279
rect 40325 8245 40359 8279
rect 40785 8245 40819 8279
rect 42073 8245 42107 8279
rect 42441 8245 42475 8279
rect 11713 8041 11747 8075
rect 11989 8041 12023 8075
rect 21833 8041 21867 8075
rect 23305 8041 23339 8075
rect 23949 8041 23983 8075
rect 26709 8041 26743 8075
rect 27537 8041 27571 8075
rect 29745 8041 29779 8075
rect 31217 8041 31251 8075
rect 41889 8041 41923 8075
rect 12633 7973 12667 8007
rect 28365 7973 28399 8007
rect 36461 7973 36495 8007
rect 37013 7973 37047 8007
rect 12357 7905 12391 7939
rect 12449 7905 12483 7939
rect 13093 7905 13127 7939
rect 19349 7905 19383 7939
rect 19809 7905 19843 7939
rect 27261 7905 27295 7939
rect 28089 7905 28123 7939
rect 28733 7905 28767 7939
rect 34713 7905 34747 7939
rect 39865 7905 39899 7939
rect 12173 7837 12207 7871
rect 12541 7837 12575 7871
rect 12909 7837 12943 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 19717 7837 19751 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 20361 7837 20395 7871
rect 21649 7837 21683 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 27077 7837 27111 7871
rect 27905 7837 27939 7871
rect 28549 7837 28583 7871
rect 31125 7837 31159 7871
rect 31309 7837 31343 7871
rect 36553 7837 36587 7871
rect 36737 7837 36771 7871
rect 36829 7837 36863 7871
rect 39313 7837 39347 7871
rect 39497 7837 39531 7871
rect 39681 7837 39715 7871
rect 43637 7837 43671 7871
rect 11805 7769 11839 7803
rect 13277 7769 13311 7803
rect 19993 7769 20027 7803
rect 21465 7769 21499 7803
rect 22017 7769 22051 7803
rect 27169 7769 27203 7803
rect 29929 7769 29963 7803
rect 34989 7769 35023 7803
rect 37013 7769 37047 7803
rect 39589 7769 39623 7803
rect 40141 7769 40175 7803
rect 43361 7769 43395 7803
rect 13369 7701 13403 7735
rect 17693 7701 17727 7735
rect 19441 7701 19475 7735
rect 19533 7701 19567 7735
rect 20545 7701 20579 7735
rect 27997 7701 28031 7735
rect 29561 7701 29595 7735
rect 29729 7701 29763 7735
rect 36829 7701 36863 7735
rect 37473 7701 37507 7735
rect 37565 7701 37599 7735
rect 37749 7701 37783 7735
rect 39129 7701 39163 7735
rect 41613 7701 41647 7735
rect 13298 7497 13332 7531
rect 13737 7497 13771 7531
rect 14841 7497 14875 7531
rect 15485 7497 15519 7531
rect 17417 7497 17451 7531
rect 19533 7497 19567 7531
rect 22937 7497 22971 7531
rect 24869 7497 24903 7531
rect 26985 7497 27019 7531
rect 27353 7497 27387 7531
rect 27445 7497 27479 7531
rect 37013 7497 37047 7531
rect 42625 7497 42659 7531
rect 44281 7497 44315 7531
rect 11161 7429 11195 7463
rect 11805 7429 11839 7463
rect 12357 7429 12391 7463
rect 13093 7429 13127 7463
rect 14657 7429 14691 7463
rect 19257 7429 19291 7463
rect 19809 7429 19843 7463
rect 20177 7429 20211 7463
rect 20361 7429 20395 7463
rect 22017 7429 22051 7463
rect 40233 7429 40267 7463
rect 42993 7429 43027 7463
rect 11069 7361 11103 7395
rect 11345 7361 11379 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12725 7361 12759 7395
rect 13553 7361 13587 7395
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 16957 7361 16991 7395
rect 17509 7361 17543 7395
rect 17693 7361 17727 7395
rect 17969 7361 18003 7395
rect 18153 7361 18187 7395
rect 18429 7361 18463 7395
rect 18613 7361 18647 7395
rect 21189 7361 21223 7395
rect 21925 7361 21959 7395
rect 22109 7361 22143 7395
rect 23489 7361 23523 7395
rect 24869 7361 24903 7395
rect 25513 7361 25547 7395
rect 35817 7361 35851 7395
rect 36185 7361 36219 7395
rect 36737 7361 36771 7395
rect 36921 7361 36955 7395
rect 37105 7361 37139 7395
rect 39129 7361 39163 7395
rect 39313 7361 39347 7395
rect 39681 7361 39715 7395
rect 39957 7361 39991 7395
rect 40417 7361 40451 7395
rect 41337 7361 41371 7395
rect 41521 7361 41555 7395
rect 41797 7361 41831 7395
rect 41981 7361 42015 7395
rect 42257 7361 42291 7395
rect 42441 7361 42475 7395
rect 42717 7361 42751 7395
rect 6929 7293 6963 7327
rect 15117 7293 15151 7327
rect 17049 7293 17083 7327
rect 17141 7293 17175 7327
rect 17233 7293 17267 7327
rect 18245 7293 18279 7327
rect 18521 7293 18555 7327
rect 18705 7293 18739 7327
rect 20913 7293 20947 7327
rect 21097 7293 21131 7327
rect 23213 7293 23247 7327
rect 25789 7293 25823 7327
rect 27537 7293 27571 7327
rect 35449 7293 35483 7327
rect 35909 7293 35943 7327
rect 37289 7293 37323 7327
rect 38761 7293 38795 7327
rect 39037 7293 39071 7327
rect 40601 7293 40635 7327
rect 13461 7225 13495 7259
rect 21557 7225 21591 7259
rect 41337 7225 41371 7259
rect 41613 7225 41647 7259
rect 42441 7225 42475 7259
rect 7573 7157 7607 7191
rect 11345 7157 11379 7191
rect 13277 7157 13311 7191
rect 20453 7157 20487 7191
rect 23397 7157 23431 7191
rect 39589 7157 39623 7191
rect 41797 7157 41831 7191
rect 7959 6953 7993 6987
rect 8953 6953 8987 6987
rect 12633 6953 12667 6987
rect 16037 6953 16071 6987
rect 17049 6953 17083 6987
rect 17417 6953 17451 6987
rect 17969 6953 18003 6987
rect 18797 6953 18831 6987
rect 21281 6953 21315 6987
rect 24041 6953 24075 6987
rect 27353 6953 27387 6987
rect 33805 6953 33839 6987
rect 35068 6953 35102 6987
rect 37289 6953 37323 6987
rect 39037 6953 39071 6987
rect 14381 6885 14415 6919
rect 16221 6885 16255 6919
rect 42809 6885 42843 6919
rect 6469 6817 6503 6851
rect 11897 6817 11931 6851
rect 13553 6817 13587 6851
rect 15577 6817 15611 6851
rect 17877 6817 17911 6851
rect 19901 6817 19935 6851
rect 20177 6817 20211 6851
rect 21097 6817 21131 6851
rect 23029 6817 23063 6851
rect 25421 6817 25455 6851
rect 31585 6817 31619 6851
rect 36553 6817 36587 6851
rect 36737 6817 36771 6851
rect 37565 6817 37599 6851
rect 42441 6817 42475 6851
rect 42901 6817 42935 6851
rect 43085 6817 43119 6851
rect 43361 6817 43395 6851
rect 5733 6749 5767 6783
rect 8217 6749 8251 6783
rect 9505 6749 9539 6783
rect 9965 6749 9999 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 12173 6749 12207 6783
rect 14105 6749 14139 6783
rect 14657 6749 14691 6783
rect 14933 6749 14967 6783
rect 15669 6749 15703 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16209 6749 16243 6783
rect 16405 6749 16439 6783
rect 16497 6749 16531 6783
rect 16589 6749 16623 6783
rect 16773 6749 16807 6783
rect 16865 6749 16899 6783
rect 17325 6749 17359 6783
rect 17601 6749 17635 6783
rect 17693 6749 17727 6783
rect 18153 6749 18187 6783
rect 18245 6749 18279 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 19257 6749 19291 6783
rect 19441 6749 19475 6783
rect 20294 6749 20328 6783
rect 20453 6749 20487 6783
rect 21189 6749 21223 6783
rect 21373 6749 21407 6783
rect 23213 6749 23247 6783
rect 23397 6749 23431 6783
rect 23489 6749 23523 6783
rect 23857 6749 23891 6783
rect 24041 6749 24075 6783
rect 24961 6749 24995 6783
rect 25237 6749 25271 6783
rect 26433 6749 26467 6783
rect 26893 6749 26927 6783
rect 27261 6749 27295 6783
rect 30941 6749 30975 6783
rect 31401 6749 31435 6783
rect 34069 6749 34103 6783
rect 34805 6749 34839 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 39405 6749 39439 6783
rect 11713 6681 11747 6715
rect 12357 6681 12391 6715
rect 12541 6681 12575 6715
rect 13093 6681 13127 6715
rect 13737 6681 13771 6715
rect 13921 6681 13955 6715
rect 18705 6681 18739 6715
rect 26801 6681 26835 6715
rect 31217 6681 31251 6715
rect 39589 6681 39623 6715
rect 6377 6613 6411 6647
rect 9781 6613 9815 6647
rect 13369 6613 13403 6647
rect 23673 6613 23707 6647
rect 25053 6613 25087 6647
rect 31033 6613 31067 6647
rect 32321 6613 32355 6647
rect 38209 6613 38243 6647
rect 38301 6613 38335 6647
rect 39313 6613 39347 6647
rect 44833 6613 44867 6647
rect 4445 6409 4479 6443
rect 8171 6409 8205 6443
rect 14933 6409 14967 6443
rect 15393 6409 15427 6443
rect 17325 6409 17359 6443
rect 19073 6409 19107 6443
rect 23857 6409 23891 6443
rect 37289 6409 37323 6443
rect 37926 6409 37960 6443
rect 42441 6409 42475 6443
rect 43085 6409 43119 6443
rect 44649 6409 44683 6443
rect 14289 6341 14323 6375
rect 15209 6341 15243 6375
rect 17509 6341 17543 6375
rect 19257 6341 19291 6375
rect 19901 6341 19935 6375
rect 24041 6341 24075 6375
rect 24869 6341 24903 6375
rect 24961 6341 24995 6375
rect 33793 6341 33827 6375
rect 37105 6341 37139 6375
rect 37457 6341 37491 6375
rect 37657 6341 37691 6375
rect 38025 6341 38059 6375
rect 6745 6273 6779 6307
rect 13645 6273 13679 6307
rect 14473 6273 14507 6307
rect 14565 6273 14599 6307
rect 15025 6273 15059 6307
rect 15117 6273 15151 6307
rect 15301 6273 15335 6307
rect 16313 6273 16347 6307
rect 17141 6273 17175 6307
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 19073 6273 19107 6307
rect 19349 6273 19383 6307
rect 19993 6273 20027 6307
rect 23581 6273 23615 6307
rect 23765 6273 23799 6307
rect 24409 6273 24443 6307
rect 24685 6273 24719 6307
rect 25053 6273 25087 6307
rect 25789 6273 25823 6307
rect 34069 6273 34103 6307
rect 36921 6273 36955 6307
rect 37749 6273 37783 6307
rect 37841 6273 37875 6307
rect 38117 6273 38151 6307
rect 38209 6273 38243 6307
rect 42625 6273 42659 6307
rect 42717 6273 42751 6307
rect 42809 6273 42843 6307
rect 43361 6273 43395 6307
rect 43545 6273 43579 6307
rect 44833 6273 44867 6307
rect 5917 6205 5951 6239
rect 6193 6205 6227 6239
rect 6377 6205 6411 6239
rect 8309 6205 8343 6239
rect 8585 6205 8619 6239
rect 10057 6205 10091 6239
rect 10241 6205 10275 6239
rect 13001 6205 13035 6239
rect 15577 6205 15611 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 16129 6205 16163 6239
rect 16957 6205 16991 6239
rect 18797 6205 18831 6239
rect 29469 6205 29503 6239
rect 30205 6205 30239 6239
rect 31677 6205 31711 6239
rect 31953 6205 31987 6239
rect 36737 6205 36771 6239
rect 38393 6205 38427 6239
rect 43269 6205 43303 6239
rect 43453 6205 43487 6239
rect 13369 6137 13403 6171
rect 13461 6137 13495 6171
rect 16497 6137 16531 6171
rect 18981 6137 19015 6171
rect 25329 6137 25363 6171
rect 38117 6137 38151 6171
rect 42993 6137 43027 6171
rect 10885 6069 10919 6103
rect 13921 6069 13955 6103
rect 23765 6069 23799 6103
rect 24041 6069 24075 6103
rect 25237 6069 25271 6103
rect 25697 6069 25731 6103
rect 30113 6069 30147 6103
rect 32321 6069 32355 6103
rect 37473 6069 37507 6103
rect 6377 5865 6411 5899
rect 6745 5865 6779 5899
rect 8953 5865 8987 5899
rect 13553 5865 13587 5899
rect 14657 5865 14691 5899
rect 15393 5865 15427 5899
rect 15945 5865 15979 5899
rect 17969 5865 18003 5899
rect 21005 5865 21039 5899
rect 24409 5865 24443 5899
rect 25770 5865 25804 5899
rect 29377 5865 29411 5899
rect 31309 5865 31343 5899
rect 32229 5865 32263 5899
rect 32321 5865 32355 5899
rect 33701 5865 33735 5899
rect 34069 5865 34103 5899
rect 37841 5865 37875 5899
rect 11851 5797 11885 5831
rect 33241 5797 33275 5831
rect 7021 5729 7055 5763
rect 8769 5729 8803 5763
rect 10057 5729 10091 5763
rect 15025 5729 15059 5763
rect 16129 5729 16163 5763
rect 16405 5729 16439 5763
rect 24869 5729 24903 5763
rect 25053 5729 25087 5763
rect 27629 5729 27663 5763
rect 29837 5729 29871 5763
rect 33517 5729 33551 5763
rect 43085 5729 43119 5763
rect 3801 5661 3835 5695
rect 4169 5661 4203 5695
rect 5595 5661 5629 5695
rect 5733 5661 5767 5695
rect 9505 5661 9539 5695
rect 10425 5661 10459 5695
rect 13737 5661 13771 5695
rect 13921 5661 13955 5695
rect 14289 5661 14323 5695
rect 14565 5661 14599 5695
rect 15485 5661 15519 5695
rect 15669 5661 15703 5695
rect 16221 5661 16255 5695
rect 16589 5661 16623 5695
rect 17785 5661 17819 5695
rect 20913 5661 20947 5695
rect 23765 5661 23799 5695
rect 24041 5661 24075 5695
rect 25237 5661 25271 5695
rect 25421 5661 25455 5695
rect 25513 5661 25547 5695
rect 27537 5661 27571 5695
rect 29561 5661 29595 5695
rect 31585 5661 31619 5695
rect 32505 5661 32539 5695
rect 32597 5661 32631 5695
rect 33609 5661 33643 5695
rect 37841 5661 37875 5695
rect 38025 5661 38059 5695
rect 6837 5593 6871 5627
rect 7297 5593 7331 5627
rect 16313 5593 16347 5627
rect 17601 5593 17635 5627
rect 24225 5593 24259 5627
rect 27905 5593 27939 5627
rect 32321 5593 32355 5627
rect 43361 5593 43395 5627
rect 14197 5525 14231 5559
rect 16497 5525 16531 5559
rect 23857 5525 23891 5559
rect 24777 5525 24811 5559
rect 25329 5525 25363 5559
rect 33057 5525 33091 5559
rect 44833 5525 44867 5559
rect 4445 5321 4479 5355
rect 10885 5321 10919 5355
rect 14381 5321 14415 5355
rect 14565 5321 14599 5355
rect 31309 5321 31343 5355
rect 38577 5321 38611 5355
rect 41245 5321 41279 5355
rect 42165 5321 42199 5355
rect 43177 5321 43211 5355
rect 2513 5253 2547 5287
rect 2881 5253 2915 5287
rect 7021 5253 7055 5287
rect 8769 5253 8803 5287
rect 14197 5253 14231 5287
rect 19809 5253 19843 5287
rect 37289 5253 37323 5287
rect 10333 5185 10367 5219
rect 10701 5185 10735 5219
rect 11069 5185 11103 5219
rect 12173 5185 12207 5219
rect 17509 5185 17543 5219
rect 22017 5185 22051 5219
rect 22569 5185 22603 5219
rect 23397 5185 23431 5219
rect 23489 5185 23523 5219
rect 23765 5185 23799 5219
rect 24317 5185 24351 5219
rect 24685 5185 24719 5219
rect 24777 5185 24811 5219
rect 24961 5185 24995 5219
rect 25329 5185 25363 5219
rect 25789 5185 25823 5219
rect 27077 5185 27111 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 36369 5185 36403 5219
rect 41429 5185 41463 5219
rect 41797 5185 41831 5219
rect 41889 5185 41923 5219
rect 42073 5185 42107 5219
rect 42257 5185 42291 5219
rect 42809 5185 42843 5219
rect 43913 5185 43947 5219
rect 1869 5117 1903 5151
rect 2605 5117 2639 5151
rect 4353 5117 4387 5151
rect 4997 5117 5031 5151
rect 17601 5117 17635 5151
rect 21281 5117 21315 5151
rect 21649 5117 21683 5151
rect 25145 5117 25179 5151
rect 25513 5117 25547 5151
rect 25605 5117 25639 5151
rect 29561 5117 29595 5151
rect 29837 5117 29871 5151
rect 36093 5117 36127 5151
rect 39313 5117 39347 5151
rect 39589 5117 39623 5151
rect 41061 5117 41095 5151
rect 42717 5117 42751 5151
rect 44465 5117 44499 5151
rect 17877 5049 17911 5083
rect 24869 5049 24903 5083
rect 25421 5049 25455 5083
rect 27353 5049 27387 5083
rect 36277 5049 36311 5083
rect 8907 4981 8941 5015
rect 11989 4981 12023 5015
rect 14381 4981 14415 5015
rect 21925 4981 21959 5015
rect 23213 4981 23247 5015
rect 23673 4981 23707 5015
rect 23857 4981 23891 5015
rect 24225 4981 24259 5015
rect 24501 4981 24535 5015
rect 34713 4981 34747 5015
rect 36185 4981 36219 5015
rect 41521 4981 41555 5015
rect 1639 4777 1673 4811
rect 21189 4777 21223 4811
rect 23581 4777 23615 4811
rect 23765 4777 23799 4811
rect 35712 4777 35746 4811
rect 37841 4777 37875 4811
rect 38025 4777 38059 4811
rect 38485 4777 38519 4811
rect 39957 4777 39991 4811
rect 40785 4777 40819 4811
rect 40969 4777 41003 4811
rect 42073 4777 42107 4811
rect 13047 4709 13081 4743
rect 13185 4709 13219 4743
rect 18797 4709 18831 4743
rect 20913 4709 20947 4743
rect 42257 4709 42291 4743
rect 3433 4641 3467 4675
rect 9229 4641 9263 4675
rect 11253 4641 11287 4675
rect 11621 4641 11655 4675
rect 13737 4641 13771 4675
rect 18981 4641 19015 4675
rect 19349 4641 19383 4675
rect 20361 4641 20395 4675
rect 20453 4641 20487 4675
rect 21833 4641 21867 4675
rect 22201 4641 22235 4675
rect 33057 4641 33091 4675
rect 35449 4641 35483 4675
rect 39037 4641 39071 4675
rect 40325 4641 40359 4675
rect 3065 4573 3099 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 18705 4573 18739 4607
rect 19257 4573 19291 4607
rect 19441 4573 19475 4607
rect 20545 4573 20579 4607
rect 21005 4573 21039 4607
rect 24041 4573 24075 4607
rect 29561 4573 29595 4607
rect 31309 4573 31343 4607
rect 32781 4573 32815 4607
rect 35265 4573 35299 4607
rect 37381 4573 37415 4607
rect 37473 4573 37507 4607
rect 37841 4573 37875 4607
rect 39865 4573 39899 4607
rect 40049 4573 40083 4607
rect 40141 4573 40175 4607
rect 40509 4573 40543 4607
rect 40693 4573 40727 4607
rect 41245 4573 41279 4607
rect 41337 4573 41371 4607
rect 41429 4573 41463 4607
rect 42698 4573 42732 4607
rect 42993 4573 43027 4607
rect 16865 4505 16899 4539
rect 18613 4505 18647 4539
rect 23765 4505 23799 4539
rect 34713 4505 34747 4539
rect 38301 4505 38335 4539
rect 41153 4505 41187 4539
rect 41889 4505 41923 4539
rect 42105 4505 42139 4539
rect 42349 4505 42383 4539
rect 42533 4505 42567 4539
rect 7849 4437 7883 4471
rect 8953 4437 8987 4471
rect 13553 4437 13587 4471
rect 13645 4437 13679 4471
rect 18981 4437 19015 4471
rect 23949 4437 23983 4471
rect 34529 4437 34563 4471
rect 37197 4437 37231 4471
rect 38501 4437 38535 4471
rect 38669 4437 38703 4471
rect 39681 4437 39715 4471
rect 40943 4437 40977 4471
rect 42809 4437 42843 4471
rect 3801 4233 3835 4267
rect 12633 4233 12667 4267
rect 34897 4233 34931 4267
rect 36527 4233 36561 4267
rect 37289 4233 37323 4267
rect 38669 4233 38703 4267
rect 40877 4233 40911 4267
rect 41613 4233 41647 4267
rect 16773 4165 16807 4199
rect 18521 4165 18555 4199
rect 34437 4165 34471 4199
rect 36277 4165 36311 4199
rect 36737 4165 36771 4199
rect 40141 4165 40175 4199
rect 6377 4097 6411 4131
rect 9321 4097 9355 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 15025 4097 15059 4131
rect 17417 4097 17451 4131
rect 20269 4097 20303 4131
rect 25605 4097 25639 4131
rect 26985 4097 27019 4131
rect 27445 4097 27479 4131
rect 32965 4097 32999 4131
rect 33149 4097 33183 4131
rect 34161 4097 34195 4131
rect 34621 4097 34655 4131
rect 34713 4097 34747 4131
rect 35173 4097 35207 4131
rect 35357 4097 35391 4131
rect 36001 4097 36035 4131
rect 36093 4097 36127 4131
rect 36921 4097 36955 4131
rect 37105 4097 37139 4131
rect 38209 4097 38243 4131
rect 40509 4097 40543 4131
rect 40601 4097 40635 4131
rect 40693 4097 40727 4131
rect 40785 4097 40819 4131
rect 40969 4097 41003 4131
rect 41061 4097 41095 4131
rect 41245 4097 41279 4131
rect 4445 4029 4479 4063
rect 5549 4029 5583 4063
rect 6653 4029 6687 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 9597 4029 9631 4063
rect 11069 4029 11103 4063
rect 12081 4029 12115 4063
rect 13093 4029 13127 4063
rect 13277 4029 13311 4063
rect 14289 4029 14323 4063
rect 17509 4029 17543 4063
rect 18245 4029 18279 4063
rect 20177 4029 20211 4063
rect 20637 4029 20671 4063
rect 28549 4029 28583 4063
rect 28825 4029 28859 4063
rect 30297 4029 30331 4063
rect 33885 4029 33919 4063
rect 34345 4029 34379 4063
rect 37841 4029 37875 4063
rect 38025 4029 38059 4063
rect 40417 4029 40451 4063
rect 42165 4029 42199 4063
rect 42441 4029 42475 4063
rect 42717 4029 42751 4063
rect 44189 4029 44223 4063
rect 15209 3961 15243 3995
rect 19993 3961 20027 3995
rect 33149 3961 33183 3995
rect 36277 3961 36311 3995
rect 36921 3961 36955 3995
rect 6193 3893 6227 3927
rect 8217 3893 8251 3927
rect 11529 3893 11563 3927
rect 14565 3893 14599 3927
rect 17049 3893 17083 3927
rect 17693 3893 17727 3927
rect 25789 3893 25823 3927
rect 27169 3893 27203 3927
rect 27261 3893 27295 3927
rect 33241 3893 33275 3927
rect 33977 3893 34011 3927
rect 34437 3893 34471 3927
rect 35173 3893 35207 3927
rect 36369 3893 36403 3927
rect 36553 3893 36587 3927
rect 38393 3893 38427 3927
rect 41245 3893 41279 3927
rect 7959 3689 7993 3723
rect 8953 3689 8987 3723
rect 9597 3689 9631 3723
rect 13185 3689 13219 3723
rect 16267 3689 16301 3723
rect 26782 3689 26816 3723
rect 29193 3689 29227 3723
rect 29837 3689 29871 3723
rect 32676 3689 32710 3723
rect 34529 3689 34563 3723
rect 37749 3689 37783 3723
rect 39497 3689 39531 3723
rect 28273 3621 28307 3655
rect 3893 3553 3927 3587
rect 4261 3553 4295 3587
rect 8217 3553 8251 3587
rect 9413 3553 9447 3587
rect 10149 3553 10183 3587
rect 10609 3553 10643 3587
rect 10977 3553 11011 3587
rect 12909 3553 12943 3587
rect 14105 3553 14139 3587
rect 18061 3553 18095 3587
rect 18613 3553 18647 3587
rect 23949 3553 23983 3587
rect 24409 3553 24443 3587
rect 26525 3553 26559 3587
rect 28549 3553 28583 3587
rect 30481 3553 30515 3587
rect 32413 3553 32447 3587
rect 35265 3553 35299 3587
rect 35449 3553 35483 3587
rect 35909 3553 35943 3587
rect 37197 3553 37231 3587
rect 39405 3553 39439 3587
rect 39589 3553 39623 3587
rect 9321 3485 9355 3519
rect 12817 3485 12851 3519
rect 13737 3485 13771 3519
rect 16129 3485 16163 3519
rect 17693 3485 17727 3519
rect 18521 3485 18555 3519
rect 23857 3485 23891 3519
rect 26433 3485 26467 3519
rect 30021 3485 30055 3519
rect 30849 3485 30883 3519
rect 34253 3485 34287 3519
rect 34345 3485 34379 3519
rect 35817 3485 35851 3519
rect 36553 3485 36587 3519
rect 38301 3485 38335 3519
rect 38485 3485 38519 3519
rect 38669 3485 38703 3519
rect 39313 3485 39347 3519
rect 5687 3417 5721 3451
rect 15853 3417 15887 3451
rect 24685 3417 24719 3451
rect 34529 3417 34563 3451
rect 34713 3417 34747 3451
rect 6469 3349 6503 3383
rect 12403 3349 12437 3383
rect 13921 3349 13955 3383
rect 18153 3349 18187 3383
rect 24225 3349 24259 3383
rect 32275 3349 32309 3383
rect 34161 3349 34195 3383
rect 38577 3349 38611 3383
rect 4445 3145 4479 3179
rect 12817 3145 12851 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 16957 3145 16991 3179
rect 17325 3145 17359 3179
rect 26065 3145 26099 3179
rect 26709 3145 26743 3179
rect 28825 3145 28859 3179
rect 30665 3145 30699 3179
rect 31401 3145 31435 3179
rect 34713 3145 34747 3179
rect 35005 3145 35039 3179
rect 37105 3145 37139 3179
rect 37565 3145 37599 3179
rect 42073 3145 42107 3179
rect 5917 3077 5951 3111
rect 17417 3077 17451 3111
rect 27261 3077 27295 3111
rect 34805 3077 34839 3111
rect 35633 3077 35667 3111
rect 40601 3077 40635 3111
rect 6193 3009 6227 3043
rect 7665 3009 7699 3043
rect 12173 3009 12207 3043
rect 12633 3009 12667 3043
rect 16313 3009 16347 3043
rect 26985 3009 27019 3043
rect 30573 3009 30607 3043
rect 31493 3009 31527 3043
rect 32781 3009 32815 3043
rect 32965 3009 32999 3043
rect 35357 3009 35391 3043
rect 39313 3009 39347 3043
rect 40325 3009 40359 3043
rect 6929 2941 6963 2975
rect 7573 2941 7607 2975
rect 8033 2941 8067 2975
rect 10241 2941 10275 2975
rect 12265 2941 12299 2975
rect 12541 2941 12575 2975
rect 14841 2941 14875 2975
rect 15025 2941 15059 2975
rect 17601 2941 17635 2975
rect 25605 2941 25639 2975
rect 26249 2941 26283 2975
rect 28733 2941 28767 2975
rect 30297 2941 30331 2975
rect 31125 2941 31159 2975
rect 33241 2941 33275 2975
rect 39037 2941 39071 2975
rect 9459 2873 9493 2907
rect 10517 2873 10551 2907
rect 10701 2873 10735 2907
rect 16497 2873 16531 2907
rect 25881 2873 25915 2907
rect 26617 2873 26651 2907
rect 30849 2873 30883 2907
rect 32597 2805 32631 2839
rect 34989 2805 35023 2839
rect 35173 2805 35207 2839
rect 1593 2601 1627 2635
rect 8493 2601 8527 2635
rect 8769 2601 8803 2635
rect 17693 2601 17727 2635
rect 26709 2601 26743 2635
rect 30205 2601 30239 2635
rect 32689 2601 32723 2635
rect 43913 2601 43947 2635
rect 7205 2465 7239 2499
rect 8217 2465 8251 2499
rect 29561 2465 29595 2499
rect 32229 2465 32263 2499
rect 1409 2397 1443 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 8585 2397 8619 2431
rect 17509 2397 17543 2431
rect 26525 2397 26559 2431
rect 32321 2397 32355 2431
rect 44097 2397 44131 2431
<< metal1 >>
rect 1104 46266 45172 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 45172 46266
rect 1104 46192 45172 46214
rect 14826 46112 14832 46164
rect 14884 46112 14890 46164
rect 934 45976 940 46028
rect 992 46016 998 46028
rect 1397 46019 1455 46025
rect 1397 46016 1409 46019
rect 992 45988 1409 46016
rect 992 45976 998 45988
rect 1397 45985 1409 45988
rect 1443 45985 1455 46019
rect 14844 46016 14872 46112
rect 14844 45988 14964 46016
rect 1397 45979 1455 45985
rect 1670 45908 1676 45960
rect 1728 45908 1734 45960
rect 6454 45908 6460 45960
rect 6512 45948 6518 45960
rect 6549 45951 6607 45957
rect 6549 45948 6561 45951
rect 6512 45920 6561 45948
rect 6512 45908 6518 45920
rect 6549 45917 6561 45920
rect 6595 45917 6607 45951
rect 6549 45911 6607 45917
rect 9858 45908 9864 45960
rect 9916 45908 9922 45960
rect 14826 45908 14832 45960
rect 14884 45908 14890 45960
rect 14936 45957 14964 45988
rect 21818 45976 21824 46028
rect 21876 45976 21882 46028
rect 22281 46019 22339 46025
rect 22281 45985 22293 46019
rect 22327 46016 22339 46019
rect 24118 46016 24124 46028
rect 22327 45988 24124 46016
rect 22327 45985 22339 45988
rect 22281 45979 22339 45985
rect 24118 45976 24124 45988
rect 24176 45976 24182 46028
rect 14921 45951 14979 45957
rect 14921 45917 14933 45951
rect 14967 45917 14979 45951
rect 14921 45911 14979 45917
rect 22186 45908 22192 45960
rect 22244 45908 22250 45960
rect 23842 45908 23848 45960
rect 23900 45948 23906 45960
rect 23937 45951 23995 45957
rect 23937 45948 23949 45951
rect 23900 45920 23949 45948
rect 23900 45908 23906 45920
rect 23937 45917 23949 45920
rect 23983 45917 23995 45951
rect 23937 45911 23995 45917
rect 27617 45951 27675 45957
rect 27617 45917 27629 45951
rect 27663 45917 27675 45951
rect 27617 45911 27675 45917
rect 14553 45883 14611 45889
rect 14553 45849 14565 45883
rect 14599 45880 14611 45883
rect 15930 45880 15936 45892
rect 14599 45852 15936 45880
rect 14599 45849 14611 45852
rect 14553 45843 14611 45849
rect 15930 45840 15936 45852
rect 15988 45840 15994 45892
rect 27632 45880 27660 45911
rect 27890 45908 27896 45960
rect 27948 45948 27954 45960
rect 28353 45951 28411 45957
rect 28353 45948 28365 45951
rect 27948 45920 28365 45948
rect 27948 45908 27954 45920
rect 28353 45917 28365 45920
rect 28399 45917 28411 45951
rect 28353 45911 28411 45917
rect 33134 45908 33140 45960
rect 33192 45908 33198 45960
rect 41874 45908 41880 45960
rect 41932 45948 41938 45960
rect 42153 45951 42211 45957
rect 42153 45948 42165 45951
rect 41932 45920 42165 45948
rect 41932 45908 41938 45920
rect 42153 45917 42165 45920
rect 42199 45917 42211 45951
rect 42153 45911 42211 45917
rect 27632 45852 28212 45880
rect 6733 45815 6791 45821
rect 6733 45781 6745 45815
rect 6779 45812 6791 45815
rect 7466 45812 7472 45824
rect 6779 45784 7472 45812
rect 6779 45781 6791 45784
rect 6733 45775 6791 45781
rect 7466 45772 7472 45784
rect 7524 45772 7530 45824
rect 8846 45772 8852 45824
rect 8904 45812 8910 45824
rect 9309 45815 9367 45821
rect 9309 45812 9321 45815
rect 8904 45784 9321 45812
rect 8904 45772 8910 45784
rect 9309 45781 9321 45784
rect 9355 45781 9367 45815
rect 9309 45775 9367 45781
rect 13998 45772 14004 45824
rect 14056 45812 14062 45824
rect 15105 45815 15163 45821
rect 15105 45812 15117 45815
rect 14056 45784 15117 45812
rect 14056 45772 14062 45784
rect 15105 45781 15117 45784
rect 15151 45781 15163 45815
rect 15105 45775 15163 45781
rect 24121 45815 24179 45821
rect 24121 45781 24133 45815
rect 24167 45812 24179 45815
rect 24946 45812 24952 45824
rect 24167 45784 24952 45812
rect 24167 45781 24179 45784
rect 24121 45775 24179 45781
rect 24946 45772 24952 45784
rect 25004 45772 25010 45824
rect 27522 45772 27528 45824
rect 27580 45772 27586 45824
rect 28184 45821 28212 45852
rect 41966 45840 41972 45892
rect 42024 45840 42030 45892
rect 28169 45815 28227 45821
rect 28169 45781 28181 45815
rect 28215 45812 28227 45815
rect 29086 45812 29092 45824
rect 28215 45784 29092 45812
rect 28215 45781 28227 45784
rect 28169 45775 28227 45781
rect 29086 45772 29092 45784
rect 29144 45772 29150 45824
rect 32030 45772 32036 45824
rect 32088 45812 32094 45824
rect 32953 45815 33011 45821
rect 32953 45812 32965 45815
rect 32088 45784 32965 45812
rect 32088 45772 32094 45784
rect 32953 45781 32965 45784
rect 32999 45781 33011 45815
rect 32953 45775 33011 45781
rect 1104 45722 45172 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 45172 45722
rect 1104 45648 45172 45670
rect 22186 45568 22192 45620
rect 22244 45608 22250 45620
rect 27890 45617 27896 45620
rect 22925 45611 22983 45617
rect 22925 45608 22937 45611
rect 22244 45580 22937 45608
rect 22244 45568 22250 45580
rect 22925 45577 22937 45580
rect 22971 45577 22983 45611
rect 22925 45571 22983 45577
rect 27709 45611 27767 45617
rect 27709 45577 27721 45611
rect 27755 45608 27767 45611
rect 27877 45611 27896 45617
rect 27755 45580 27789 45608
rect 27755 45577 27767 45580
rect 27709 45571 27767 45577
rect 27877 45577 27889 45611
rect 27877 45571 27896 45577
rect 9493 45543 9551 45549
rect 9493 45509 9505 45543
rect 9539 45540 9551 45543
rect 10042 45540 10048 45552
rect 9539 45512 10048 45540
rect 9539 45509 9551 45512
rect 9493 45503 9551 45509
rect 10042 45500 10048 45512
rect 10100 45500 10106 45552
rect 13722 45540 13728 45552
rect 13280 45512 13728 45540
rect 8849 45475 8907 45481
rect 8849 45441 8861 45475
rect 8895 45472 8907 45475
rect 9585 45475 9643 45481
rect 8895 45444 9168 45472
rect 8895 45441 8907 45444
rect 8849 45435 8907 45441
rect 9140 45345 9168 45444
rect 9585 45441 9597 45475
rect 9631 45472 9643 45475
rect 10134 45472 10140 45484
rect 9631 45444 10140 45472
rect 9631 45441 9643 45444
rect 9585 45435 9643 45441
rect 10134 45432 10140 45444
rect 10192 45472 10198 45484
rect 10597 45475 10655 45481
rect 10597 45472 10609 45475
rect 10192 45444 10609 45472
rect 10192 45432 10198 45444
rect 10597 45441 10609 45444
rect 10643 45441 10655 45475
rect 10597 45435 10655 45441
rect 11698 45432 11704 45484
rect 11756 45432 11762 45484
rect 13280 45481 13308 45512
rect 13722 45500 13728 45512
rect 13780 45500 13786 45552
rect 15841 45543 15899 45549
rect 15841 45509 15853 45543
rect 15887 45540 15899 45543
rect 15930 45540 15936 45552
rect 15887 45512 15936 45540
rect 15887 45509 15899 45512
rect 15841 45503 15899 45509
rect 15930 45500 15936 45512
rect 15988 45540 15994 45552
rect 16298 45540 16304 45552
rect 15988 45512 16304 45540
rect 15988 45500 15994 45512
rect 16298 45500 16304 45512
rect 16356 45500 16362 45552
rect 16482 45500 16488 45552
rect 16540 45540 16546 45552
rect 25409 45543 25467 45549
rect 25409 45540 25421 45543
rect 16540 45512 17264 45540
rect 16540 45500 16546 45512
rect 13538 45481 13544 45484
rect 13265 45475 13323 45481
rect 13265 45441 13277 45475
rect 13311 45441 13323 45475
rect 13265 45435 13323 45441
rect 13532 45435 13544 45481
rect 13538 45432 13544 45435
rect 13596 45432 13602 45484
rect 16025 45475 16083 45481
rect 16025 45441 16037 45475
rect 16071 45472 16083 45475
rect 16071 45444 16712 45472
rect 16071 45441 16083 45444
rect 16025 45435 16083 45441
rect 9769 45407 9827 45413
rect 9769 45373 9781 45407
rect 9815 45373 9827 45407
rect 9769 45367 9827 45373
rect 9125 45339 9183 45345
rect 9125 45305 9137 45339
rect 9171 45305 9183 45339
rect 9784 45336 9812 45367
rect 9950 45364 9956 45416
rect 10008 45364 10014 45416
rect 12526 45364 12532 45416
rect 12584 45364 12590 45416
rect 15289 45407 15347 45413
rect 15289 45404 15301 45407
rect 14660 45376 15301 45404
rect 12544 45336 12572 45364
rect 14660 45345 14688 45376
rect 15289 45373 15301 45376
rect 15335 45373 15347 45407
rect 15289 45367 15347 45373
rect 9784 45308 12572 45336
rect 14645 45339 14703 45345
rect 9125 45299 9183 45305
rect 14645 45305 14657 45339
rect 14691 45305 14703 45339
rect 16574 45336 16580 45348
rect 14645 45299 14703 45305
rect 15764 45308 16580 45336
rect 9030 45228 9036 45280
rect 9088 45228 9094 45280
rect 11514 45228 11520 45280
rect 11572 45228 11578 45280
rect 14734 45228 14740 45280
rect 14792 45228 14798 45280
rect 15764 45277 15792 45308
rect 16574 45296 16580 45308
rect 16632 45296 16638 45348
rect 16684 45345 16712 45444
rect 16850 45432 16856 45484
rect 16908 45472 16914 45484
rect 17037 45475 17095 45481
rect 17037 45472 17049 45475
rect 16908 45444 17049 45472
rect 16908 45432 16914 45444
rect 17037 45441 17049 45444
rect 17083 45441 17095 45475
rect 17037 45435 17095 45441
rect 17236 45413 17264 45512
rect 23400 45512 25421 45540
rect 23400 45484 23428 45512
rect 25409 45509 25421 45512
rect 25455 45509 25467 45543
rect 25409 45503 25467 45509
rect 25866 45500 25872 45552
rect 25924 45540 25930 45552
rect 27724 45540 27752 45571
rect 27890 45568 27896 45571
rect 27948 45568 27954 45620
rect 25924 45512 27752 45540
rect 25924 45500 25930 45512
rect 28074 45500 28080 45552
rect 28132 45500 28138 45552
rect 18414 45432 18420 45484
rect 18472 45432 18478 45484
rect 22002 45432 22008 45484
rect 22060 45432 22066 45484
rect 23382 45432 23388 45484
rect 23440 45432 23446 45484
rect 23934 45432 23940 45484
rect 23992 45472 23998 45484
rect 24029 45475 24087 45481
rect 24029 45472 24041 45475
rect 23992 45444 24041 45472
rect 23992 45432 23998 45444
rect 24029 45441 24041 45444
rect 24075 45441 24087 45475
rect 24029 45435 24087 45441
rect 24118 45432 24124 45484
rect 24176 45472 24182 45484
rect 24213 45475 24271 45481
rect 24213 45472 24225 45475
rect 24176 45444 24225 45472
rect 24176 45432 24182 45444
rect 24213 45441 24225 45444
rect 24259 45441 24271 45475
rect 24213 45435 24271 45441
rect 25133 45475 25191 45481
rect 25133 45441 25145 45475
rect 25179 45441 25191 45475
rect 25133 45435 25191 45441
rect 17129 45407 17187 45413
rect 17129 45404 17141 45407
rect 17052 45376 17141 45404
rect 16669 45339 16727 45345
rect 16669 45305 16681 45339
rect 16715 45305 16727 45339
rect 16669 45299 16727 45305
rect 17052 45280 17080 45376
rect 17129 45373 17141 45376
rect 17175 45373 17187 45407
rect 17129 45367 17187 45373
rect 17221 45407 17279 45413
rect 17221 45373 17233 45407
rect 17267 45373 17279 45407
rect 17221 45367 17279 45373
rect 17310 45364 17316 45416
rect 17368 45404 17374 45416
rect 18049 45407 18107 45413
rect 18049 45404 18061 45407
rect 17368 45376 18061 45404
rect 17368 45364 17374 45376
rect 18049 45373 18061 45376
rect 18095 45373 18107 45407
rect 18049 45367 18107 45373
rect 23474 45364 23480 45416
rect 23532 45364 23538 45416
rect 25148 45404 25176 45435
rect 28534 45432 28540 45484
rect 28592 45432 28598 45484
rect 25148 45376 25544 45404
rect 25516 45280 25544 45376
rect 26694 45364 26700 45416
rect 26752 45404 26758 45416
rect 27525 45407 27583 45413
rect 27525 45404 27537 45407
rect 26752 45376 27537 45404
rect 26752 45364 26758 45376
rect 27525 45373 27537 45376
rect 27571 45373 27583 45407
rect 27525 45367 27583 45373
rect 29638 45364 29644 45416
rect 29696 45364 29702 45416
rect 29914 45364 29920 45416
rect 29972 45364 29978 45416
rect 30561 45407 30619 45413
rect 30561 45373 30573 45407
rect 30607 45373 30619 45407
rect 30561 45367 30619 45373
rect 30576 45336 30604 45367
rect 29840 45308 30604 45336
rect 15749 45271 15807 45277
rect 15749 45237 15761 45271
rect 15795 45237 15807 45271
rect 15749 45231 15807 45237
rect 16206 45228 16212 45280
rect 16264 45228 16270 45280
rect 17034 45228 17040 45280
rect 17092 45268 17098 45280
rect 17497 45271 17555 45277
rect 17497 45268 17509 45271
rect 17092 45240 17509 45268
rect 17092 45228 17098 45240
rect 17497 45237 17509 45240
rect 17543 45237 17555 45271
rect 17497 45231 17555 45237
rect 18230 45228 18236 45280
rect 18288 45228 18294 45280
rect 22370 45228 22376 45280
rect 22428 45268 22434 45280
rect 22649 45271 22707 45277
rect 22649 45268 22661 45271
rect 22428 45240 22661 45268
rect 22428 45228 22434 45240
rect 22649 45237 22661 45240
rect 22695 45237 22707 45271
rect 22649 45231 22707 45237
rect 24026 45228 24032 45280
rect 24084 45228 24090 45280
rect 25041 45271 25099 45277
rect 25041 45237 25053 45271
rect 25087 45268 25099 45271
rect 25130 45268 25136 45280
rect 25087 45240 25136 45268
rect 25087 45237 25099 45240
rect 25041 45231 25099 45237
rect 25130 45228 25136 45240
rect 25188 45228 25194 45280
rect 25498 45228 25504 45280
rect 25556 45228 25562 45280
rect 26418 45228 26424 45280
rect 26476 45268 26482 45280
rect 26973 45271 27031 45277
rect 26973 45268 26985 45271
rect 26476 45240 26985 45268
rect 26476 45228 26482 45240
rect 26973 45237 26985 45240
rect 27019 45237 27031 45271
rect 26973 45231 27031 45237
rect 27154 45228 27160 45280
rect 27212 45268 27218 45280
rect 27893 45271 27951 45277
rect 27893 45268 27905 45271
rect 27212 45240 27905 45268
rect 27212 45228 27218 45240
rect 27893 45237 27905 45240
rect 27939 45268 27951 45271
rect 28169 45271 28227 45277
rect 28169 45268 28181 45271
rect 27939 45240 28181 45268
rect 27939 45237 27951 45240
rect 27893 45231 27951 45237
rect 28169 45237 28181 45240
rect 28215 45268 28227 45271
rect 29840 45268 29868 45308
rect 28215 45240 29868 45268
rect 28215 45237 28227 45240
rect 28169 45231 28227 45237
rect 30006 45228 30012 45280
rect 30064 45228 30070 45280
rect 1104 45178 45172 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 45172 45178
rect 1104 45104 45172 45126
rect 9030 45024 9036 45076
rect 9088 45064 9094 45076
rect 9198 45067 9256 45073
rect 9198 45064 9210 45067
rect 9088 45036 9210 45064
rect 9088 45024 9094 45036
rect 9198 45033 9210 45036
rect 9244 45033 9256 45067
rect 9198 45027 9256 45033
rect 11320 45067 11378 45073
rect 11320 45033 11332 45067
rect 11366 45064 11378 45067
rect 11514 45064 11520 45076
rect 11366 45036 11520 45064
rect 11366 45033 11378 45036
rect 11320 45027 11378 45033
rect 11514 45024 11520 45036
rect 11572 45024 11578 45076
rect 13538 45024 13544 45076
rect 13596 45064 13602 45076
rect 13633 45067 13691 45073
rect 13633 45064 13645 45067
rect 13596 45036 13645 45064
rect 13596 45024 13602 45036
rect 13633 45033 13645 45036
rect 13679 45033 13691 45067
rect 13633 45027 13691 45033
rect 14292 45036 15332 45064
rect 8938 44888 8944 44940
rect 8996 44928 9002 44940
rect 11057 44931 11115 44937
rect 11057 44928 11069 44931
rect 8996 44900 11069 44928
rect 8996 44888 9002 44900
rect 11057 44897 11069 44900
rect 11103 44928 11115 44931
rect 11974 44928 11980 44940
rect 11103 44900 11980 44928
rect 11103 44897 11115 44900
rect 11057 44891 11115 44897
rect 11974 44888 11980 44900
rect 12032 44888 12038 44940
rect 12805 44931 12863 44937
rect 12805 44897 12817 44931
rect 12851 44928 12863 44931
rect 12894 44928 12900 44940
rect 12851 44900 12900 44928
rect 12851 44897 12863 44900
rect 12805 44891 12863 44897
rect 12894 44888 12900 44900
rect 12952 44928 12958 44940
rect 14292 44937 14320 45036
rect 14458 44956 14464 45008
rect 14516 44996 14522 45008
rect 14921 44999 14979 45005
rect 14921 44996 14933 44999
rect 14516 44968 14933 44996
rect 14516 44956 14522 44968
rect 14921 44965 14933 44968
rect 14967 44965 14979 44999
rect 14921 44959 14979 44965
rect 15304 44940 15332 45036
rect 16298 45024 16304 45076
rect 16356 45064 16362 45076
rect 17576 45067 17634 45073
rect 16356 45036 17448 45064
rect 16356 45024 16362 45036
rect 13449 44931 13507 44937
rect 13449 44928 13461 44931
rect 12952 44900 13461 44928
rect 12952 44888 12958 44900
rect 13449 44897 13461 44900
rect 13495 44897 13507 44931
rect 13449 44891 13507 44897
rect 14277 44931 14335 44937
rect 14277 44897 14289 44931
rect 14323 44897 14335 44931
rect 14277 44891 14335 44897
rect 14369 44931 14427 44937
rect 14369 44897 14381 44931
rect 14415 44928 14427 44931
rect 14734 44928 14740 44940
rect 14415 44900 14740 44928
rect 14415 44897 14427 44900
rect 14369 44891 14427 44897
rect 14734 44888 14740 44900
rect 14792 44888 14798 44940
rect 15286 44888 15292 44940
rect 15344 44888 15350 44940
rect 16206 44888 16212 44940
rect 16264 44928 16270 44940
rect 16945 44931 17003 44937
rect 16945 44928 16957 44931
rect 16264 44900 16957 44928
rect 16264 44888 16270 44900
rect 16945 44897 16957 44900
rect 16991 44897 17003 44931
rect 17420 44928 17448 45036
rect 17576 45033 17588 45067
rect 17622 45064 17634 45067
rect 18230 45064 18236 45076
rect 17622 45036 18236 45064
rect 17622 45033 17634 45036
rect 17576 45027 17634 45033
rect 18230 45024 18236 45036
rect 18288 45024 18294 45076
rect 24026 45024 24032 45076
rect 24084 45024 24090 45076
rect 27985 45067 28043 45073
rect 27985 45033 27997 45067
rect 28031 45064 28043 45067
rect 28074 45064 28080 45076
rect 28031 45036 28080 45064
rect 28031 45033 28043 45036
rect 27985 45027 28043 45033
rect 28074 45024 28080 45036
rect 28132 45024 28138 45076
rect 29365 45067 29423 45073
rect 29365 45033 29377 45067
rect 29411 45064 29423 45067
rect 29638 45064 29644 45076
rect 29411 45036 29644 45064
rect 29411 45033 29423 45036
rect 29365 45027 29423 45033
rect 29638 45024 29644 45036
rect 29696 45024 29702 45076
rect 30006 45024 30012 45076
rect 30064 45024 30070 45076
rect 23566 44956 23572 45008
rect 23624 44996 23630 45008
rect 23937 44999 23995 45005
rect 23937 44996 23949 44999
rect 23624 44968 23949 44996
rect 23624 44956 23630 44968
rect 23937 44965 23949 44968
rect 23983 44965 23995 44999
rect 23937 44959 23995 44965
rect 21637 44931 21695 44937
rect 17420 44900 18828 44928
rect 16945 44891 17003 44897
rect 8757 44863 8815 44869
rect 8757 44829 8769 44863
rect 8803 44860 8815 44863
rect 8846 44860 8852 44872
rect 8803 44832 8852 44860
rect 8803 44829 8815 44832
rect 8757 44823 8815 44829
rect 8846 44820 8852 44832
rect 8904 44820 8910 44872
rect 13814 44820 13820 44872
rect 13872 44820 13878 44872
rect 15105 44863 15163 44869
rect 15105 44860 15117 44863
rect 14844 44832 15117 44860
rect 10502 44792 10508 44804
rect 10442 44764 10508 44792
rect 10502 44752 10508 44764
rect 10560 44792 10566 44804
rect 10560 44764 11822 44792
rect 10560 44752 10566 44764
rect 8570 44684 8576 44736
rect 8628 44684 8634 44736
rect 10042 44684 10048 44736
rect 10100 44724 10106 44736
rect 10689 44727 10747 44733
rect 10689 44724 10701 44727
rect 10100 44696 10701 44724
rect 10100 44684 10106 44696
rect 10689 44693 10701 44696
rect 10735 44693 10747 44727
rect 10689 44687 10747 44693
rect 12158 44684 12164 44736
rect 12216 44724 12222 44736
rect 12897 44727 12955 44733
rect 12897 44724 12909 44727
rect 12216 44696 12909 44724
rect 12216 44684 12222 44696
rect 12897 44693 12909 44696
rect 12943 44693 12955 44727
rect 12897 44687 12955 44693
rect 13262 44684 13268 44736
rect 13320 44724 13326 44736
rect 14844 44733 14872 44832
rect 15105 44829 15117 44832
rect 15151 44829 15163 44863
rect 15105 44823 15163 44829
rect 17221 44863 17279 44869
rect 17221 44829 17233 44863
rect 17267 44860 17279 44863
rect 17313 44863 17371 44869
rect 17313 44860 17325 44863
rect 17267 44832 17325 44860
rect 17267 44829 17279 44832
rect 17221 44823 17279 44829
rect 17313 44829 17325 44832
rect 17359 44829 17371 44863
rect 17313 44823 17371 44829
rect 16666 44792 16672 44804
rect 16514 44764 16672 44792
rect 16666 44752 16672 44764
rect 16724 44752 16730 44804
rect 17328 44792 17356 44823
rect 17862 44792 17868 44804
rect 17328 44764 17868 44792
rect 17862 44752 17868 44764
rect 17920 44752 17926 44804
rect 18800 44792 18828 44900
rect 21637 44897 21649 44931
rect 21683 44928 21695 44931
rect 22186 44928 22192 44940
rect 21683 44900 22192 44928
rect 21683 44897 21695 44900
rect 21637 44891 21695 44897
rect 22186 44888 22192 44900
rect 22244 44888 22250 44940
rect 23109 44931 23167 44937
rect 23109 44897 23121 44931
rect 23155 44928 23167 44931
rect 24044 44928 24072 45024
rect 24673 44931 24731 44937
rect 24673 44928 24685 44931
rect 23155 44900 23336 44928
rect 24044 44900 24685 44928
rect 23155 44897 23167 44900
rect 23109 44891 23167 44897
rect 21174 44820 21180 44872
rect 21232 44860 21238 44872
rect 23308 44869 23336 44900
rect 24673 44897 24685 44900
rect 24719 44897 24731 44931
rect 28092 44928 28120 45024
rect 28629 44931 28687 44937
rect 28629 44928 28641 44931
rect 28092 44900 28641 44928
rect 24673 44891 24731 44897
rect 28629 44897 28641 44900
rect 28675 44897 28687 44931
rect 28629 44891 28687 44897
rect 29086 44888 29092 44940
rect 29144 44888 29150 44940
rect 21361 44863 21419 44869
rect 21361 44860 21373 44863
rect 21232 44832 21373 44860
rect 21232 44820 21238 44832
rect 21361 44829 21373 44832
rect 21407 44829 21419 44863
rect 21361 44823 21419 44829
rect 23293 44863 23351 44869
rect 23293 44829 23305 44863
rect 23339 44860 23351 44863
rect 23658 44860 23664 44872
rect 23339 44832 23664 44860
rect 23339 44829 23351 44832
rect 23293 44823 23351 44829
rect 23658 44820 23664 44832
rect 23716 44820 23722 44872
rect 24118 44860 24124 44872
rect 23768 44832 24124 44860
rect 23768 44804 23796 44832
rect 24118 44820 24124 44832
rect 24176 44860 24182 44872
rect 24213 44863 24271 44869
rect 24213 44860 24225 44863
rect 24176 44832 24225 44860
rect 24176 44820 24182 44832
rect 24213 44829 24225 44832
rect 24259 44829 24271 44863
rect 24213 44823 24271 44829
rect 24394 44820 24400 44872
rect 24452 44820 24458 44872
rect 26234 44820 26240 44872
rect 26292 44820 26298 44872
rect 28997 44863 29055 44869
rect 28997 44829 29009 44863
rect 29043 44860 29055 44863
rect 30024 44860 30052 45024
rect 29043 44832 30052 44860
rect 29043 44829 29055 44832
rect 28997 44823 29055 44829
rect 20622 44792 20628 44804
rect 18800 44778 20628 44792
rect 18814 44764 20628 44778
rect 20622 44752 20628 44764
rect 20680 44752 20686 44804
rect 22646 44752 22652 44804
rect 22704 44752 22710 44804
rect 23750 44752 23756 44804
rect 23808 44752 23814 44804
rect 23845 44795 23903 44801
rect 23845 44761 23857 44795
rect 23891 44792 23903 44795
rect 23937 44795 23995 44801
rect 23937 44792 23949 44795
rect 23891 44764 23949 44792
rect 23891 44761 23903 44764
rect 23845 44755 23903 44761
rect 23937 44761 23949 44764
rect 23983 44761 23995 44795
rect 23937 44755 23995 44761
rect 25130 44752 25136 44804
rect 25188 44752 25194 44804
rect 26510 44752 26516 44804
rect 26568 44752 26574 44804
rect 28534 44792 28540 44804
rect 27738 44764 28540 44792
rect 28534 44752 28540 44764
rect 28592 44752 28598 44804
rect 14461 44727 14519 44733
rect 14461 44724 14473 44727
rect 13320 44696 14473 44724
rect 13320 44684 13326 44696
rect 14461 44693 14473 44696
rect 14507 44693 14519 44727
rect 14461 44687 14519 44693
rect 14829 44727 14887 44733
rect 14829 44693 14841 44727
rect 14875 44693 14887 44727
rect 14829 44687 14887 44693
rect 15473 44727 15531 44733
rect 15473 44693 15485 44727
rect 15519 44724 15531 44727
rect 16850 44724 16856 44736
rect 15519 44696 16856 44724
rect 15519 44693 15531 44696
rect 15473 44687 15531 44693
rect 16850 44684 16856 44696
rect 16908 44684 16914 44736
rect 19058 44684 19064 44736
rect 19116 44684 19122 44736
rect 23474 44684 23480 44736
rect 23532 44724 23538 44736
rect 24121 44727 24179 44733
rect 24121 44724 24133 44727
rect 23532 44696 24133 44724
rect 23532 44684 23538 44696
rect 24121 44693 24133 44696
rect 24167 44693 24179 44727
rect 24121 44687 24179 44693
rect 25682 44684 25688 44736
rect 25740 44724 25746 44736
rect 26145 44727 26203 44733
rect 26145 44724 26157 44727
rect 25740 44696 26157 44724
rect 25740 44684 25746 44696
rect 26145 44693 26157 44696
rect 26191 44693 26203 44727
rect 26145 44687 26203 44693
rect 28074 44684 28080 44736
rect 28132 44684 28138 44736
rect 1104 44634 45172 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 45172 44634
rect 1104 44560 45172 44582
rect 8938 44480 8944 44532
rect 8996 44480 9002 44532
rect 9677 44523 9735 44529
rect 9677 44489 9689 44523
rect 9723 44489 9735 44523
rect 9677 44483 9735 44489
rect 9769 44523 9827 44529
rect 9769 44489 9781 44523
rect 9815 44520 9827 44523
rect 9858 44520 9864 44532
rect 9815 44492 9864 44520
rect 9815 44489 9827 44492
rect 9769 44483 9827 44489
rect 8956 44452 8984 44480
rect 8312 44424 8984 44452
rect 9692 44452 9720 44483
rect 9858 44480 9864 44492
rect 9916 44480 9922 44532
rect 9950 44480 9956 44532
rect 10008 44480 10014 44532
rect 10134 44480 10140 44532
rect 10192 44480 10198 44532
rect 10965 44523 11023 44529
rect 10965 44520 10977 44523
rect 10796 44492 10977 44520
rect 9968 44452 9996 44480
rect 9692 44424 9996 44452
rect 8312 44393 8340 44424
rect 8570 44393 8576 44396
rect 8297 44387 8355 44393
rect 8297 44353 8309 44387
rect 8343 44353 8355 44387
rect 8564 44384 8576 44393
rect 8531 44356 8576 44384
rect 8297 44347 8355 44353
rect 8564 44347 8576 44356
rect 8570 44344 8576 44347
rect 8628 44344 8634 44396
rect 10686 44344 10692 44396
rect 10744 44384 10750 44396
rect 10796 44384 10824 44492
rect 10965 44489 10977 44492
rect 11011 44489 11023 44523
rect 10965 44483 11023 44489
rect 11333 44523 11391 44529
rect 11333 44489 11345 44523
rect 11379 44489 11391 44523
rect 11333 44483 11391 44489
rect 11609 44523 11667 44529
rect 11609 44489 11621 44523
rect 11655 44520 11667 44523
rect 11698 44520 11704 44532
rect 11655 44492 11704 44520
rect 11655 44489 11667 44492
rect 11609 44483 11667 44489
rect 10873 44455 10931 44461
rect 10873 44421 10885 44455
rect 10919 44452 10931 44455
rect 11238 44452 11244 44464
rect 10919 44424 11244 44452
rect 10919 44421 10931 44424
rect 10873 44415 10931 44421
rect 11238 44412 11244 44424
rect 11296 44412 11302 44464
rect 11348 44384 11376 44483
rect 11698 44480 11704 44492
rect 11756 44480 11762 44532
rect 11977 44523 12035 44529
rect 11977 44489 11989 44523
rect 12023 44520 12035 44523
rect 12158 44520 12164 44532
rect 12023 44492 12164 44520
rect 12023 44489 12035 44492
rect 11977 44483 12035 44489
rect 12158 44480 12164 44492
rect 12216 44480 12222 44532
rect 12894 44480 12900 44532
rect 12952 44480 12958 44532
rect 14642 44480 14648 44532
rect 14700 44520 14706 44532
rect 14826 44520 14832 44532
rect 14700 44492 14832 44520
rect 14700 44480 14706 44492
rect 14826 44480 14832 44492
rect 14884 44480 14890 44532
rect 16485 44523 16543 44529
rect 16485 44489 16497 44523
rect 16531 44489 16543 44523
rect 16485 44483 16543 44489
rect 12912 44393 12940 44480
rect 16500 44452 16528 44483
rect 17034 44480 17040 44532
rect 17092 44480 17098 44532
rect 17310 44480 17316 44532
rect 17368 44480 17374 44532
rect 18233 44523 18291 44529
rect 18233 44489 18245 44523
rect 18279 44489 18291 44523
rect 18233 44483 18291 44489
rect 17328 44452 17356 44480
rect 14030 44424 15516 44452
rect 16500 44424 17356 44452
rect 18248 44452 18276 44483
rect 22370 44480 22376 44532
rect 22428 44480 22434 44532
rect 23474 44480 23480 44532
rect 23532 44520 23538 44532
rect 23569 44523 23627 44529
rect 23569 44520 23581 44523
rect 23532 44492 23581 44520
rect 23532 44480 23538 44492
rect 23569 44489 23581 44492
rect 23615 44489 23627 44523
rect 23569 44483 23627 44489
rect 23845 44523 23903 44529
rect 23845 44489 23857 44523
rect 23891 44520 23903 44523
rect 23934 44520 23940 44532
rect 23891 44492 23940 44520
rect 23891 44489 23903 44492
rect 23845 44483 23903 44489
rect 23934 44480 23940 44492
rect 23992 44480 23998 44532
rect 24210 44480 24216 44532
rect 24268 44520 24274 44532
rect 25409 44523 25467 44529
rect 25409 44520 25421 44523
rect 24268 44492 25421 44520
rect 24268 44480 24274 44492
rect 25409 44489 25421 44492
rect 25455 44489 25467 44523
rect 25409 44483 25467 44489
rect 25961 44523 26019 44529
rect 25961 44489 25973 44523
rect 26007 44520 26019 44523
rect 26510 44520 26516 44532
rect 26007 44492 26516 44520
rect 26007 44489 26019 44492
rect 25961 44483 26019 44489
rect 26510 44480 26516 44492
rect 26568 44480 26574 44532
rect 26694 44529 26700 44532
rect 26690 44520 26700 44529
rect 26655 44492 26700 44520
rect 26690 44483 26700 44492
rect 26694 44480 26700 44483
rect 26752 44480 26758 44532
rect 28074 44520 28080 44532
rect 26804 44492 28080 44520
rect 18570 44455 18628 44461
rect 18570 44452 18582 44455
rect 18248 44424 18582 44452
rect 15378 44393 15384 44396
rect 12621 44387 12679 44393
rect 12621 44384 12633 44387
rect 10744 44356 11192 44384
rect 11348 44356 12633 44384
rect 10744 44344 10750 44356
rect 9306 44276 9312 44328
rect 9364 44316 9370 44328
rect 10229 44319 10287 44325
rect 10229 44316 10241 44319
rect 9364 44288 10241 44316
rect 9364 44276 9370 44288
rect 10229 44285 10241 44288
rect 10275 44285 10287 44319
rect 10229 44279 10287 44285
rect 10413 44319 10471 44325
rect 10413 44285 10425 44319
rect 10459 44316 10471 44319
rect 10781 44319 10839 44325
rect 10781 44316 10793 44319
rect 10459 44288 10793 44316
rect 10459 44285 10471 44288
rect 10413 44279 10471 44285
rect 10781 44285 10793 44288
rect 10827 44285 10839 44319
rect 11164 44316 11192 44356
rect 12621 44353 12633 44356
rect 12667 44353 12679 44387
rect 12621 44347 12679 44353
rect 12897 44387 12955 44393
rect 12897 44353 12909 44387
rect 12943 44353 12955 44387
rect 12897 44347 12955 44353
rect 13004 44356 13308 44384
rect 12069 44319 12127 44325
rect 12069 44316 12081 44319
rect 11164 44288 12081 44316
rect 10781 44279 10839 44285
rect 12069 44285 12081 44288
rect 12115 44285 12127 44319
rect 12069 44279 12127 44285
rect 12253 44319 12311 44325
rect 12253 44285 12265 44319
rect 12299 44316 12311 44319
rect 12526 44316 12532 44328
rect 12299 44288 12532 44316
rect 12299 44285 12311 44288
rect 12253 44279 12311 44285
rect 10502 44208 10508 44260
rect 10560 44208 10566 44260
rect 10796 44248 10824 44279
rect 12526 44276 12532 44288
rect 12584 44276 12590 44328
rect 12805 44319 12863 44325
rect 12805 44285 12817 44319
rect 12851 44316 12863 44319
rect 13004 44316 13032 44356
rect 12851 44288 13032 44316
rect 12851 44285 12863 44288
rect 12805 44279 12863 44285
rect 13170 44276 13176 44328
rect 13228 44276 13234 44328
rect 13280 44316 13308 44356
rect 15372 44347 15384 44393
rect 15378 44344 15384 44347
rect 15436 44344 15442 44396
rect 15488 44384 15516 44424
rect 18570 44421 18582 44424
rect 18616 44421 18628 44455
rect 18570 44415 18628 44421
rect 22097 44455 22155 44461
rect 22097 44421 22109 44455
rect 22143 44452 22155 44455
rect 22388 44452 22416 44480
rect 22143 44424 22416 44452
rect 22143 44421 22155 44424
rect 22097 44415 22155 44421
rect 22646 44412 22652 44464
rect 22704 44412 22710 44464
rect 24121 44455 24179 44461
rect 24121 44452 24133 44455
rect 23768 44424 24133 44452
rect 16666 44384 16672 44396
rect 15488 44356 16672 44384
rect 16666 44344 16672 44356
rect 16724 44384 16730 44396
rect 17494 44384 17500 44396
rect 16724 44356 17500 44384
rect 16724 44344 16730 44356
rect 17494 44344 17500 44356
rect 17552 44344 17558 44396
rect 18049 44387 18107 44393
rect 18049 44353 18061 44387
rect 18095 44384 18107 44387
rect 18874 44384 18880 44396
rect 18095 44356 18880 44384
rect 18095 44353 18107 44356
rect 18049 44347 18107 44353
rect 18874 44344 18880 44356
rect 18932 44344 18938 44396
rect 23768 44393 23796 44424
rect 24121 44421 24133 44424
rect 24167 44421 24179 44455
rect 24121 44415 24179 44421
rect 24857 44455 24915 44461
rect 24857 44421 24869 44455
rect 24903 44452 24915 44455
rect 26418 44452 26424 44464
rect 24903 44424 26004 44452
rect 24903 44421 24915 44424
rect 24857 44415 24915 44421
rect 23753 44387 23811 44393
rect 19536 44356 20484 44384
rect 13446 44316 13452 44328
rect 13280 44288 13452 44316
rect 13446 44276 13452 44288
rect 13504 44276 13510 44328
rect 14458 44276 14464 44328
rect 14516 44276 14522 44328
rect 14737 44319 14795 44325
rect 14737 44285 14749 44319
rect 14783 44316 14795 44319
rect 15105 44319 15163 44325
rect 15105 44316 15117 44319
rect 14783 44288 15117 44316
rect 14783 44285 14795 44288
rect 14737 44279 14795 44285
rect 15105 44285 15117 44288
rect 15151 44285 15163 44319
rect 15105 44279 15163 44285
rect 13188 44248 13216 44276
rect 10796 44220 13216 44248
rect 8202 44140 8208 44192
rect 8260 44180 8266 44192
rect 10520 44180 10548 44208
rect 8260 44152 10548 44180
rect 8260 44140 8266 44152
rect 12434 44140 12440 44192
rect 12492 44140 12498 44192
rect 12989 44183 13047 44189
rect 12989 44149 13001 44183
rect 13035 44180 13047 44183
rect 13262 44180 13268 44192
rect 13035 44152 13268 44180
rect 13035 44149 13047 44152
rect 12989 44143 13047 44149
rect 13262 44140 13268 44152
rect 13320 44140 13326 44192
rect 13722 44140 13728 44192
rect 13780 44180 13786 44192
rect 14752 44180 14780 44279
rect 17126 44276 17132 44328
rect 17184 44276 17190 44328
rect 17310 44276 17316 44328
rect 17368 44276 17374 44328
rect 18325 44319 18383 44325
rect 18325 44285 18337 44319
rect 18371 44285 18383 44319
rect 18325 44279 18383 44285
rect 14826 44208 14832 44260
rect 14884 44208 14890 44260
rect 16546 44220 16804 44248
rect 13780 44152 14780 44180
rect 14844 44180 14872 44208
rect 16546 44180 16574 44220
rect 14844 44152 16574 44180
rect 13780 44140 13786 44152
rect 16666 44140 16672 44192
rect 16724 44140 16730 44192
rect 16776 44180 16804 44220
rect 18046 44208 18052 44260
rect 18104 44248 18110 44260
rect 18340 44248 18368 44279
rect 18104 44220 18368 44248
rect 18104 44208 18110 44220
rect 19536 44180 19564 44356
rect 20349 44319 20407 44325
rect 20349 44285 20361 44319
rect 20395 44285 20407 44319
rect 20349 44279 20407 44285
rect 19705 44251 19763 44257
rect 19705 44217 19717 44251
rect 19751 44248 19763 44251
rect 20364 44248 20392 44279
rect 19751 44220 20392 44248
rect 19751 44217 19763 44220
rect 19705 44211 19763 44217
rect 16776 44152 19564 44180
rect 19610 44140 19616 44192
rect 19668 44180 19674 44192
rect 19797 44183 19855 44189
rect 19797 44180 19809 44183
rect 19668 44152 19809 44180
rect 19668 44140 19674 44152
rect 19797 44149 19809 44152
rect 19843 44149 19855 44183
rect 20456 44180 20484 44356
rect 23753 44353 23765 44387
rect 23799 44353 23811 44387
rect 23753 44347 23811 44353
rect 23937 44387 23995 44393
rect 23937 44353 23949 44387
rect 23983 44384 23995 44387
rect 25593 44387 25651 44393
rect 25593 44384 25605 44387
rect 23983 44356 25605 44384
rect 23983 44353 23995 44356
rect 23937 44347 23995 44353
rect 25593 44353 25605 44356
rect 25639 44384 25651 44387
rect 25866 44384 25872 44396
rect 25639 44356 25872 44384
rect 25639 44353 25651 44356
rect 25593 44347 25651 44353
rect 25866 44344 25872 44356
rect 25924 44344 25930 44396
rect 21174 44276 21180 44328
rect 21232 44316 21238 44328
rect 21821 44319 21879 44325
rect 21821 44316 21833 44319
rect 21232 44288 21833 44316
rect 21232 44276 21238 44288
rect 21821 44285 21833 44288
rect 21867 44285 21879 44319
rect 21821 44279 21879 44285
rect 24765 44319 24823 44325
rect 24765 44285 24777 44319
rect 24811 44316 24823 44319
rect 25682 44316 25688 44328
rect 24811 44288 25688 44316
rect 24811 44285 24823 44288
rect 24765 44279 24823 44285
rect 25682 44276 25688 44288
rect 25740 44316 25746 44328
rect 25777 44319 25835 44325
rect 25777 44316 25789 44319
rect 25740 44288 25789 44316
rect 25740 44276 25746 44288
rect 25777 44285 25789 44288
rect 25823 44285 25835 44319
rect 25777 44279 25835 44285
rect 25130 44208 25136 44260
rect 25188 44208 25194 44260
rect 25976 44248 26004 44424
rect 26206 44424 26424 44452
rect 26053 44387 26111 44393
rect 26053 44353 26065 44387
rect 26099 44384 26111 44387
rect 26206 44384 26234 44424
rect 26418 44412 26424 44424
rect 26476 44412 26482 44464
rect 26804 44461 26832 44492
rect 28074 44480 28080 44492
rect 28132 44480 28138 44532
rect 26789 44455 26847 44461
rect 26789 44421 26801 44455
rect 26835 44421 26847 44455
rect 27154 44452 27160 44464
rect 26789 44415 26847 44421
rect 26988 44424 27160 44452
rect 26099 44356 26234 44384
rect 26099 44353 26111 44356
rect 26053 44347 26111 44353
rect 26510 44344 26516 44396
rect 26568 44344 26574 44396
rect 26605 44387 26663 44393
rect 26605 44353 26617 44387
rect 26651 44384 26663 44387
rect 26988 44384 27016 44424
rect 27154 44412 27160 44424
rect 27212 44412 27218 44464
rect 27249 44455 27307 44461
rect 27249 44421 27261 44455
rect 27295 44452 27307 44455
rect 27522 44452 27528 44464
rect 27295 44424 27528 44452
rect 27295 44421 27307 44424
rect 27249 44415 27307 44421
rect 27522 44412 27528 44424
rect 27580 44412 27586 44464
rect 28534 44384 28540 44396
rect 26651 44356 27016 44384
rect 28382 44356 28540 44384
rect 26651 44353 26663 44356
rect 26605 44347 26663 44353
rect 28534 44344 28540 44356
rect 28592 44344 28598 44396
rect 44821 44387 44879 44393
rect 44821 44353 44833 44387
rect 44867 44384 44879 44387
rect 45278 44384 45284 44396
rect 44867 44356 45284 44384
rect 44867 44353 44879 44356
rect 44821 44347 44879 44353
rect 45278 44344 45284 44356
rect 45336 44344 45342 44396
rect 26970 44276 26976 44328
rect 27028 44276 27034 44328
rect 44358 44316 44364 44328
rect 27080 44288 44364 44316
rect 27080 44248 27108 44288
rect 44358 44276 44364 44288
rect 44416 44316 44422 44328
rect 44545 44319 44603 44325
rect 44545 44316 44557 44319
rect 44416 44288 44557 44316
rect 44416 44276 44422 44288
rect 44545 44285 44557 44288
rect 44591 44285 44603 44319
rect 44545 44279 44603 44285
rect 25976 44220 27108 44248
rect 23382 44180 23388 44192
rect 20456 44152 23388 44180
rect 19797 44143 19855 44149
rect 23382 44140 23388 44152
rect 23440 44140 23446 44192
rect 25314 44140 25320 44192
rect 25372 44140 25378 44192
rect 26510 44140 26516 44192
rect 26568 44180 26574 44192
rect 27890 44180 27896 44192
rect 26568 44152 27896 44180
rect 26568 44140 26574 44152
rect 27890 44140 27896 44152
rect 27948 44180 27954 44192
rect 28721 44183 28779 44189
rect 28721 44180 28733 44183
rect 27948 44152 28733 44180
rect 27948 44140 27954 44152
rect 28721 44149 28733 44152
rect 28767 44149 28779 44183
rect 28721 44143 28779 44149
rect 1104 44090 45172 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 45172 44090
rect 1104 44016 45172 44038
rect 7377 43979 7435 43985
rect 7377 43945 7389 43979
rect 7423 43976 7435 43979
rect 8202 43976 8208 43988
rect 7423 43948 8208 43976
rect 7423 43945 7435 43948
rect 7377 43939 7435 43945
rect 8202 43936 8208 43948
rect 8260 43936 8266 43988
rect 10505 43979 10563 43985
rect 10505 43945 10517 43979
rect 10551 43976 10563 43979
rect 10686 43976 10692 43988
rect 10551 43948 10692 43976
rect 10551 43945 10563 43948
rect 10505 43939 10563 43945
rect 10686 43936 10692 43948
rect 10744 43936 10750 43988
rect 13814 43936 13820 43988
rect 13872 43976 13878 43988
rect 14093 43979 14151 43985
rect 14093 43976 14105 43979
rect 13872 43948 14105 43976
rect 13872 43936 13878 43948
rect 14093 43945 14105 43948
rect 14139 43945 14151 43979
rect 14093 43939 14151 43945
rect 15378 43936 15384 43988
rect 15436 43976 15442 43988
rect 15749 43979 15807 43985
rect 15749 43976 15761 43979
rect 15436 43948 15761 43976
rect 15436 43936 15442 43948
rect 15749 43945 15761 43948
rect 15795 43945 15807 43979
rect 15749 43939 15807 43945
rect 18325 43979 18383 43985
rect 18325 43945 18337 43979
rect 18371 43976 18383 43979
rect 18414 43976 18420 43988
rect 18371 43948 18420 43976
rect 18371 43945 18383 43948
rect 18325 43939 18383 43945
rect 18414 43936 18420 43948
rect 18472 43936 18478 43988
rect 18874 43936 18880 43988
rect 18932 43976 18938 43988
rect 19245 43979 19303 43985
rect 19245 43976 19257 43979
rect 18932 43948 19257 43976
rect 18932 43936 18938 43948
rect 19245 43945 19257 43948
rect 19291 43945 19303 43979
rect 19245 43939 19303 43945
rect 22186 43936 22192 43988
rect 22244 43936 22250 43988
rect 23658 43936 23664 43988
rect 23716 43936 23722 43988
rect 10597 43911 10655 43917
rect 10597 43908 10609 43911
rect 9968 43880 10609 43908
rect 9968 43849 9996 43880
rect 10597 43877 10609 43880
rect 10643 43877 10655 43911
rect 10597 43871 10655 43877
rect 9953 43843 10011 43849
rect 9953 43809 9965 43843
rect 9999 43809 10011 43843
rect 9953 43803 10011 43809
rect 13170 43800 13176 43852
rect 13228 43840 13234 43852
rect 14645 43843 14703 43849
rect 14645 43840 14657 43843
rect 13228 43812 14657 43840
rect 13228 43800 13234 43812
rect 14645 43809 14657 43812
rect 14691 43840 14703 43843
rect 14691 43812 15240 43840
rect 14691 43809 14703 43812
rect 14645 43803 14703 43809
rect 11974 43732 11980 43784
rect 12032 43732 12038 43784
rect 12434 43732 12440 43784
rect 12492 43732 12498 43784
rect 14461 43775 14519 43781
rect 14461 43741 14473 43775
rect 14507 43772 14519 43775
rect 14734 43772 14740 43784
rect 14507 43744 14740 43772
rect 14507 43741 14519 43744
rect 14461 43735 14519 43741
rect 14734 43732 14740 43744
rect 14792 43732 14798 43784
rect 7101 43707 7159 43713
rect 7101 43673 7113 43707
rect 7147 43704 7159 43707
rect 11732 43707 11790 43713
rect 7147 43676 8064 43704
rect 7147 43673 7159 43676
rect 7101 43667 7159 43673
rect 8036 43648 8064 43676
rect 11732 43673 11744 43707
rect 11778 43704 11790 43707
rect 12452 43704 12480 43732
rect 11778 43676 12480 43704
rect 11778 43673 11790 43676
rect 11732 43667 11790 43673
rect 12526 43664 12532 43716
rect 12584 43704 12590 43716
rect 12894 43704 12900 43716
rect 12584 43676 12900 43704
rect 12584 43664 12590 43676
rect 12894 43664 12900 43676
rect 12952 43704 12958 43716
rect 15105 43707 15163 43713
rect 15105 43704 15117 43707
rect 12952 43676 15117 43704
rect 12952 43664 12958 43676
rect 15105 43673 15117 43676
rect 15151 43673 15163 43707
rect 15212 43704 15240 43812
rect 15286 43800 15292 43852
rect 15344 43840 15350 43852
rect 16482 43840 16488 43852
rect 15344 43812 16488 43840
rect 15344 43800 15350 43812
rect 15396 43781 15424 43812
rect 16482 43800 16488 43812
rect 16540 43840 16546 43852
rect 18874 43840 18880 43852
rect 16540 43812 18880 43840
rect 16540 43800 16546 43812
rect 18874 43800 18880 43812
rect 18932 43800 18938 43852
rect 19797 43843 19855 43849
rect 19797 43809 19809 43843
rect 19843 43809 19855 43843
rect 22741 43843 22799 43849
rect 22741 43840 22753 43843
rect 19797 43803 19855 43809
rect 22204 43812 22753 43840
rect 15381 43775 15439 43781
rect 15381 43741 15393 43775
rect 15427 43741 15439 43775
rect 15381 43735 15439 43741
rect 15933 43775 15991 43781
rect 15933 43741 15945 43775
rect 15979 43772 15991 43775
rect 16666 43772 16672 43784
rect 15979 43744 16672 43772
rect 15979 43741 15991 43744
rect 15933 43735 15991 43741
rect 16666 43732 16672 43744
rect 16724 43732 16730 43784
rect 18785 43775 18843 43781
rect 18785 43741 18797 43775
rect 18831 43772 18843 43775
rect 19610 43772 19616 43784
rect 18831 43744 19616 43772
rect 18831 43741 18843 43744
rect 18785 43735 18843 43741
rect 19610 43732 19616 43744
rect 19668 43732 19674 43784
rect 17310 43704 17316 43716
rect 15212 43676 17316 43704
rect 15105 43667 15163 43673
rect 17310 43664 17316 43676
rect 17368 43704 17374 43716
rect 19812 43704 19840 43803
rect 22204 43781 22232 43812
rect 22741 43809 22753 43812
rect 22787 43809 22799 43843
rect 22741 43803 22799 43809
rect 23385 43843 23443 43849
rect 23385 43809 23397 43843
rect 23431 43840 23443 43843
rect 23566 43840 23572 43852
rect 23431 43812 23572 43840
rect 23431 43809 23443 43812
rect 23385 43803 23443 43809
rect 23566 43800 23572 43812
rect 23624 43800 23630 43852
rect 25961 43843 26019 43849
rect 25961 43809 25973 43843
rect 26007 43840 26019 43843
rect 26234 43840 26240 43852
rect 26007 43812 26240 43840
rect 26007 43809 26019 43812
rect 25961 43803 26019 43809
rect 26234 43800 26240 43812
rect 26292 43840 26298 43852
rect 26970 43840 26976 43852
rect 26292 43812 26976 43840
rect 26292 43800 26298 43812
rect 26970 43800 26976 43812
rect 27028 43800 27034 43852
rect 29914 43800 29920 43852
rect 29972 43840 29978 43852
rect 30285 43843 30343 43849
rect 30285 43840 30297 43843
rect 29972 43812 30297 43840
rect 29972 43800 29978 43812
rect 30285 43809 30297 43812
rect 30331 43809 30343 43843
rect 30285 43803 30343 43809
rect 31846 43800 31852 43852
rect 31904 43840 31910 43852
rect 32125 43843 32183 43849
rect 32125 43840 32137 43843
rect 31904 43812 32137 43840
rect 31904 43800 31910 43812
rect 32125 43809 32137 43812
rect 32171 43809 32183 43843
rect 32125 43803 32183 43809
rect 33042 43800 33048 43852
rect 33100 43840 33106 43852
rect 33597 43843 33655 43849
rect 33597 43840 33609 43843
rect 33100 43812 33609 43840
rect 33100 43800 33106 43812
rect 33597 43809 33609 43812
rect 33643 43809 33655 43843
rect 33597 43803 33655 43809
rect 22189 43775 22247 43781
rect 22189 43741 22201 43775
rect 22235 43741 22247 43775
rect 22189 43735 22247 43741
rect 22373 43775 22431 43781
rect 22373 43741 22385 43775
rect 22419 43741 22431 43775
rect 22373 43735 22431 43741
rect 20438 43704 20444 43716
rect 17368 43676 20444 43704
rect 17368 43664 17374 43676
rect 20438 43664 20444 43676
rect 20496 43664 20502 43716
rect 8018 43596 8024 43648
rect 8076 43636 8082 43648
rect 14458 43636 14464 43648
rect 8076 43608 14464 43636
rect 8076 43596 8082 43608
rect 14458 43596 14464 43608
rect 14516 43596 14522 43648
rect 14550 43596 14556 43648
rect 14608 43596 14614 43648
rect 18414 43596 18420 43648
rect 18472 43636 18478 43648
rect 18693 43639 18751 43645
rect 18693 43636 18705 43639
rect 18472 43608 18705 43636
rect 18472 43596 18478 43608
rect 18693 43605 18705 43608
rect 18739 43636 18751 43639
rect 19058 43636 19064 43648
rect 18739 43608 19064 43636
rect 18739 43605 18751 43608
rect 18693 43599 18751 43605
rect 19058 43596 19064 43608
rect 19116 43596 19122 43648
rect 19705 43639 19763 43645
rect 19705 43605 19717 43639
rect 19751 43636 19763 43639
rect 20070 43636 20076 43648
rect 19751 43608 20076 43636
rect 19751 43605 19763 43608
rect 19705 43599 19763 43605
rect 20070 43596 20076 43608
rect 20128 43596 20134 43648
rect 22388 43636 22416 43735
rect 23474 43732 23480 43784
rect 23532 43772 23538 43784
rect 25225 43775 25283 43781
rect 23532 43744 23888 43772
rect 23532 43732 23538 43744
rect 23645 43707 23703 43713
rect 23645 43673 23657 43707
rect 23691 43704 23703 43707
rect 23750 43704 23756 43716
rect 23691 43676 23756 43704
rect 23691 43673 23703 43676
rect 23645 43667 23703 43673
rect 23750 43664 23756 43676
rect 23808 43664 23814 43716
rect 23860 43713 23888 43744
rect 25225 43741 25237 43775
rect 25271 43772 25283 43775
rect 25314 43772 25320 43784
rect 25271 43744 25320 43772
rect 25271 43741 25283 43744
rect 25225 43735 25283 43741
rect 25314 43732 25320 43744
rect 25372 43732 25378 43784
rect 33873 43775 33931 43781
rect 33873 43741 33885 43775
rect 33919 43772 33931 43775
rect 33919 43744 34008 43772
rect 33919 43741 33931 43744
rect 33873 43735 33931 43741
rect 23845 43707 23903 43713
rect 23845 43673 23857 43707
rect 23891 43673 23903 43707
rect 23845 43667 23903 43673
rect 26237 43707 26295 43713
rect 26237 43673 26249 43707
rect 26283 43673 26295 43707
rect 30561 43707 30619 43713
rect 27462 43676 28580 43704
rect 26237 43667 26295 43673
rect 22646 43636 22652 43648
rect 22388 43608 22652 43636
rect 22646 43596 22652 43608
rect 22704 43636 22710 43648
rect 23477 43639 23535 43645
rect 23477 43636 23489 43639
rect 22704 43608 23489 43636
rect 22704 43596 22710 43608
rect 23477 43605 23489 43608
rect 23523 43605 23535 43639
rect 23477 43599 23535 43605
rect 25409 43639 25467 43645
rect 25409 43605 25421 43639
rect 25455 43636 25467 43639
rect 26252 43636 26280 43667
rect 28552 43648 28580 43676
rect 30561 43673 30573 43707
rect 30607 43704 30619 43707
rect 30834 43704 30840 43716
rect 30607 43676 30840 43704
rect 30607 43673 30619 43676
rect 30561 43667 30619 43673
rect 30834 43664 30840 43676
rect 30892 43664 30898 43716
rect 31786 43676 32430 43704
rect 25455 43608 26280 43636
rect 25455 43605 25467 43608
rect 25409 43599 25467 43605
rect 27706 43596 27712 43648
rect 27764 43596 27770 43648
rect 28534 43596 28540 43648
rect 28592 43636 28598 43648
rect 31864 43636 31892 43676
rect 33980 43648 34008 43744
rect 28592 43608 31892 43636
rect 28592 43596 28598 43608
rect 31938 43596 31944 43648
rect 31996 43636 32002 43648
rect 32033 43639 32091 43645
rect 32033 43636 32045 43639
rect 31996 43608 32045 43636
rect 31996 43596 32002 43608
rect 32033 43605 32045 43608
rect 32079 43605 32091 43639
rect 32033 43599 32091 43605
rect 33962 43596 33968 43648
rect 34020 43596 34026 43648
rect 1104 43546 45172 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 45172 43546
rect 1104 43472 45172 43494
rect 7742 43392 7748 43444
rect 7800 43432 7806 43444
rect 8018 43432 8024 43444
rect 7800 43404 8024 43432
rect 7800 43392 7806 43404
rect 8018 43392 8024 43404
rect 8076 43392 8082 43444
rect 29914 43392 29920 43444
rect 29972 43392 29978 43444
rect 7466 43324 7472 43376
rect 7524 43364 7530 43376
rect 7653 43367 7711 43373
rect 7653 43364 7665 43367
rect 7524 43336 7665 43364
rect 7524 43324 7530 43336
rect 7653 43333 7665 43336
rect 7699 43364 7711 43367
rect 7926 43364 7932 43376
rect 7699 43336 7932 43364
rect 7699 43333 7711 43336
rect 7653 43327 7711 43333
rect 7926 43324 7932 43336
rect 7984 43324 7990 43376
rect 8389 43367 8447 43373
rect 8389 43333 8401 43367
rect 8435 43364 8447 43367
rect 8846 43364 8852 43376
rect 8435 43336 8852 43364
rect 8435 43333 8447 43336
rect 8389 43327 8447 43333
rect 8846 43324 8852 43336
rect 8904 43364 8910 43376
rect 9306 43364 9312 43376
rect 8904 43336 9312 43364
rect 8904 43324 8910 43336
rect 9306 43324 9312 43336
rect 9364 43324 9370 43376
rect 27433 43367 27491 43373
rect 27433 43364 27445 43367
rect 26804 43336 27445 43364
rect 26804 43308 26832 43336
rect 27433 43333 27445 43336
rect 27479 43333 27491 43367
rect 29932 43364 29960 43392
rect 32214 43364 32220 43376
rect 29932 43336 32220 43364
rect 27433 43327 27491 43333
rect 32214 43324 32220 43336
rect 32272 43324 32278 43376
rect 8294 43305 8300 43308
rect 8292 43296 8300 43305
rect 8255 43268 8300 43296
rect 8292 43259 8300 43268
rect 8294 43256 8300 43259
rect 8352 43256 8358 43308
rect 8478 43256 8484 43308
rect 8536 43256 8542 43308
rect 8664 43299 8722 43305
rect 8664 43265 8676 43299
rect 8710 43265 8722 43299
rect 8664 43259 8722 43265
rect 6914 43188 6920 43240
rect 6972 43188 6978 43240
rect 8680 43228 8708 43259
rect 8754 43256 8760 43308
rect 8812 43256 8818 43308
rect 13354 43256 13360 43308
rect 13412 43256 13418 43308
rect 20717 43299 20775 43305
rect 20717 43265 20729 43299
rect 20763 43296 20775 43299
rect 20806 43296 20812 43308
rect 20763 43268 20812 43296
rect 20763 43265 20775 43268
rect 20717 43259 20775 43265
rect 20806 43256 20812 43268
rect 20864 43256 20870 43308
rect 26786 43256 26792 43308
rect 26844 43256 26850 43308
rect 26878 43256 26884 43308
rect 26936 43296 26942 43308
rect 27249 43299 27307 43305
rect 27249 43296 27261 43299
rect 26936 43268 27261 43296
rect 26936 43256 26942 43268
rect 27249 43265 27261 43268
rect 27295 43265 27307 43299
rect 27249 43259 27307 43265
rect 9493 43231 9551 43237
rect 9493 43228 9505 43231
rect 8680 43200 9505 43228
rect 9493 43197 9505 43200
rect 9539 43197 9551 43231
rect 9493 43191 9551 43197
rect 10137 43231 10195 43237
rect 10137 43197 10149 43231
rect 10183 43228 10195 43231
rect 10686 43228 10692 43240
rect 10183 43200 10692 43228
rect 10183 43197 10195 43200
rect 10137 43191 10195 43197
rect 10686 43188 10692 43200
rect 10744 43188 10750 43240
rect 16666 43188 16672 43240
rect 16724 43188 16730 43240
rect 32232 43228 32260 43324
rect 33870 43256 33876 43308
rect 33928 43256 33934 43308
rect 33962 43228 33968 43240
rect 32232 43200 33968 43228
rect 33962 43188 33968 43200
rect 34020 43188 34026 43240
rect 34238 43188 34244 43240
rect 34296 43188 34302 43240
rect 35360 43228 35388 43282
rect 35526 43256 35532 43308
rect 35584 43296 35590 43308
rect 35805 43299 35863 43305
rect 35805 43296 35817 43299
rect 35584 43268 35817 43296
rect 35584 43256 35590 43268
rect 35805 43265 35817 43268
rect 35851 43265 35863 43299
rect 35805 43259 35863 43265
rect 35360 43200 36032 43228
rect 31726 43132 32720 43160
rect 31726 43104 31754 43132
rect 7466 43052 7472 43104
rect 7524 43052 7530 43104
rect 8110 43052 8116 43104
rect 8168 43052 8174 43104
rect 13170 43052 13176 43104
rect 13228 43052 13234 43104
rect 17310 43052 17316 43104
rect 17368 43052 17374 43104
rect 19150 43052 19156 43104
rect 19208 43092 19214 43104
rect 19429 43095 19487 43101
rect 19429 43092 19441 43095
rect 19208 43064 19441 43092
rect 19208 43052 19214 43064
rect 19429 43061 19441 43064
rect 19475 43092 19487 43095
rect 21174 43092 21180 43104
rect 19475 43064 21180 43092
rect 19475 43061 19487 43064
rect 19429 43055 19487 43061
rect 21174 43052 21180 43064
rect 21232 43052 21238 43104
rect 26970 43052 26976 43104
rect 27028 43092 27034 43104
rect 27065 43095 27123 43101
rect 27065 43092 27077 43095
rect 27028 43064 27077 43092
rect 27028 43052 27034 43064
rect 27065 43061 27077 43064
rect 27111 43061 27123 43095
rect 27065 43055 27123 43061
rect 31662 43052 31668 43104
rect 31720 43064 31754 43104
rect 31720 43052 31726 43064
rect 32214 43052 32220 43104
rect 32272 43092 32278 43104
rect 32401 43095 32459 43101
rect 32401 43092 32413 43095
rect 32272 43064 32413 43092
rect 32272 43052 32278 43064
rect 32401 43061 32413 43064
rect 32447 43061 32459 43095
rect 32692 43092 32720 43132
rect 35526 43092 35532 43104
rect 32692 43064 35532 43092
rect 32401 43055 32459 43061
rect 35526 43052 35532 43064
rect 35584 43052 35590 43104
rect 35710 43052 35716 43104
rect 35768 43052 35774 43104
rect 36004 43101 36032 43200
rect 35989 43095 36047 43101
rect 35989 43061 36001 43095
rect 36035 43092 36047 43095
rect 36906 43092 36912 43104
rect 36035 43064 36912 43092
rect 36035 43061 36047 43064
rect 35989 43055 36047 43061
rect 36906 43052 36912 43064
rect 36964 43052 36970 43104
rect 1104 43002 45172 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 45172 43002
rect 1104 42928 45172 42950
rect 7119 42891 7177 42897
rect 7119 42857 7131 42891
rect 7165 42888 7177 42891
rect 7466 42888 7472 42900
rect 7165 42860 7472 42888
rect 7165 42857 7177 42860
rect 7119 42851 7177 42857
rect 7466 42848 7472 42860
rect 7524 42848 7530 42900
rect 14550 42848 14556 42900
rect 14608 42888 14614 42900
rect 14829 42891 14887 42897
rect 14829 42888 14841 42891
rect 14608 42860 14841 42888
rect 14608 42848 14614 42860
rect 14829 42857 14841 42860
rect 14875 42857 14887 42891
rect 14829 42851 14887 42857
rect 16209 42891 16267 42897
rect 16209 42857 16221 42891
rect 16255 42888 16267 42891
rect 16666 42888 16672 42900
rect 16255 42860 16672 42888
rect 16255 42857 16267 42860
rect 16209 42851 16267 42857
rect 16666 42848 16672 42860
rect 16724 42848 16730 42900
rect 17310 42848 17316 42900
rect 17368 42888 17374 42900
rect 17785 42891 17843 42897
rect 17785 42888 17797 42891
rect 17368 42860 17797 42888
rect 17368 42848 17374 42860
rect 17785 42857 17797 42860
rect 17831 42857 17843 42891
rect 17785 42851 17843 42857
rect 25222 42848 25228 42900
rect 25280 42888 25286 42900
rect 28534 42888 28540 42900
rect 25280 42860 28540 42888
rect 25280 42848 25286 42860
rect 28534 42848 28540 42860
rect 28592 42848 28598 42900
rect 31938 42888 31944 42900
rect 30760 42860 31944 42888
rect 17972 42792 18184 42820
rect 7561 42755 7619 42761
rect 7561 42752 7573 42755
rect 6012 42724 7573 42752
rect 3878 42644 3884 42696
rect 3936 42644 3942 42696
rect 4065 42687 4123 42693
rect 4065 42653 4077 42687
rect 4111 42684 4123 42687
rect 4111 42656 4200 42684
rect 4111 42653 4123 42656
rect 4065 42647 4123 42653
rect 4172 42560 4200 42656
rect 4890 42644 4896 42696
rect 4948 42644 4954 42696
rect 5350 42644 5356 42696
rect 5408 42684 5414 42696
rect 6012 42684 6040 42724
rect 7561 42721 7573 42724
rect 7607 42752 7619 42755
rect 8018 42752 8024 42764
rect 7607 42724 8024 42752
rect 7607 42721 7619 42724
rect 7561 42715 7619 42721
rect 8018 42712 8024 42724
rect 8076 42712 8082 42764
rect 8110 42712 8116 42764
rect 8168 42712 8174 42764
rect 8294 42712 8300 42764
rect 8352 42752 8358 42764
rect 11790 42752 11796 42764
rect 8352 42724 11796 42752
rect 8352 42712 8358 42724
rect 11790 42712 11796 42724
rect 11848 42712 11854 42764
rect 12621 42755 12679 42761
rect 12621 42721 12633 42755
rect 12667 42752 12679 42755
rect 13817 42755 13875 42761
rect 12667 42724 13768 42752
rect 12667 42721 12679 42724
rect 12621 42715 12679 42721
rect 13740 42696 13768 42724
rect 13817 42721 13829 42755
rect 13863 42752 13875 42755
rect 14734 42752 14740 42764
rect 13863 42724 14740 42752
rect 13863 42721 13875 42724
rect 13817 42715 13875 42721
rect 14734 42712 14740 42724
rect 14792 42712 14798 42764
rect 16301 42755 16359 42761
rect 16301 42752 16313 42755
rect 15948 42724 16313 42752
rect 5408 42670 6040 42684
rect 7377 42687 7435 42693
rect 5408 42656 6026 42670
rect 5408 42644 5414 42656
rect 7377 42653 7389 42687
rect 7423 42684 7435 42687
rect 7423 42656 7512 42684
rect 7423 42653 7435 42656
rect 7377 42647 7435 42653
rect 7484 42560 7512 42656
rect 7834 42644 7840 42696
rect 7892 42684 7898 42696
rect 8202 42684 8208 42696
rect 7892 42656 8208 42684
rect 7892 42644 7898 42656
rect 8202 42644 8208 42656
rect 8260 42644 8266 42696
rect 10594 42644 10600 42696
rect 10652 42684 10658 42696
rect 10652 42656 11270 42684
rect 10652 42644 10658 42656
rect 12802 42644 12808 42696
rect 12860 42684 12866 42696
rect 13265 42687 13323 42693
rect 13265 42684 13277 42687
rect 12860 42656 13277 42684
rect 12860 42644 12866 42656
rect 13265 42653 13277 42656
rect 13311 42653 13323 42687
rect 13265 42647 13323 42653
rect 13449 42687 13507 42693
rect 13449 42653 13461 42687
rect 13495 42653 13507 42687
rect 13633 42687 13691 42693
rect 13633 42684 13645 42687
rect 13449 42647 13507 42653
rect 13556 42656 13645 42684
rect 9030 42576 9036 42628
rect 9088 42576 9094 42628
rect 10781 42619 10839 42625
rect 10781 42585 10793 42619
rect 10827 42616 10839 42619
rect 11054 42616 11060 42628
rect 10827 42588 11060 42616
rect 10827 42585 10839 42588
rect 10781 42579 10839 42585
rect 11054 42576 11060 42588
rect 11112 42576 11118 42628
rect 12345 42619 12403 42625
rect 12345 42585 12357 42619
rect 12391 42616 12403 42619
rect 12713 42619 12771 42625
rect 12713 42616 12725 42619
rect 12391 42588 12725 42616
rect 12391 42585 12403 42588
rect 12345 42579 12403 42585
rect 12713 42585 12725 42588
rect 12759 42585 12771 42619
rect 12713 42579 12771 42585
rect 4154 42508 4160 42560
rect 4212 42508 4218 42560
rect 4249 42551 4307 42557
rect 4249 42517 4261 42551
rect 4295 42548 4307 42551
rect 4614 42548 4620 42560
rect 4295 42520 4620 42548
rect 4295 42517 4307 42520
rect 4249 42511 4307 42517
rect 4614 42508 4620 42520
rect 4672 42508 4678 42560
rect 5442 42508 5448 42560
rect 5500 42508 5506 42560
rect 5629 42551 5687 42557
rect 5629 42517 5641 42551
rect 5675 42548 5687 42551
rect 6454 42548 6460 42560
rect 5675 42520 6460 42548
rect 5675 42517 5687 42520
rect 5629 42511 5687 42517
rect 6454 42508 6460 42520
rect 6512 42508 6518 42560
rect 7466 42508 7472 42560
rect 7524 42508 7530 42560
rect 8757 42551 8815 42557
rect 8757 42517 8769 42551
rect 8803 42548 8815 42551
rect 9122 42548 9128 42560
rect 8803 42520 9128 42548
rect 8803 42517 8815 42520
rect 8757 42511 8815 42517
rect 9122 42508 9128 42520
rect 9180 42508 9186 42560
rect 10873 42551 10931 42557
rect 10873 42517 10885 42551
rect 10919 42548 10931 42551
rect 11698 42548 11704 42560
rect 10919 42520 11704 42548
rect 10919 42517 10931 42520
rect 10873 42511 10931 42517
rect 11698 42508 11704 42520
rect 11756 42548 11762 42560
rect 13464 42548 13492 42647
rect 13556 42560 13584 42656
rect 13633 42653 13645 42656
rect 13679 42653 13691 42687
rect 13633 42647 13691 42653
rect 13722 42644 13728 42696
rect 13780 42644 13786 42696
rect 14642 42644 14648 42696
rect 14700 42644 14706 42696
rect 15381 42687 15439 42693
rect 15381 42653 15393 42687
rect 15427 42653 15439 42687
rect 15381 42647 15439 42653
rect 13906 42576 13912 42628
rect 13964 42616 13970 42628
rect 15396 42616 15424 42647
rect 15562 42644 15568 42696
rect 15620 42644 15626 42696
rect 15713 42687 15771 42693
rect 15713 42653 15725 42687
rect 15759 42684 15771 42687
rect 15948 42684 15976 42724
rect 16301 42721 16313 42724
rect 16347 42752 16359 42755
rect 17972 42752 18000 42792
rect 16347 42724 18000 42752
rect 16347 42721 16359 42724
rect 16301 42715 16359 42721
rect 15759 42656 15976 42684
rect 16071 42687 16129 42693
rect 15759 42653 15771 42656
rect 15713 42647 15771 42653
rect 16071 42653 16083 42687
rect 16117 42684 16129 42687
rect 16117 42656 16528 42684
rect 16117 42653 16129 42656
rect 16071 42647 16129 42653
rect 16500 42628 16528 42656
rect 18046 42644 18052 42696
rect 18104 42644 18110 42696
rect 18156 42693 18184 42792
rect 18248 42724 22600 42752
rect 18141 42687 18199 42693
rect 18141 42653 18153 42687
rect 18187 42653 18199 42687
rect 18141 42647 18199 42653
rect 15838 42616 15844 42628
rect 13964 42588 15424 42616
rect 15488 42588 15844 42616
rect 13964 42576 13970 42588
rect 11756 42520 13492 42548
rect 11756 42508 11762 42520
rect 13538 42508 13544 42560
rect 13596 42508 13602 42560
rect 14090 42508 14096 42560
rect 14148 42508 14154 42560
rect 14182 42508 14188 42560
rect 14240 42548 14246 42560
rect 15488 42548 15516 42588
rect 15838 42576 15844 42588
rect 15896 42576 15902 42628
rect 15933 42619 15991 42625
rect 15933 42585 15945 42619
rect 15979 42585 15991 42619
rect 15933 42579 15991 42585
rect 14240 42520 15516 42548
rect 14240 42508 14246 42520
rect 15746 42508 15752 42560
rect 15804 42548 15810 42560
rect 15948 42548 15976 42579
rect 16482 42576 16488 42628
rect 16540 42576 16546 42628
rect 17494 42616 17500 42628
rect 17342 42588 17500 42616
rect 17494 42576 17500 42588
rect 17552 42616 17558 42628
rect 18248 42616 18276 42724
rect 22572 42696 22600 42724
rect 22830 42712 22836 42764
rect 22888 42752 22894 42764
rect 23017 42755 23075 42761
rect 23017 42752 23029 42755
rect 22888 42724 23029 42752
rect 22888 42712 22894 42724
rect 23017 42721 23029 42724
rect 23063 42752 23075 42755
rect 23201 42755 23259 42761
rect 23201 42752 23213 42755
rect 23063 42724 23213 42752
rect 23063 42721 23075 42724
rect 23017 42715 23075 42721
rect 23201 42721 23213 42724
rect 23247 42721 23259 42755
rect 23201 42715 23259 42721
rect 24394 42712 24400 42764
rect 24452 42752 24458 42764
rect 26234 42752 26240 42764
rect 24452 42724 26240 42752
rect 24452 42712 24458 42724
rect 26234 42712 26240 42724
rect 26292 42752 26298 42764
rect 26694 42752 26700 42764
rect 26292 42724 26700 42752
rect 26292 42712 26298 42724
rect 26694 42712 26700 42724
rect 26752 42712 26758 42764
rect 30193 42755 30251 42761
rect 30193 42721 30205 42755
rect 30239 42721 30251 42755
rect 30760 42752 30788 42860
rect 31938 42848 31944 42860
rect 31996 42888 32002 42900
rect 32769 42891 32827 42897
rect 31996 42860 32076 42888
rect 31996 42848 32002 42860
rect 31938 42752 31944 42764
rect 30193 42715 30251 42721
rect 30300 42724 30788 42752
rect 30852 42724 31944 42752
rect 18325 42687 18383 42693
rect 18325 42653 18337 42687
rect 18371 42653 18383 42687
rect 18325 42647 18383 42653
rect 17552 42588 18276 42616
rect 18340 42616 18368 42647
rect 18782 42644 18788 42696
rect 18840 42644 18846 42696
rect 19334 42644 19340 42696
rect 19392 42644 19398 42696
rect 21174 42644 21180 42696
rect 21232 42684 21238 42696
rect 21269 42687 21327 42693
rect 21269 42684 21281 42687
rect 21232 42656 21281 42684
rect 21232 42644 21238 42656
rect 21269 42653 21281 42656
rect 21315 42653 21327 42687
rect 21269 42647 21327 42653
rect 22554 42644 22560 42696
rect 22612 42684 22618 42696
rect 22612 42656 22678 42684
rect 22612 42644 22618 42656
rect 24026 42644 24032 42696
rect 24084 42644 24090 42696
rect 25976 42656 29960 42684
rect 18340 42588 21496 42616
rect 17552 42576 17558 42588
rect 17126 42548 17132 42560
rect 15804 42520 17132 42548
rect 15804 42508 15810 42520
rect 17126 42508 17132 42520
rect 17184 42508 17190 42560
rect 17586 42508 17592 42560
rect 17644 42548 17650 42560
rect 18340 42548 18368 42588
rect 17644 42520 18368 42548
rect 17644 42508 17650 42520
rect 18506 42508 18512 42560
rect 18564 42508 18570 42560
rect 18601 42551 18659 42557
rect 18601 42517 18613 42551
rect 18647 42548 18659 42551
rect 18690 42548 18696 42560
rect 18647 42520 18696 42548
rect 18647 42517 18659 42520
rect 18601 42511 18659 42517
rect 18690 42508 18696 42520
rect 18748 42508 18754 42560
rect 19978 42508 19984 42560
rect 20036 42508 20042 42560
rect 21468 42548 21496 42588
rect 21542 42576 21548 42628
rect 21600 42576 21606 42628
rect 24673 42619 24731 42625
rect 24673 42585 24685 42619
rect 24719 42585 24731 42619
rect 24673 42579 24731 42585
rect 23474 42548 23480 42560
rect 21468 42520 23480 42548
rect 23474 42508 23480 42520
rect 23532 42508 23538 42560
rect 23842 42508 23848 42560
rect 23900 42508 23906 42560
rect 24213 42551 24271 42557
rect 24213 42517 24225 42551
rect 24259 42548 24271 42551
rect 24688 42548 24716 42579
rect 25222 42576 25228 42628
rect 25280 42576 25286 42628
rect 24259 42520 24716 42548
rect 24259 42517 24271 42520
rect 24213 42511 24271 42517
rect 25498 42508 25504 42560
rect 25556 42548 25562 42560
rect 25976 42548 26004 42656
rect 27982 42576 27988 42628
rect 28040 42576 28046 42628
rect 25556 42520 26004 42548
rect 25556 42508 25562 42520
rect 26142 42508 26148 42560
rect 26200 42508 26206 42560
rect 26694 42508 26700 42560
rect 26752 42508 26758 42560
rect 29932 42548 29960 42656
rect 30006 42576 30012 42628
rect 30064 42616 30070 42628
rect 30208 42616 30236 42715
rect 30300 42693 30328 42724
rect 30285 42687 30343 42693
rect 30285 42653 30297 42687
rect 30331 42653 30343 42687
rect 30745 42687 30803 42693
rect 30745 42684 30757 42687
rect 30285 42647 30343 42653
rect 30576 42656 30757 42684
rect 30576 42616 30604 42656
rect 30745 42653 30757 42656
rect 30791 42684 30803 42687
rect 30852 42684 30880 42724
rect 31938 42712 31944 42724
rect 31996 42712 32002 42764
rect 30791 42656 30880 42684
rect 30929 42687 30987 42693
rect 30791 42653 30803 42656
rect 30745 42647 30803 42653
rect 30929 42653 30941 42687
rect 30975 42684 30987 42687
rect 31018 42684 31024 42696
rect 30975 42656 31024 42684
rect 30975 42653 30987 42656
rect 30929 42647 30987 42653
rect 31018 42644 31024 42656
rect 31076 42684 31082 42696
rect 31846 42684 31852 42696
rect 31076 42656 31852 42684
rect 31076 42644 31082 42656
rect 31846 42644 31852 42656
rect 31904 42644 31910 42696
rect 32048 42693 32076 42860
rect 32769 42857 32781 42891
rect 32815 42888 32827 42891
rect 33042 42888 33048 42900
rect 32815 42860 33048 42888
rect 32815 42857 32827 42860
rect 32769 42851 32827 42857
rect 33042 42848 33048 42860
rect 33100 42848 33106 42900
rect 32490 42780 32496 42832
rect 32548 42820 32554 42832
rect 32548 42792 33640 42820
rect 32548 42780 32554 42792
rect 32784 42724 33180 42752
rect 32033 42687 32091 42693
rect 32033 42653 32045 42687
rect 32079 42684 32091 42687
rect 32674 42684 32680 42696
rect 32079 42656 32680 42684
rect 32079 42653 32091 42656
rect 32033 42647 32091 42653
rect 32674 42644 32680 42656
rect 32732 42644 32738 42696
rect 31389 42619 31447 42625
rect 31389 42616 31401 42619
rect 30064 42588 30604 42616
rect 30760 42588 31401 42616
rect 30064 42576 30070 42588
rect 30760 42560 30788 42588
rect 31389 42585 31401 42588
rect 31435 42585 31447 42619
rect 31389 42579 31447 42585
rect 30374 42548 30380 42560
rect 29932 42520 30380 42548
rect 30374 42508 30380 42520
rect 30432 42508 30438 42560
rect 30650 42508 30656 42560
rect 30708 42508 30714 42560
rect 30742 42508 30748 42560
rect 30800 42508 30806 42560
rect 30929 42551 30987 42557
rect 30929 42517 30941 42551
rect 30975 42548 30987 42551
rect 31754 42548 31760 42560
rect 30975 42520 31760 42548
rect 30975 42517 30987 42520
rect 30929 42511 30987 42517
rect 31754 42508 31760 42520
rect 31812 42508 31818 42560
rect 31864 42548 31892 42644
rect 32582 42576 32588 42628
rect 32640 42616 32646 42628
rect 32784 42616 32812 42724
rect 33152 42693 33180 42724
rect 32953 42687 33011 42693
rect 32953 42684 32965 42687
rect 32640 42588 32812 42616
rect 32876 42656 32965 42684
rect 32640 42576 32646 42588
rect 32490 42548 32496 42560
rect 31864 42520 32496 42548
rect 32490 42508 32496 42520
rect 32548 42508 32554 42560
rect 32876 42548 32904 42656
rect 32953 42653 32965 42656
rect 32999 42653 33011 42687
rect 32953 42647 33011 42653
rect 33137 42687 33195 42693
rect 33137 42653 33149 42687
rect 33183 42653 33195 42687
rect 33137 42647 33195 42653
rect 33226 42644 33232 42696
rect 33284 42693 33290 42696
rect 33284 42687 33313 42693
rect 33301 42653 33313 42687
rect 33284 42647 33313 42653
rect 33413 42687 33471 42693
rect 33413 42653 33425 42687
rect 33459 42684 33471 42687
rect 33505 42687 33563 42693
rect 33505 42684 33517 42687
rect 33459 42656 33517 42684
rect 33459 42653 33471 42656
rect 33413 42647 33471 42653
rect 33505 42653 33517 42656
rect 33551 42653 33563 42687
rect 33612 42684 33640 42792
rect 35250 42712 35256 42764
rect 35308 42752 35314 42764
rect 35710 42752 35716 42764
rect 35308 42724 35716 42752
rect 35308 42712 35314 42724
rect 35710 42712 35716 42724
rect 35768 42712 35774 42764
rect 34057 42687 34115 42693
rect 34057 42684 34069 42687
rect 33612 42656 34069 42684
rect 33505 42647 33563 42653
rect 34057 42653 34069 42656
rect 34103 42653 34115 42687
rect 34057 42647 34115 42653
rect 33284 42644 33290 42647
rect 33045 42619 33103 42625
rect 33045 42585 33057 42619
rect 33091 42616 33103 42619
rect 33091 42588 34928 42616
rect 33091 42585 33103 42588
rect 33045 42579 33103 42585
rect 34900 42560 34928 42588
rect 33134 42548 33140 42560
rect 32876 42520 33140 42548
rect 33134 42508 33140 42520
rect 33192 42508 33198 42560
rect 33318 42508 33324 42560
rect 33376 42548 33382 42560
rect 34701 42551 34759 42557
rect 34701 42548 34713 42551
rect 33376 42520 34713 42548
rect 33376 42508 33382 42520
rect 34701 42517 34713 42520
rect 34747 42517 34759 42551
rect 34701 42511 34759 42517
rect 34882 42508 34888 42560
rect 34940 42508 34946 42560
rect 1104 42458 45172 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 45172 42458
rect 1104 42384 45172 42406
rect 3878 42304 3884 42356
rect 3936 42304 3942 42356
rect 5442 42304 5448 42356
rect 5500 42344 5506 42356
rect 5500 42316 5856 42344
rect 5500 42304 5506 42316
rect 3697 42211 3755 42217
rect 3697 42177 3709 42211
rect 3743 42208 3755 42211
rect 3896 42208 3924 42304
rect 5350 42236 5356 42288
rect 5408 42236 5414 42288
rect 5828 42285 5856 42316
rect 6454 42304 6460 42356
rect 6512 42304 6518 42356
rect 6914 42304 6920 42356
rect 6972 42344 6978 42356
rect 7009 42347 7067 42353
rect 7009 42344 7021 42347
rect 6972 42316 7021 42344
rect 6972 42304 6978 42316
rect 7009 42313 7021 42316
rect 7055 42313 7067 42347
rect 8478 42344 8484 42356
rect 7009 42307 7067 42313
rect 7392 42316 8484 42344
rect 5813 42279 5871 42285
rect 5813 42245 5825 42279
rect 5859 42245 5871 42279
rect 5813 42239 5871 42245
rect 3743 42180 3924 42208
rect 3743 42177 3755 42180
rect 3697 42171 3755 42177
rect 6362 42168 6368 42220
rect 6420 42168 6426 42220
rect 6472 42217 6500 42304
rect 6641 42279 6699 42285
rect 6641 42245 6653 42279
rect 6687 42276 6699 42279
rect 7392 42276 7420 42316
rect 8478 42304 8484 42316
rect 8536 42304 8542 42356
rect 8846 42304 8852 42356
rect 8904 42304 8910 42356
rect 11054 42344 11060 42356
rect 8956 42316 11060 42344
rect 8956 42276 8984 42316
rect 11054 42304 11060 42316
rect 11112 42304 11118 42356
rect 11238 42304 11244 42356
rect 11296 42344 11302 42356
rect 11882 42344 11888 42356
rect 11296 42316 11888 42344
rect 11296 42304 11302 42316
rect 11882 42304 11888 42316
rect 11940 42344 11946 42356
rect 12161 42347 12219 42353
rect 12161 42344 12173 42347
rect 11940 42316 12173 42344
rect 11940 42304 11946 42316
rect 12161 42313 12173 42316
rect 12207 42313 12219 42347
rect 12161 42307 12219 42313
rect 13633 42347 13691 42353
rect 13633 42313 13645 42347
rect 13679 42344 13691 42347
rect 13906 42344 13912 42356
rect 13679 42316 13912 42344
rect 13679 42313 13691 42316
rect 13633 42307 13691 42313
rect 13906 42304 13912 42316
rect 13964 42304 13970 42356
rect 14090 42304 14096 42356
rect 14148 42304 14154 42356
rect 15562 42304 15568 42356
rect 15620 42304 15626 42356
rect 16669 42347 16727 42353
rect 16669 42313 16681 42347
rect 16715 42344 16727 42347
rect 17126 42344 17132 42356
rect 16715 42316 17132 42344
rect 16715 42313 16727 42316
rect 16669 42307 16727 42313
rect 17126 42304 17132 42316
rect 17184 42304 17190 42356
rect 19794 42304 19800 42356
rect 19852 42344 19858 42356
rect 20901 42347 20959 42353
rect 20901 42344 20913 42347
rect 19852 42316 20913 42344
rect 19852 42304 19858 42316
rect 20901 42313 20913 42316
rect 20947 42313 20959 42347
rect 20901 42307 20959 42313
rect 6687 42248 7420 42276
rect 7668 42248 8984 42276
rect 6687 42245 6699 42248
rect 6641 42239 6699 42245
rect 6458 42211 6516 42217
rect 6458 42177 6470 42211
rect 6504 42177 6516 42211
rect 6458 42171 6516 42177
rect 6730 42168 6736 42220
rect 6788 42168 6794 42220
rect 6871 42211 6929 42217
rect 6871 42177 6883 42211
rect 6917 42208 6929 42211
rect 6917 42180 7420 42208
rect 6917 42177 6929 42180
rect 6871 42171 6929 42177
rect 3326 42100 3332 42152
rect 3384 42140 3390 42152
rect 5350 42140 5356 42152
rect 3384 42112 5356 42140
rect 3384 42100 3390 42112
rect 5350 42100 5356 42112
rect 5408 42100 5414 42152
rect 6086 42100 6092 42152
rect 6144 42100 6150 42152
rect 4706 42072 4712 42084
rect 4264 42044 4712 42072
rect 4264 42013 4292 42044
rect 4706 42032 4712 42044
rect 4764 42032 4770 42084
rect 4249 42007 4307 42013
rect 4249 41973 4261 42007
rect 4295 41973 4307 42007
rect 4249 41967 4307 41973
rect 4341 42007 4399 42013
rect 4341 41973 4353 42007
rect 4387 42004 4399 42007
rect 5350 42004 5356 42016
rect 4387 41976 5356 42004
rect 4387 41973 4399 41976
rect 4341 41967 4399 41973
rect 5350 41964 5356 41976
rect 5408 41964 5414 42016
rect 5442 41964 5448 42016
rect 5500 42004 5506 42016
rect 7392 42004 7420 42180
rect 7466 42168 7472 42220
rect 7524 42208 7530 42220
rect 7668 42208 7696 42248
rect 7524 42180 7696 42208
rect 7736 42211 7794 42217
rect 7524 42168 7530 42180
rect 7736 42177 7748 42211
rect 7782 42208 7794 42211
rect 8294 42208 8300 42220
rect 7782 42180 8300 42208
rect 7782 42177 7794 42180
rect 7736 42171 7794 42177
rect 8294 42168 8300 42180
rect 8352 42168 8358 42220
rect 8478 42168 8484 42220
rect 8536 42168 8542 42220
rect 8956 42217 8984 42248
rect 9122 42236 9128 42288
rect 9180 42276 9186 42288
rect 9217 42279 9275 42285
rect 9217 42276 9229 42279
rect 9180 42248 9229 42276
rect 9180 42236 9186 42248
rect 9217 42245 9229 42248
rect 9263 42245 9275 42279
rect 10594 42276 10600 42288
rect 10442 42248 10600 42276
rect 9217 42239 9275 42245
rect 10594 42236 10600 42248
rect 10652 42236 10658 42288
rect 10778 42236 10784 42288
rect 10836 42276 10842 42288
rect 12520 42279 12578 42285
rect 10836 42248 12434 42276
rect 10836 42236 10842 42248
rect 10980 42217 11008 42248
rect 8941 42211 8999 42217
rect 8941 42177 8953 42211
rect 8987 42177 8999 42211
rect 10965 42211 11023 42217
rect 8941 42171 8999 42177
rect 10612 42180 10916 42208
rect 8496 42140 8524 42168
rect 10612 42140 10640 42180
rect 10781 42143 10839 42149
rect 10781 42140 10793 42143
rect 8496 42112 10640 42140
rect 10704 42112 10793 42140
rect 10704 42016 10732 42112
rect 10781 42109 10793 42112
rect 10827 42109 10839 42143
rect 10781 42103 10839 42109
rect 10888 42072 10916 42180
rect 10965 42177 10977 42211
rect 11011 42177 11023 42211
rect 10965 42171 11023 42177
rect 11054 42168 11060 42220
rect 11112 42208 11118 42220
rect 11974 42208 11980 42220
rect 11112 42180 11980 42208
rect 11112 42168 11118 42180
rect 11974 42168 11980 42180
rect 12032 42208 12038 42220
rect 12253 42211 12311 42217
rect 12253 42208 12265 42211
rect 12032 42180 12265 42208
rect 12032 42168 12038 42180
rect 12253 42177 12265 42180
rect 12299 42177 12311 42211
rect 12406 42208 12434 42248
rect 12520 42245 12532 42279
rect 12566 42276 12578 42279
rect 13170 42276 13176 42288
rect 12566 42248 13176 42276
rect 12566 42245 12578 42248
rect 12520 42239 12578 42245
rect 13170 42236 13176 42248
rect 13228 42236 13234 42288
rect 14001 42279 14059 42285
rect 14001 42245 14013 42279
rect 14047 42276 14059 42279
rect 14108 42276 14136 42304
rect 14047 42248 14136 42276
rect 14047 42245 14059 42248
rect 14001 42239 14059 42245
rect 14458 42236 14464 42288
rect 14516 42236 14522 42288
rect 18046 42276 18052 42288
rect 17696 42248 18052 42276
rect 13538 42208 13544 42220
rect 12406 42180 13544 42208
rect 12253 42171 12311 42177
rect 13538 42168 13544 42180
rect 13596 42168 13602 42220
rect 15749 42211 15807 42217
rect 15749 42208 15761 42211
rect 15212 42180 15761 42208
rect 11514 42100 11520 42152
rect 11572 42100 11578 42152
rect 13556 42072 13584 42168
rect 13722 42100 13728 42152
rect 13780 42100 13786 42152
rect 15212 42140 15240 42180
rect 15749 42177 15761 42180
rect 15795 42208 15807 42211
rect 17586 42208 17592 42220
rect 15795 42180 17592 42208
rect 15795 42177 15807 42180
rect 15749 42171 15807 42177
rect 17586 42168 17592 42180
rect 17644 42168 17650 42220
rect 17696 42217 17724 42248
rect 18046 42236 18052 42248
rect 18104 42276 18110 42288
rect 20916 42276 20944 42307
rect 21542 42304 21548 42356
rect 21600 42344 21606 42356
rect 22005 42347 22063 42353
rect 22005 42344 22017 42347
rect 21600 42316 22017 42344
rect 21600 42304 21606 42316
rect 22005 42313 22017 42316
rect 22051 42313 22063 42347
rect 22005 42307 22063 42313
rect 22112 42316 23612 42344
rect 22112 42276 22140 42316
rect 23584 42288 23612 42316
rect 23842 42304 23848 42356
rect 23900 42304 23906 42356
rect 24026 42304 24032 42356
rect 24084 42344 24090 42356
rect 24673 42347 24731 42353
rect 24673 42344 24685 42347
rect 24084 42316 24685 42344
rect 24084 42304 24090 42316
rect 24673 42313 24685 42316
rect 24719 42313 24731 42347
rect 24673 42307 24731 42313
rect 26694 42304 26700 42356
rect 26752 42344 26758 42356
rect 31478 42344 31484 42356
rect 26752 42316 28856 42344
rect 26752 42304 26758 42316
rect 23017 42279 23075 42285
rect 23017 42276 23029 42279
rect 18104 42248 19196 42276
rect 20916 42248 22140 42276
rect 22388 42248 23029 42276
rect 18104 42236 18110 42248
rect 17681 42211 17739 42217
rect 17681 42177 17693 42211
rect 17727 42177 17739 42211
rect 17681 42171 17739 42177
rect 17948 42211 18006 42217
rect 17948 42177 17960 42211
rect 17994 42208 18006 42211
rect 18690 42208 18696 42220
rect 17994 42180 18696 42208
rect 17994 42177 18006 42180
rect 17948 42171 18006 42177
rect 18690 42168 18696 42180
rect 18748 42168 18754 42220
rect 19168 42152 19196 42248
rect 21913 42211 21971 42217
rect 20562 42180 20668 42208
rect 20640 42152 20668 42180
rect 21913 42177 21925 42211
rect 21959 42177 21971 42211
rect 21913 42171 21971 42177
rect 22097 42211 22155 42217
rect 22097 42177 22109 42211
rect 22143 42208 22155 42211
rect 22189 42211 22247 42217
rect 22189 42208 22201 42211
rect 22143 42180 22201 42208
rect 22143 42177 22155 42180
rect 22097 42171 22155 42177
rect 22189 42177 22201 42180
rect 22235 42208 22247 42211
rect 22278 42208 22284 42220
rect 22235 42180 22284 42208
rect 22235 42177 22247 42180
rect 22189 42171 22247 42177
rect 15933 42143 15991 42149
rect 15933 42140 15945 42143
rect 13832 42112 15240 42140
rect 15488 42112 15945 42140
rect 13832 42072 13860 42112
rect 10888 42044 12296 42072
rect 13556 42044 13860 42072
rect 12268 42016 12296 42044
rect 8386 42004 8392 42016
rect 5500 41976 8392 42004
rect 5500 41964 5506 41976
rect 8386 41964 8392 41976
rect 8444 41964 8450 42016
rect 10686 41964 10692 42016
rect 10744 41964 10750 42016
rect 11146 41964 11152 42016
rect 11204 41964 11210 42016
rect 12250 41964 12256 42016
rect 12308 42004 12314 42016
rect 14182 42004 14188 42016
rect 12308 41976 14188 42004
rect 12308 41964 12314 41976
rect 14182 41964 14188 41976
rect 14240 41964 14246 42016
rect 15286 41964 15292 42016
rect 15344 42004 15350 42016
rect 15488 42013 15516 42112
rect 15933 42109 15945 42112
rect 15979 42109 15991 42143
rect 15933 42103 15991 42109
rect 17310 42100 17316 42152
rect 17368 42100 17374 42152
rect 19150 42100 19156 42152
rect 19208 42100 19214 42152
rect 19429 42143 19487 42149
rect 19429 42109 19441 42143
rect 19475 42140 19487 42143
rect 19978 42140 19984 42152
rect 19475 42112 19984 42140
rect 19475 42109 19487 42112
rect 19429 42103 19487 42109
rect 19978 42100 19984 42112
rect 20036 42100 20042 42152
rect 20622 42100 20628 42152
rect 20680 42100 20686 42152
rect 15838 42032 15844 42084
rect 15896 42072 15902 42084
rect 21928 42072 21956 42171
rect 22278 42168 22284 42180
rect 22336 42168 22342 42220
rect 22388 42217 22416 42248
rect 23017 42245 23029 42248
rect 23063 42245 23075 42279
rect 23017 42239 23075 42245
rect 23566 42236 23572 42288
rect 23624 42236 23630 42288
rect 22373 42211 22431 42217
rect 22373 42177 22385 42211
rect 22419 42177 22431 42211
rect 22373 42171 22431 42177
rect 22646 42168 22652 42220
rect 22704 42168 22710 42220
rect 22830 42168 22836 42220
rect 22888 42208 22894 42220
rect 23106 42208 23112 42220
rect 22888 42180 23112 42208
rect 22888 42168 22894 42180
rect 23106 42168 23112 42180
rect 23164 42168 23170 42220
rect 23753 42211 23811 42217
rect 23753 42208 23765 42211
rect 23216 42180 23765 42208
rect 22664 42140 22692 42168
rect 22922 42140 22928 42152
rect 22664 42112 22928 42140
rect 22922 42100 22928 42112
rect 22980 42140 22986 42152
rect 23216 42140 23244 42180
rect 23753 42177 23765 42180
rect 23799 42177 23811 42211
rect 23860 42208 23888 42304
rect 25133 42279 25191 42285
rect 25133 42245 25145 42279
rect 25179 42276 25191 42279
rect 26326 42276 26332 42288
rect 25179 42248 26332 42276
rect 25179 42245 25191 42248
rect 25133 42239 25191 42245
rect 26326 42236 26332 42248
rect 26384 42276 26390 42288
rect 26384 42248 26740 42276
rect 26384 42236 26390 42248
rect 26712 42220 26740 42248
rect 26878 42236 26884 42288
rect 26936 42236 26942 42288
rect 23937 42211 23995 42217
rect 23937 42208 23949 42211
rect 23860 42180 23949 42208
rect 23753 42171 23811 42177
rect 23937 42177 23949 42180
rect 23983 42177 23995 42211
rect 23937 42171 23995 42177
rect 25038 42168 25044 42220
rect 25096 42168 25102 42220
rect 26142 42168 26148 42220
rect 26200 42208 26206 42220
rect 26605 42211 26663 42217
rect 26605 42208 26617 42211
rect 26200 42180 26617 42208
rect 26200 42168 26206 42180
rect 26605 42177 26617 42180
rect 26651 42177 26663 42211
rect 26605 42171 26663 42177
rect 22980 42112 23244 42140
rect 22980 42100 22986 42112
rect 23290 42100 23296 42152
rect 23348 42140 23354 42152
rect 23569 42143 23627 42149
rect 23569 42140 23581 42143
rect 23348 42112 23581 42140
rect 23348 42100 23354 42112
rect 23569 42109 23581 42112
rect 23615 42109 23627 42143
rect 23569 42103 23627 42109
rect 25317 42143 25375 42149
rect 25317 42109 25329 42143
rect 25363 42140 25375 42143
rect 26160 42140 26188 42168
rect 25363 42112 26188 42140
rect 26620 42140 26648 42171
rect 26694 42168 26700 42220
rect 26752 42168 26758 42220
rect 26789 42211 26847 42217
rect 26789 42177 26801 42211
rect 26835 42208 26847 42211
rect 26896 42208 26924 42236
rect 26988 42217 27016 42316
rect 28534 42276 28540 42288
rect 28474 42248 28540 42276
rect 28534 42236 28540 42248
rect 28592 42236 28598 42288
rect 28828 42217 28856 42316
rect 30484 42316 31484 42344
rect 30374 42276 30380 42288
rect 30314 42248 30380 42276
rect 30374 42236 30380 42248
rect 30432 42276 30438 42288
rect 30484 42276 30512 42316
rect 31478 42304 31484 42316
rect 31536 42344 31542 42356
rect 31662 42344 31668 42356
rect 31536 42316 31668 42344
rect 31536 42304 31542 42316
rect 31662 42304 31668 42316
rect 31720 42304 31726 42356
rect 31754 42304 31760 42356
rect 31812 42304 31818 42356
rect 32582 42304 32588 42356
rect 32640 42344 32646 42356
rect 33778 42344 33784 42356
rect 32640 42316 33784 42344
rect 32640 42304 32646 42316
rect 30432 42248 30512 42276
rect 30432 42236 30438 42248
rect 30558 42236 30564 42288
rect 30616 42276 30622 42288
rect 33226 42276 33232 42288
rect 30616 42248 33232 42276
rect 30616 42236 30622 42248
rect 33226 42236 33232 42248
rect 33284 42276 33290 42288
rect 33612 42285 33640 42316
rect 33778 42304 33784 42316
rect 33836 42304 33842 42356
rect 33965 42347 34023 42353
rect 33965 42313 33977 42347
rect 34011 42344 34023 42347
rect 34238 42344 34244 42356
rect 34011 42316 34244 42344
rect 34011 42313 34023 42316
rect 33965 42307 34023 42313
rect 34238 42304 34244 42316
rect 34296 42304 34302 42356
rect 34882 42304 34888 42356
rect 34940 42304 34946 42356
rect 33459 42279 33517 42285
rect 33459 42276 33471 42279
rect 33284 42248 33471 42276
rect 33284 42236 33290 42248
rect 33459 42245 33471 42248
rect 33505 42245 33517 42279
rect 33459 42239 33517 42245
rect 33597 42279 33655 42285
rect 33597 42245 33609 42279
rect 33643 42245 33655 42279
rect 33597 42239 33655 42245
rect 33686 42236 33692 42288
rect 33744 42236 33750 42288
rect 34146 42276 34152 42288
rect 33796 42248 34152 42276
rect 26835 42180 26924 42208
rect 26835 42177 26847 42180
rect 26789 42171 26847 42177
rect 26620 42112 26832 42140
rect 25363 42109 25375 42112
rect 25317 42103 25375 42109
rect 26804 42084 26832 42112
rect 23753 42075 23811 42081
rect 23753 42072 23765 42075
rect 15896 42044 16574 42072
rect 21928 42044 23765 42072
rect 15896 42032 15902 42044
rect 15473 42007 15531 42013
rect 15473 42004 15485 42007
rect 15344 41976 15485 42004
rect 15344 41964 15350 41976
rect 15473 41973 15485 41976
rect 15519 41973 15531 42007
rect 16546 42004 16574 42044
rect 23753 42041 23765 42044
rect 23799 42041 23811 42075
rect 23753 42035 23811 42041
rect 26786 42032 26792 42084
rect 26844 42032 26850 42084
rect 18966 42004 18972 42016
rect 16546 41976 18972 42004
rect 15473 41967 15531 41973
rect 18966 41964 18972 41976
rect 19024 41964 19030 42016
rect 19061 42007 19119 42013
rect 19061 41973 19073 42007
rect 19107 42004 19119 42007
rect 20530 42004 20536 42016
rect 19107 41976 20536 42004
rect 19107 41973 19119 41976
rect 19061 41967 19119 41973
rect 20530 41964 20536 41976
rect 20588 41964 20594 42016
rect 22186 41964 22192 42016
rect 22244 41964 22250 42016
rect 22278 41964 22284 42016
rect 22336 42004 22342 42016
rect 22465 42007 22523 42013
rect 22465 42004 22477 42007
rect 22336 41976 22477 42004
rect 22336 41964 22342 41976
rect 22465 41973 22477 41976
rect 22511 42004 22523 42007
rect 22830 42004 22836 42016
rect 22511 41976 22836 42004
rect 22511 41973 22523 41976
rect 22465 41967 22523 41973
rect 22830 41964 22836 41976
rect 22888 41964 22894 42016
rect 26694 41964 26700 42016
rect 26752 41964 26758 42016
rect 26896 42004 26924 42180
rect 26973 42211 27031 42217
rect 26973 42177 26985 42211
rect 27019 42177 27031 42211
rect 26973 42171 27031 42177
rect 28813 42211 28871 42217
rect 28813 42177 28825 42211
rect 28859 42177 28871 42211
rect 28813 42171 28871 42177
rect 30650 42168 30656 42220
rect 30708 42208 30714 42220
rect 31573 42211 31631 42217
rect 31573 42208 31585 42211
rect 30708 42180 31585 42208
rect 30708 42168 30714 42180
rect 31573 42177 31585 42180
rect 31619 42177 31631 42211
rect 31573 42171 31631 42177
rect 27246 42100 27252 42152
rect 27304 42100 27310 42152
rect 29086 42100 29092 42152
rect 29144 42100 29150 42152
rect 30561 42143 30619 42149
rect 30561 42140 30573 42143
rect 30208 42112 30573 42140
rect 30208 42084 30236 42112
rect 30561 42109 30573 42112
rect 30607 42140 30619 42143
rect 31205 42143 31263 42149
rect 31205 42140 31217 42143
rect 30607 42112 31217 42140
rect 30607 42109 30619 42112
rect 30561 42103 30619 42109
rect 31205 42109 31217 42112
rect 31251 42109 31263 42143
rect 31588 42140 31616 42171
rect 31846 42168 31852 42220
rect 31904 42168 31910 42220
rect 32125 42211 32183 42217
rect 32125 42177 32137 42211
rect 32171 42177 32183 42211
rect 32125 42171 32183 42177
rect 32309 42211 32367 42217
rect 32309 42177 32321 42211
rect 32355 42177 32367 42211
rect 32309 42171 32367 42177
rect 31662 42140 31668 42152
rect 31588 42112 31668 42140
rect 31205 42103 31263 42109
rect 31662 42100 31668 42112
rect 31720 42140 31726 42152
rect 32140 42140 32168 42171
rect 31720 42112 32168 42140
rect 31720 42100 31726 42112
rect 30190 42032 30196 42084
rect 30248 42032 30254 42084
rect 30466 42032 30472 42084
rect 30524 42072 30530 42084
rect 31389 42075 31447 42081
rect 31389 42072 31401 42075
rect 30524 42044 31401 42072
rect 30524 42032 30530 42044
rect 31389 42041 31401 42044
rect 31435 42041 31447 42075
rect 32324 42072 32352 42171
rect 33318 42168 33324 42220
rect 33376 42168 33382 42220
rect 33796 42217 33824 42248
rect 34146 42236 34152 42248
rect 34204 42276 34210 42288
rect 34204 42248 34376 42276
rect 34204 42236 34210 42248
rect 33781 42211 33839 42217
rect 33781 42177 33793 42211
rect 33827 42177 33839 42211
rect 33781 42171 33839 42177
rect 34241 42211 34299 42217
rect 34241 42177 34253 42211
rect 34287 42177 34299 42211
rect 34348 42208 34376 42248
rect 34698 42236 34704 42288
rect 34756 42236 34762 42288
rect 34790 42236 34796 42288
rect 34848 42276 34854 42288
rect 34848 42248 35020 42276
rect 34848 42236 34854 42248
rect 34992 42217 35020 42248
rect 34885 42211 34943 42217
rect 34885 42208 34897 42211
rect 34348 42180 34897 42208
rect 34241 42171 34299 42177
rect 34885 42177 34897 42180
rect 34931 42177 34943 42211
rect 34885 42171 34943 42177
rect 34977 42211 35035 42217
rect 34977 42177 34989 42211
rect 35023 42177 35035 42211
rect 34977 42171 35035 42177
rect 34149 42143 34207 42149
rect 34149 42140 34161 42143
rect 31389 42035 31447 42041
rect 31680 42044 32352 42072
rect 32784 42112 34161 42140
rect 28350 42004 28356 42016
rect 26896 41976 28356 42004
rect 28350 41964 28356 41976
rect 28408 42004 28414 42016
rect 28721 42007 28779 42013
rect 28721 42004 28733 42007
rect 28408 41976 28733 42004
rect 28408 41964 28414 41976
rect 28721 41973 28733 41976
rect 28767 41973 28779 42007
rect 28721 41967 28779 41973
rect 30650 41964 30656 42016
rect 30708 41964 30714 42016
rect 31202 41964 31208 42016
rect 31260 42004 31266 42016
rect 31680 42004 31708 42044
rect 32784 42016 32812 42112
rect 34149 42109 34161 42112
rect 34195 42109 34207 42143
rect 34256 42140 34284 42171
rect 35250 42168 35256 42220
rect 35308 42168 35314 42220
rect 35268 42140 35296 42168
rect 34256 42112 35296 42140
rect 34149 42103 34207 42109
rect 31260 41976 31708 42004
rect 31260 41964 31266 41976
rect 31754 41964 31760 42016
rect 31812 42004 31818 42016
rect 32125 42007 32183 42013
rect 32125 42004 32137 42007
rect 31812 41976 32137 42004
rect 31812 41964 31818 41976
rect 32125 41973 32137 41976
rect 32171 41973 32183 42007
rect 32125 41967 32183 41973
rect 32766 41964 32772 42016
rect 32824 41964 32830 42016
rect 33502 41964 33508 42016
rect 33560 42004 33566 42016
rect 34440 42004 34468 42112
rect 34609 42075 34667 42081
rect 34609 42041 34621 42075
rect 34655 42072 34667 42075
rect 34698 42072 34704 42084
rect 34655 42044 34704 42072
rect 34655 42041 34667 42044
rect 34609 42035 34667 42041
rect 34698 42032 34704 42044
rect 34756 42032 34762 42084
rect 33560 41976 34468 42004
rect 33560 41964 33566 41976
rect 1104 41914 45172 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 45172 41914
rect 1104 41840 45172 41862
rect 3605 41803 3663 41809
rect 3605 41769 3617 41803
rect 3651 41800 3663 41803
rect 3878 41800 3884 41812
rect 3651 41772 3884 41800
rect 3651 41769 3663 41772
rect 3605 41763 3663 41769
rect 3878 41760 3884 41772
rect 3936 41760 3942 41812
rect 4614 41760 4620 41812
rect 4672 41760 4678 41812
rect 4890 41760 4896 41812
rect 4948 41800 4954 41812
rect 4985 41803 5043 41809
rect 4985 41800 4997 41803
rect 4948 41772 4997 41800
rect 4948 41760 4954 41772
rect 4985 41769 4997 41772
rect 5031 41769 5043 41803
rect 4985 41763 5043 41769
rect 5350 41760 5356 41812
rect 5408 41760 5414 41812
rect 6362 41760 6368 41812
rect 6420 41800 6426 41812
rect 6457 41803 6515 41809
rect 6457 41800 6469 41803
rect 6420 41772 6469 41800
rect 6420 41760 6426 41772
rect 6457 41769 6469 41772
rect 6503 41769 6515 41803
rect 6457 41763 6515 41769
rect 8294 41760 8300 41812
rect 8352 41760 8358 41812
rect 8754 41760 8760 41812
rect 8812 41760 8818 41812
rect 10778 41800 10784 41812
rect 8864 41772 10784 41800
rect 4338 41732 4344 41744
rect 3804 41704 4344 41732
rect 2133 41667 2191 41673
rect 2133 41633 2145 41667
rect 2179 41664 2191 41667
rect 2774 41664 2780 41676
rect 2179 41636 2780 41664
rect 2179 41633 2191 41636
rect 2133 41627 2191 41633
rect 2774 41624 2780 41636
rect 2832 41624 2838 41676
rect 3326 41624 3332 41676
rect 3384 41624 3390 41676
rect 3804 41673 3832 41704
rect 4338 41692 4344 41704
rect 4396 41692 4402 41744
rect 3789 41667 3847 41673
rect 3789 41633 3801 41667
rect 3835 41633 3847 41667
rect 4632 41664 4660 41760
rect 4798 41732 4804 41744
rect 3789 41627 3847 41633
rect 4356 41636 4660 41664
rect 4724 41704 4804 41732
rect 1854 41556 1860 41608
rect 1912 41556 1918 41608
rect 3344 41596 3372 41624
rect 4356 41605 4384 41636
rect 3266 41568 3372 41596
rect 3973 41599 4031 41605
rect 3973 41565 3985 41599
rect 4019 41596 4031 41599
rect 4341 41599 4399 41605
rect 4019 41568 4292 41596
rect 4019 41565 4031 41568
rect 3973 41559 4031 41565
rect 4264 41540 4292 41568
rect 4341 41565 4353 41599
rect 4387 41565 4399 41599
rect 4341 41559 4399 41565
rect 4489 41599 4547 41605
rect 4489 41565 4501 41599
rect 4535 41596 4547 41599
rect 4724 41596 4752 41704
rect 4798 41692 4804 41704
rect 4856 41692 4862 41744
rect 5368 41673 5396 41760
rect 7745 41735 7803 41741
rect 7745 41701 7757 41735
rect 7791 41732 7803 41735
rect 8772 41732 8800 41760
rect 7791 41704 8800 41732
rect 7791 41701 7803 41704
rect 7745 41695 7803 41701
rect 5353 41667 5411 41673
rect 5353 41633 5365 41667
rect 5399 41633 5411 41667
rect 5353 41627 5411 41633
rect 5442 41624 5448 41676
rect 5500 41664 5506 41676
rect 5500 41636 6316 41664
rect 5500 41624 5506 41636
rect 4535 41565 4568 41596
rect 4489 41559 4568 41565
rect 4246 41488 4252 41540
rect 4304 41488 4310 41540
rect 4154 41420 4160 41472
rect 4212 41420 4218 41472
rect 4540 41460 4568 41559
rect 4632 41568 4752 41596
rect 4847 41599 4905 41605
rect 4632 41537 4660 41568
rect 4847 41565 4859 41599
rect 4893 41596 4905 41599
rect 4982 41596 4988 41608
rect 4893 41568 4988 41596
rect 4893 41565 4905 41568
rect 4847 41559 4905 41565
rect 4982 41556 4988 41568
rect 5040 41596 5046 41608
rect 5534 41596 5540 41608
rect 5040 41568 5540 41596
rect 5040 41556 5046 41568
rect 5534 41556 5540 41568
rect 5592 41556 5598 41608
rect 6288 41605 6316 41636
rect 6454 41624 6460 41676
rect 6512 41664 6518 41676
rect 7377 41667 7435 41673
rect 7377 41664 7389 41667
rect 6512 41636 7389 41664
rect 6512 41624 6518 41636
rect 7377 41633 7389 41636
rect 7423 41633 7435 41667
rect 8864 41664 8892 41772
rect 10778 41760 10784 41772
rect 10836 41760 10842 41812
rect 11146 41760 11152 41812
rect 11204 41760 11210 41812
rect 11514 41760 11520 41812
rect 11572 41760 11578 41812
rect 11698 41760 11704 41812
rect 11756 41760 11762 41812
rect 12253 41803 12311 41809
rect 12253 41769 12265 41803
rect 12299 41800 12311 41803
rect 12802 41800 12808 41812
rect 12299 41772 12808 41800
rect 12299 41769 12311 41772
rect 12253 41763 12311 41769
rect 12802 41760 12808 41772
rect 12860 41760 12866 41812
rect 13081 41803 13139 41809
rect 13081 41769 13093 41803
rect 13127 41800 13139 41803
rect 13354 41800 13360 41812
rect 13127 41772 13360 41800
rect 13127 41769 13139 41772
rect 13081 41763 13139 41769
rect 13354 41760 13360 41772
rect 13412 41760 13418 41812
rect 17310 41760 17316 41812
rect 17368 41760 17374 41812
rect 18506 41760 18512 41812
rect 18564 41760 18570 41812
rect 18782 41760 18788 41812
rect 18840 41800 18846 41812
rect 19061 41803 19119 41809
rect 19061 41800 19073 41803
rect 18840 41772 19073 41800
rect 18840 41760 18846 41772
rect 19061 41769 19073 41772
rect 19107 41769 19119 41803
rect 19061 41763 19119 41769
rect 19245 41803 19303 41809
rect 19245 41769 19257 41803
rect 19291 41800 19303 41803
rect 19334 41800 19340 41812
rect 19291 41772 19340 41800
rect 19291 41769 19303 41772
rect 19245 41763 19303 41769
rect 19334 41760 19340 41772
rect 19392 41760 19398 41812
rect 19981 41803 20039 41809
rect 19536 41772 19932 41800
rect 7377 41627 7435 41633
rect 7576 41636 8892 41664
rect 9493 41667 9551 41673
rect 7576 41605 7604 41636
rect 9493 41633 9505 41667
rect 9539 41633 9551 41667
rect 9493 41627 9551 41633
rect 6089 41599 6147 41605
rect 6089 41596 6101 41599
rect 6012 41568 6101 41596
rect 4617 41531 4675 41537
rect 4617 41497 4629 41531
rect 4663 41497 4675 41531
rect 4617 41491 4675 41497
rect 4709 41531 4767 41537
rect 4709 41497 4721 41531
rect 4755 41528 4767 41531
rect 5258 41528 5264 41540
rect 4755 41500 5264 41528
rect 4755 41497 4767 41500
rect 4709 41491 4767 41497
rect 5258 41488 5264 41500
rect 5316 41488 5322 41540
rect 6012 41469 6040 41568
rect 6089 41565 6101 41568
rect 6135 41565 6147 41599
rect 6089 41559 6147 41565
rect 6273 41599 6331 41605
rect 6273 41565 6285 41599
rect 6319 41596 6331 41599
rect 7561 41599 7619 41605
rect 7561 41596 7573 41599
rect 6319 41568 7573 41596
rect 6319 41565 6331 41568
rect 6273 41559 6331 41565
rect 7561 41565 7573 41568
rect 7607 41565 7619 41599
rect 7561 41559 7619 41565
rect 8481 41599 8539 41605
rect 8481 41565 8493 41599
rect 8527 41596 8539 41599
rect 8527 41568 8984 41596
rect 8527 41565 8539 41568
rect 8481 41559 8539 41565
rect 8956 41469 8984 41568
rect 9122 41488 9128 41540
rect 9180 41528 9186 41540
rect 9508 41528 9536 41627
rect 10137 41599 10195 41605
rect 10137 41565 10149 41599
rect 10183 41596 10195 41599
rect 11164 41596 11192 41760
rect 11716 41605 11744 41760
rect 11790 41692 11796 41744
rect 11848 41732 11854 41744
rect 18524 41732 18552 41760
rect 19536 41732 19564 41772
rect 11848 41704 12204 41732
rect 11848 41692 11854 41704
rect 11882 41624 11888 41676
rect 11940 41624 11946 41676
rect 12176 41664 12204 41704
rect 12406 41704 13768 41732
rect 18524 41704 19564 41732
rect 12406 41664 12434 41704
rect 12176 41636 12434 41664
rect 11609 41599 11667 41605
rect 11609 41596 11621 41599
rect 10183 41568 11100 41596
rect 11164 41568 11621 41596
rect 10183 41565 10195 41568
rect 10137 41559 10195 41565
rect 11072 41540 11100 41568
rect 11609 41565 11621 41568
rect 11655 41565 11667 41599
rect 11609 41559 11667 41565
rect 11702 41599 11760 41605
rect 11702 41565 11714 41599
rect 11748 41565 11760 41599
rect 11900 41596 11928 41624
rect 11977 41599 12035 41605
rect 11977 41596 11989 41599
rect 11900 41568 11989 41596
rect 11702 41559 11760 41565
rect 11977 41565 11989 41568
rect 12023 41565 12035 41599
rect 11977 41559 12035 41565
rect 12074 41599 12132 41605
rect 12074 41565 12086 41599
rect 12120 41596 12132 41599
rect 12176 41596 12204 41636
rect 13630 41624 13636 41676
rect 13688 41624 13694 41676
rect 13740 41664 13768 41704
rect 19794 41692 19800 41744
rect 19852 41692 19858 41744
rect 14274 41664 14280 41676
rect 13740 41636 14280 41664
rect 14274 41624 14280 41636
rect 14332 41664 14338 41676
rect 14332 41636 16068 41664
rect 14332 41624 14338 41636
rect 12120 41568 12204 41596
rect 12120 41565 12132 41568
rect 12074 41559 12132 41565
rect 12250 41556 12256 41608
rect 12308 41556 12314 41608
rect 13449 41599 13507 41605
rect 13449 41565 13461 41599
rect 13495 41596 13507 41599
rect 14550 41596 14556 41608
rect 13495 41568 14556 41596
rect 13495 41565 13507 41568
rect 13449 41559 13507 41565
rect 14550 41556 14556 41568
rect 14608 41556 14614 41608
rect 15933 41599 15991 41605
rect 15933 41565 15945 41599
rect 15979 41565 15991 41599
rect 16040 41596 16068 41636
rect 18322 41624 18328 41676
rect 18380 41664 18386 41676
rect 18417 41667 18475 41673
rect 18417 41664 18429 41667
rect 18380 41636 18429 41664
rect 18380 41624 18386 41636
rect 18417 41633 18429 41636
rect 18463 41633 18475 41667
rect 18417 41627 18475 41633
rect 16482 41596 16488 41608
rect 16040 41568 16488 41596
rect 15933 41559 15991 41565
rect 9180 41500 9536 41528
rect 9180 41488 9186 41500
rect 5997 41463 6055 41469
rect 5997 41460 6009 41463
rect 4540 41432 6009 41460
rect 5997 41429 6009 41432
rect 6043 41429 6055 41463
rect 5997 41423 6055 41429
rect 8941 41463 8999 41469
rect 8941 41429 8953 41463
rect 8987 41429 8999 41463
rect 8941 41423 8999 41429
rect 9306 41420 9312 41472
rect 9364 41420 9370 41472
rect 9398 41420 9404 41472
rect 9456 41420 9462 41472
rect 9508 41460 9536 41500
rect 10404 41531 10462 41537
rect 10404 41497 10416 41531
rect 10450 41528 10462 41531
rect 10502 41528 10508 41540
rect 10450 41500 10508 41528
rect 10450 41497 10462 41500
rect 10404 41491 10462 41497
rect 10502 41488 10508 41500
rect 10560 41488 10566 41540
rect 11054 41488 11060 41540
rect 11112 41488 11118 41540
rect 11885 41531 11943 41537
rect 11885 41497 11897 41531
rect 11931 41528 11943 41531
rect 12268 41528 12296 41556
rect 11931 41500 12296 41528
rect 14093 41531 14151 41537
rect 11931 41497 11943 41500
rect 11885 41491 11943 41497
rect 14093 41497 14105 41531
rect 14139 41528 14151 41531
rect 15470 41528 15476 41540
rect 14139 41500 15476 41528
rect 14139 41497 14151 41500
rect 14093 41491 14151 41497
rect 15470 41488 15476 41500
rect 15528 41488 15534 41540
rect 11238 41460 11244 41472
rect 9508 41432 11244 41460
rect 11238 41420 11244 41432
rect 11296 41420 11302 41472
rect 13354 41420 13360 41472
rect 13412 41460 13418 41472
rect 13541 41463 13599 41469
rect 13541 41460 13553 41463
rect 13412 41432 13553 41460
rect 13412 41420 13418 41432
rect 13541 41429 13553 41432
rect 13587 41429 13599 41463
rect 13541 41423 13599 41429
rect 13722 41420 13728 41472
rect 13780 41460 13786 41472
rect 15378 41460 15384 41472
rect 13780 41432 15384 41460
rect 13780 41420 13786 41432
rect 15378 41420 15384 41432
rect 15436 41460 15442 41472
rect 15948 41460 15976 41559
rect 16482 41556 16488 41568
rect 16540 41596 16546 41608
rect 18782 41596 18788 41608
rect 16540 41568 18788 41596
rect 16540 41556 16546 41568
rect 18782 41556 18788 41568
rect 18840 41596 18846 41608
rect 19812 41605 19840 41692
rect 19904 41605 19932 41772
rect 19981 41769 19993 41803
rect 20027 41800 20039 41803
rect 20070 41800 20076 41812
rect 20027 41772 20076 41800
rect 20027 41769 20039 41772
rect 19981 41763 20039 41769
rect 19383 41599 19441 41605
rect 19383 41596 19395 41599
rect 18840 41568 19395 41596
rect 18840 41556 18846 41568
rect 19383 41565 19395 41568
rect 19429 41565 19441 41599
rect 19383 41559 19441 41565
rect 19521 41599 19579 41605
rect 19521 41565 19533 41599
rect 19567 41596 19579 41599
rect 19796 41599 19854 41605
rect 19567 41568 19748 41596
rect 19567 41565 19579 41568
rect 19521 41559 19579 41565
rect 16022 41488 16028 41540
rect 16080 41528 16086 41540
rect 16178 41531 16236 41537
rect 16178 41528 16190 41531
rect 16080 41500 16190 41528
rect 16080 41488 16086 41500
rect 16178 41497 16190 41500
rect 16224 41497 16236 41531
rect 16178 41491 16236 41497
rect 18693 41531 18751 41537
rect 18693 41497 18705 41531
rect 18739 41528 18751 41531
rect 19536 41528 19564 41559
rect 18739 41500 19564 41528
rect 19613 41531 19671 41537
rect 18739 41497 18751 41500
rect 18693 41491 18751 41497
rect 19613 41497 19625 41531
rect 19659 41497 19671 41531
rect 19720 41528 19748 41568
rect 19796 41565 19808 41599
rect 19842 41565 19854 41599
rect 19796 41559 19854 41565
rect 19889 41599 19947 41605
rect 19889 41565 19901 41599
rect 19935 41565 19947 41599
rect 19889 41559 19947 41565
rect 19996 41528 20024 41763
rect 20070 41760 20076 41772
rect 20128 41760 20134 41812
rect 20530 41760 20536 41812
rect 20588 41760 20594 41812
rect 23201 41803 23259 41809
rect 23201 41769 23213 41803
rect 23247 41800 23259 41803
rect 23290 41800 23296 41812
rect 23247 41772 23296 41800
rect 23247 41769 23259 41772
rect 23201 41763 23259 41769
rect 20548 41673 20576 41760
rect 22925 41735 22983 41741
rect 22925 41701 22937 41735
rect 22971 41732 22983 41735
rect 23216 41732 23244 41763
rect 23290 41760 23296 41772
rect 23348 41760 23354 41812
rect 26694 41760 26700 41812
rect 26752 41760 26758 41812
rect 26789 41803 26847 41809
rect 26789 41769 26801 41803
rect 26835 41800 26847 41803
rect 27246 41800 27252 41812
rect 26835 41772 27252 41800
rect 26835 41769 26847 41772
rect 26789 41763 26847 41769
rect 27246 41760 27252 41772
rect 27304 41760 27310 41812
rect 29086 41760 29092 41812
rect 29144 41800 29150 41812
rect 29549 41803 29607 41809
rect 29549 41800 29561 41803
rect 29144 41772 29561 41800
rect 29144 41760 29150 41772
rect 29549 41769 29561 41772
rect 29595 41769 29607 41803
rect 29549 41763 29607 41769
rect 29822 41760 29828 41812
rect 29880 41800 29886 41812
rect 30374 41800 30380 41812
rect 29880 41772 30380 41800
rect 29880 41760 29886 41772
rect 30374 41760 30380 41772
rect 30432 41760 30438 41812
rect 30466 41760 30472 41812
rect 30524 41760 30530 41812
rect 30650 41760 30656 41812
rect 30708 41760 30714 41812
rect 30834 41760 30840 41812
rect 30892 41800 30898 41812
rect 30929 41803 30987 41809
rect 30929 41800 30941 41803
rect 30892 41772 30941 41800
rect 30892 41760 30898 41772
rect 30929 41769 30941 41772
rect 30975 41769 30987 41803
rect 31481 41803 31539 41809
rect 31481 41800 31493 41803
rect 30929 41763 30987 41769
rect 31036 41772 31493 41800
rect 22971 41704 23244 41732
rect 22971 41701 22983 41704
rect 22925 41695 22983 41701
rect 20533 41667 20591 41673
rect 20533 41633 20545 41667
rect 20579 41633 20591 41667
rect 23382 41664 23388 41676
rect 20533 41627 20591 41633
rect 23032 41636 23388 41664
rect 20714 41556 20720 41608
rect 20772 41596 20778 41608
rect 21174 41596 21180 41608
rect 20772 41568 21180 41596
rect 20772 41556 20778 41568
rect 21174 41556 21180 41568
rect 21232 41556 21238 41608
rect 23032 41596 23060 41636
rect 23382 41624 23388 41636
rect 23440 41664 23446 41676
rect 23934 41664 23940 41676
rect 23440 41636 23940 41664
rect 23440 41624 23446 41636
rect 23934 41624 23940 41636
rect 23992 41624 23998 41676
rect 26712 41664 26740 41760
rect 30484 41732 30512 41760
rect 30668 41732 30696 41760
rect 31036 41732 31064 41772
rect 31481 41769 31493 41772
rect 31527 41800 31539 41803
rect 31846 41800 31852 41812
rect 31527 41772 31852 41800
rect 31527 41769 31539 41772
rect 31481 41763 31539 41769
rect 31846 41760 31852 41772
rect 31904 41760 31910 41812
rect 32309 41803 32367 41809
rect 32309 41769 32321 41803
rect 32355 41800 32367 41803
rect 32355 41772 32996 41800
rect 32355 41769 32367 41772
rect 32309 41763 32367 41769
rect 32861 41735 32919 41741
rect 32861 41732 32873 41735
rect 30024 41704 30512 41732
rect 30576 41704 30696 41732
rect 30760 41704 31064 41732
rect 31128 41704 32873 41732
rect 26712 41636 27200 41664
rect 22586 41568 23060 41596
rect 23106 41556 23112 41608
rect 23164 41556 23170 41608
rect 23198 41556 23204 41608
rect 23256 41556 23262 41608
rect 23474 41556 23480 41608
rect 23532 41596 23538 41608
rect 24581 41599 24639 41605
rect 24581 41596 24593 41599
rect 23532 41568 24593 41596
rect 23532 41556 23538 41568
rect 24581 41565 24593 41568
rect 24627 41565 24639 41599
rect 24581 41559 24639 41565
rect 26970 41556 26976 41608
rect 27028 41556 27034 41608
rect 27172 41605 27200 41636
rect 28350 41624 28356 41676
rect 28408 41624 28414 41676
rect 30024 41664 30052 41704
rect 29840 41636 30052 41664
rect 29750 41609 29808 41615
rect 27157 41599 27215 41605
rect 27157 41565 27169 41599
rect 27203 41565 27215 41599
rect 27157 41559 27215 41565
rect 27433 41599 27491 41605
rect 27433 41565 27445 41599
rect 27479 41596 27491 41599
rect 27801 41599 27859 41605
rect 27801 41596 27813 41599
rect 27479 41568 27813 41596
rect 27479 41565 27491 41568
rect 27433 41559 27491 41565
rect 27801 41565 27813 41568
rect 27847 41565 27859 41599
rect 29750 41575 29762 41609
rect 29796 41606 29808 41609
rect 29840 41606 29868 41636
rect 30098 41624 30104 41676
rect 30156 41624 30162 41676
rect 30193 41667 30251 41673
rect 30193 41633 30205 41667
rect 30239 41664 30251 41667
rect 30576 41664 30604 41704
rect 30760 41664 30788 41704
rect 30239 41636 30604 41664
rect 30668 41636 30788 41664
rect 30239 41633 30251 41636
rect 30193 41627 30251 41633
rect 29796 41578 29868 41606
rect 29917 41599 29975 41605
rect 29796 41575 29808 41578
rect 29750 41569 29808 41575
rect 27801 41559 27859 41565
rect 29917 41565 29929 41599
rect 29963 41596 29975 41599
rect 30116 41596 30144 41624
rect 29963 41568 30144 41596
rect 29963 41565 29975 41568
rect 29917 41559 29975 41565
rect 30282 41556 30288 41608
rect 30340 41596 30346 41608
rect 30377 41599 30435 41605
rect 30377 41596 30389 41599
rect 30340 41568 30389 41596
rect 30340 41556 30346 41568
rect 30377 41565 30389 41568
rect 30423 41565 30435 41599
rect 30377 41559 30435 41565
rect 30561 41599 30619 41605
rect 30561 41565 30573 41599
rect 30607 41596 30619 41599
rect 30668 41596 30696 41636
rect 30926 41624 30932 41676
rect 30984 41664 30990 41676
rect 31128 41664 31156 41704
rect 32861 41701 32873 41704
rect 32907 41701 32919 41735
rect 32861 41695 32919 41701
rect 30984 41636 31156 41664
rect 30984 41624 30990 41636
rect 30607 41568 30696 41596
rect 30607 41565 30619 41568
rect 30561 41559 30619 41565
rect 30742 41556 30748 41608
rect 30800 41556 30806 41608
rect 31128 41605 31156 41636
rect 31662 41624 31668 41676
rect 31720 41624 31726 41676
rect 31938 41624 31944 41676
rect 31996 41624 32002 41676
rect 32766 41672 32772 41676
rect 32324 41664 32536 41672
rect 32692 41664 32772 41672
rect 32232 41644 32772 41664
rect 32232 41636 32352 41644
rect 32508 41636 32720 41644
rect 31021 41599 31079 41605
rect 31021 41565 31033 41599
rect 31067 41565 31079 41599
rect 31021 41559 31079 41565
rect 31113 41599 31171 41605
rect 31113 41565 31125 41599
rect 31159 41565 31171 41599
rect 31113 41559 31171 41565
rect 19720 41500 20024 41528
rect 19613 41491 19671 41497
rect 15436 41432 15976 41460
rect 15436 41420 15442 41432
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 18601 41463 18659 41469
rect 18601 41460 18613 41463
rect 18012 41432 18613 41460
rect 18012 41420 18018 41432
rect 18601 41429 18613 41432
rect 18647 41429 18659 41463
rect 18601 41423 18659 41429
rect 18966 41420 18972 41472
rect 19024 41460 19030 41472
rect 19628 41460 19656 41491
rect 21450 41488 21456 41540
rect 21508 41488 21514 41540
rect 22738 41488 22744 41540
rect 22796 41488 22802 41540
rect 22922 41488 22928 41540
rect 22980 41488 22986 41540
rect 23017 41531 23075 41537
rect 23017 41497 23029 41531
rect 23063 41528 23075 41531
rect 23124 41528 23152 41556
rect 23063 41500 23152 41528
rect 23216 41528 23244 41556
rect 27065 41531 27123 41537
rect 27065 41528 27077 41531
rect 23216 41500 23428 41528
rect 23063 41497 23075 41500
rect 23017 41491 23075 41497
rect 22756 41460 22784 41488
rect 19024 41432 22784 41460
rect 22940 41460 22968 41488
rect 23400 41469 23428 41500
rect 26206 41500 27077 41528
rect 26206 41472 26234 41500
rect 27065 41497 27077 41500
rect 27111 41528 27123 41531
rect 27111 41500 27200 41528
rect 27111 41497 27123 41500
rect 27065 41491 27123 41497
rect 23217 41463 23275 41469
rect 23217 41460 23229 41463
rect 22940 41432 23229 41460
rect 19024 41420 19030 41432
rect 23217 41429 23229 41432
rect 23263 41429 23275 41463
rect 23217 41423 23275 41429
rect 23385 41463 23443 41469
rect 23385 41429 23397 41463
rect 23431 41429 23443 41463
rect 23385 41423 23443 41429
rect 24857 41463 24915 41469
rect 24857 41429 24869 41463
rect 24903 41460 24915 41463
rect 25038 41460 25044 41472
rect 24903 41432 25044 41460
rect 24903 41429 24915 41432
rect 24857 41423 24915 41429
rect 25038 41420 25044 41432
rect 25096 41460 25102 41472
rect 26142 41460 26148 41472
rect 25096 41432 26148 41460
rect 25096 41420 25102 41432
rect 26142 41420 26148 41432
rect 26200 41432 26234 41472
rect 27172 41460 27200 41500
rect 27246 41488 27252 41540
rect 27304 41537 27310 41540
rect 27304 41531 27353 41537
rect 27304 41497 27307 41531
rect 27341 41528 27353 41531
rect 27341 41500 29776 41528
rect 27341 41497 27353 41500
rect 27304 41491 27353 41497
rect 27304 41488 27310 41491
rect 29638 41460 29644 41472
rect 27172 41432 29644 41460
rect 26200 41420 26206 41432
rect 29638 41420 29644 41432
rect 29696 41420 29702 41472
rect 29748 41460 29776 41500
rect 29822 41488 29828 41540
rect 29880 41537 29886 41540
rect 29880 41531 29894 41537
rect 29882 41528 29894 41531
rect 30055 41531 30113 41537
rect 29882 41500 29925 41528
rect 29882 41497 29894 41500
rect 29880 41491 29894 41497
rect 30055 41497 30067 41531
rect 30101 41528 30113 41531
rect 30466 41528 30472 41540
rect 30101 41500 30472 41528
rect 30101 41497 30113 41500
rect 30055 41491 30113 41497
rect 29880 41488 29886 41491
rect 30070 41460 30098 41491
rect 30466 41488 30472 41500
rect 30524 41488 30530 41540
rect 30650 41488 30656 41540
rect 30708 41488 30714 41540
rect 31036 41528 31064 41559
rect 31202 41556 31208 41608
rect 31260 41596 31266 41608
rect 31297 41599 31355 41605
rect 31297 41596 31309 41599
rect 31260 41568 31309 41596
rect 31260 41556 31266 41568
rect 31297 41565 31309 41568
rect 31343 41565 31355 41599
rect 31297 41559 31355 41565
rect 31570 41556 31576 41608
rect 31628 41556 31634 41608
rect 31680 41596 31708 41624
rect 31849 41599 31907 41605
rect 31849 41596 31861 41599
rect 31680 41568 31861 41596
rect 31849 41565 31861 41568
rect 31895 41565 31907 41599
rect 31956 41596 31984 41624
rect 32232 41605 32260 41636
rect 32766 41624 32772 41644
rect 32824 41624 32830 41676
rect 32968 41673 32996 41772
rect 33134 41760 33140 41812
rect 33192 41800 33198 41812
rect 33689 41803 33747 41809
rect 33689 41800 33701 41803
rect 33192 41772 33701 41800
rect 33192 41760 33198 41772
rect 33689 41769 33701 41772
rect 33735 41769 33747 41803
rect 33689 41763 33747 41769
rect 33778 41760 33784 41812
rect 33836 41800 33842 41812
rect 35621 41803 35679 41809
rect 35621 41800 35633 41803
rect 33836 41772 35633 41800
rect 33836 41760 33842 41772
rect 35621 41769 35633 41772
rect 35667 41769 35679 41803
rect 35621 41763 35679 41769
rect 33042 41692 33048 41744
rect 33100 41732 33106 41744
rect 34241 41735 34299 41741
rect 34241 41732 34253 41735
rect 33100 41704 34253 41732
rect 33100 41692 33106 41704
rect 34241 41701 34253 41704
rect 34287 41701 34299 41735
rect 34241 41695 34299 41701
rect 34698 41692 34704 41744
rect 34756 41692 34762 41744
rect 32953 41667 33011 41673
rect 32953 41633 32965 41667
rect 32999 41664 33011 41667
rect 34716 41664 34744 41692
rect 32999 41636 33824 41664
rect 32999 41633 33011 41636
rect 32953 41627 33011 41633
rect 33796 41608 33824 41636
rect 33888 41636 34744 41664
rect 32217 41599 32275 41605
rect 32217 41596 32229 41599
rect 31956 41568 32229 41596
rect 31849 41559 31907 41565
rect 32217 41565 32229 41568
rect 32263 41565 32275 41599
rect 32217 41559 32275 41565
rect 32401 41599 32459 41605
rect 32401 41565 32413 41599
rect 32447 41565 32459 41599
rect 32401 41559 32459 41565
rect 31386 41528 31392 41540
rect 31036 41500 31392 41528
rect 31386 41488 31392 41500
rect 31444 41488 31450 41540
rect 31665 41531 31723 41537
rect 31665 41497 31677 41531
rect 31711 41497 31723 41531
rect 32424 41528 32452 41559
rect 32490 41556 32496 41608
rect 32548 41556 32554 41608
rect 32674 41556 32680 41608
rect 32732 41556 32738 41608
rect 33045 41599 33103 41605
rect 33045 41565 33057 41599
rect 33091 41596 33103 41599
rect 33502 41596 33508 41608
rect 33091 41568 33508 41596
rect 33091 41565 33103 41568
rect 33045 41559 33103 41565
rect 33060 41528 33088 41559
rect 33502 41556 33508 41568
rect 33560 41556 33566 41608
rect 33778 41556 33784 41608
rect 33836 41556 33842 41608
rect 33888 41605 33916 41636
rect 33873 41599 33931 41605
rect 33873 41565 33885 41599
rect 33919 41565 33931 41599
rect 33873 41559 33931 41565
rect 34054 41556 34060 41608
rect 34112 41556 34118 41608
rect 34146 41556 34152 41608
rect 34204 41556 34210 41608
rect 34256 41605 34284 41636
rect 34790 41624 34796 41676
rect 34848 41664 34854 41676
rect 34848 41636 34928 41664
rect 34848 41624 34854 41636
rect 34241 41599 34299 41605
rect 34241 41565 34253 41599
rect 34287 41565 34299 41599
rect 34241 41559 34299 41565
rect 34425 41599 34483 41605
rect 34425 41565 34437 41599
rect 34471 41565 34483 41599
rect 34425 41559 34483 41565
rect 32424 41500 33088 41528
rect 31665 41491 31723 41497
rect 29748 41432 30098 41460
rect 30374 41420 30380 41472
rect 30432 41460 30438 41472
rect 31573 41463 31631 41469
rect 31573 41460 31585 41463
rect 30432 41432 31585 41460
rect 30432 41420 30438 41432
rect 31573 41429 31585 41432
rect 31619 41429 31631 41463
rect 31680 41460 31708 41491
rect 33410 41488 33416 41540
rect 33468 41488 33474 41540
rect 33594 41488 33600 41540
rect 33652 41488 33658 41540
rect 34164 41528 34192 41556
rect 34072 41500 34192 41528
rect 31846 41460 31852 41472
rect 31680 41432 31852 41460
rect 31573 41423 31631 41429
rect 31846 41420 31852 41432
rect 31904 41420 31910 41472
rect 31938 41420 31944 41472
rect 31996 41420 32002 41472
rect 33229 41463 33287 41469
rect 33229 41429 33241 41463
rect 33275 41460 33287 41463
rect 34072 41460 34100 41500
rect 34330 41488 34336 41540
rect 34388 41528 34394 41540
rect 34440 41528 34468 41559
rect 34698 41556 34704 41608
rect 34756 41556 34762 41608
rect 34900 41605 34928 41636
rect 34885 41599 34943 41605
rect 34885 41565 34897 41599
rect 34931 41565 34943 41599
rect 34885 41559 34943 41565
rect 35526 41537 35532 41540
rect 34793 41531 34851 41537
rect 34793 41528 34805 41531
rect 34388 41500 34805 41528
rect 34388 41488 34394 41500
rect 34793 41497 34805 41500
rect 34839 41497 34851 41531
rect 34793 41491 34851 41497
rect 35511 41531 35532 41537
rect 35511 41497 35523 41531
rect 35511 41491 35532 41497
rect 35526 41488 35532 41491
rect 35584 41488 35590 41540
rect 33275 41432 34100 41460
rect 33275 41429 33287 41432
rect 33229 41423 33287 41429
rect 1104 41370 45172 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 45172 41370
rect 1104 41296 45172 41318
rect 2774 41216 2780 41268
rect 2832 41256 2838 41268
rect 3053 41259 3111 41265
rect 3053 41256 3065 41259
rect 2832 41228 3065 41256
rect 2832 41216 2838 41228
rect 3053 41225 3065 41228
rect 3099 41225 3111 41259
rect 3053 41219 3111 41225
rect 4154 41216 4160 41268
rect 4212 41256 4218 41268
rect 4522 41256 4528 41268
rect 4212 41228 4528 41256
rect 4212 41216 4218 41228
rect 4522 41216 4528 41228
rect 4580 41216 4586 41268
rect 4982 41256 4988 41268
rect 4632 41228 4988 41256
rect 4632 41188 4660 41228
rect 4982 41216 4988 41228
rect 5040 41216 5046 41268
rect 9125 41259 9183 41265
rect 9125 41225 9137 41259
rect 9171 41256 9183 41259
rect 9306 41256 9312 41268
rect 9171 41228 9312 41256
rect 9171 41225 9183 41228
rect 9125 41219 9183 41225
rect 9306 41216 9312 41228
rect 9364 41216 9370 41268
rect 10502 41216 10508 41268
rect 10560 41216 10566 41268
rect 11882 41216 11888 41268
rect 11940 41216 11946 41268
rect 14182 41216 14188 41268
rect 14240 41256 14246 41268
rect 15197 41259 15255 41265
rect 14240 41228 14504 41256
rect 14240 41216 14246 41228
rect 3988 41160 4660 41188
rect 4893 41191 4951 41197
rect 3988 41129 4016 41160
rect 4893 41157 4905 41191
rect 4939 41188 4951 41191
rect 5166 41188 5172 41200
rect 4939 41160 5172 41188
rect 4939 41157 4951 41160
rect 4893 41151 4951 41157
rect 5166 41148 5172 41160
rect 5224 41148 5230 41200
rect 8018 41148 8024 41200
rect 8076 41188 8082 41200
rect 10410 41188 10416 41200
rect 8076 41160 10416 41188
rect 8076 41148 8082 41160
rect 10410 41148 10416 41160
rect 10468 41148 10474 41200
rect 11238 41148 11244 41200
rect 11296 41188 11302 41200
rect 14476 41197 14504 41228
rect 15197 41225 15209 41259
rect 15243 41256 15255 41259
rect 15243 41228 15608 41256
rect 15243 41225 15255 41228
rect 15197 41219 15255 41225
rect 14369 41191 14427 41197
rect 11296 41160 12204 41188
rect 11296 41148 11302 41160
rect 3968 41123 4026 41129
rect 3968 41089 3980 41123
rect 4014 41089 4026 41123
rect 3968 41083 4026 41089
rect 4065 41123 4123 41129
rect 4065 41089 4077 41123
rect 4111 41089 4123 41123
rect 4065 41083 4123 41089
rect 3697 41055 3755 41061
rect 3697 41021 3709 41055
rect 3743 41021 3755 41055
rect 3697 41015 3755 41021
rect 3712 40984 3740 41015
rect 3786 41012 3792 41064
rect 3844 41052 3850 41064
rect 4080 41052 4108 41083
rect 4154 41080 4160 41132
rect 4212 41080 4218 41132
rect 4338 41120 4344 41132
rect 4299 41092 4344 41120
rect 4338 41080 4344 41092
rect 4396 41080 4402 41132
rect 4433 41123 4491 41129
rect 4433 41089 4445 41123
rect 4479 41089 4491 41123
rect 4433 41083 4491 41089
rect 3844 41024 4108 41052
rect 4448 41052 4476 41083
rect 4522 41080 4528 41132
rect 4580 41080 4586 41132
rect 4706 41129 4712 41132
rect 4673 41123 4712 41129
rect 4673 41089 4685 41123
rect 4673 41083 4712 41089
rect 4706 41080 4712 41083
rect 4764 41080 4770 41132
rect 4798 41080 4804 41132
rect 4856 41080 4862 41132
rect 4982 41080 4988 41132
rect 5040 41129 5046 41132
rect 5040 41120 5048 41129
rect 5445 41123 5503 41129
rect 5040 41092 5085 41120
rect 5040 41083 5048 41092
rect 5445 41089 5457 41123
rect 5491 41089 5503 41123
rect 5445 41083 5503 41089
rect 5040 41080 5046 41083
rect 5261 41055 5319 41061
rect 5261 41052 5273 41055
rect 4448 41024 5273 41052
rect 3844 41012 3850 41024
rect 5261 41021 5273 41024
rect 5307 41021 5319 41055
rect 5261 41015 5319 41021
rect 5169 40987 5227 40993
rect 5169 40984 5181 40987
rect 3712 40956 5181 40984
rect 5169 40953 5181 40956
rect 5215 40953 5227 40987
rect 5169 40947 5227 40953
rect 5460 40928 5488 41083
rect 8846 41080 8852 41132
rect 8904 41120 8910 41132
rect 9677 41123 9735 41129
rect 9677 41120 9689 41123
rect 8904 41092 9689 41120
rect 8904 41080 8910 41092
rect 9677 41089 9689 41092
rect 9723 41089 9735 41123
rect 9677 41083 9735 41089
rect 10689 41123 10747 41129
rect 10689 41089 10701 41123
rect 10735 41120 10747 41123
rect 10735 41092 11560 41120
rect 10735 41089 10747 41092
rect 10689 41083 10747 41089
rect 5629 41055 5687 41061
rect 5629 41021 5641 41055
rect 5675 41052 5687 41055
rect 6086 41052 6092 41064
rect 5675 41024 6092 41052
rect 5675 41021 5687 41024
rect 5629 41015 5687 41021
rect 6086 41012 6092 41024
rect 6144 41012 6150 41064
rect 8110 41012 8116 41064
rect 8168 41012 8174 41064
rect 11532 40993 11560 41092
rect 12176 41064 12204 41160
rect 14369 41157 14381 41191
rect 14415 41157 14427 41191
rect 14369 41151 14427 41157
rect 14461 41191 14519 41197
rect 14461 41157 14473 41191
rect 14507 41157 14519 41191
rect 15286 41188 15292 41200
rect 14461 41151 14519 41157
rect 14660 41160 15292 41188
rect 14274 41129 14280 41132
rect 13449 41123 13507 41129
rect 13449 41089 13461 41123
rect 13495 41120 13507 41123
rect 14272 41120 14280 41129
rect 13495 41092 13676 41120
rect 14235 41092 14280 41120
rect 13495 41089 13507 41092
rect 13449 41083 13507 41089
rect 11974 41012 11980 41064
rect 12032 41012 12038 41064
rect 12158 41012 12164 41064
rect 12216 41052 12222 41064
rect 13173 41055 13231 41061
rect 13173 41052 13185 41055
rect 12216 41024 13185 41052
rect 12216 41012 12222 41024
rect 13173 41021 13185 41024
rect 13219 41021 13231 41055
rect 13173 41015 13231 41021
rect 11517 40987 11575 40993
rect 11517 40953 11529 40987
rect 11563 40953 11575 40987
rect 11517 40947 11575 40953
rect 13648 40928 13676 41092
rect 14272 41083 14280 41092
rect 14274 41080 14280 41083
rect 14332 41080 14338 41132
rect 14384 41120 14412 41151
rect 14550 41120 14556 41132
rect 14384 41092 14556 41120
rect 14550 41080 14556 41092
rect 14608 41080 14614 41132
rect 14660 41129 14688 41160
rect 15286 41148 15292 41160
rect 15344 41148 15350 41200
rect 15580 41188 15608 41228
rect 15746 41216 15752 41268
rect 15804 41216 15810 41268
rect 16022 41216 16028 41268
rect 16080 41216 16086 41268
rect 18782 41216 18788 41268
rect 18840 41216 18846 41268
rect 21174 41216 21180 41268
rect 21232 41216 21238 41268
rect 21450 41216 21456 41268
rect 21508 41256 21514 41268
rect 21545 41259 21603 41265
rect 21545 41256 21557 41259
rect 21508 41228 21557 41256
rect 21508 41216 21514 41228
rect 21545 41225 21557 41228
rect 21591 41225 21603 41259
rect 21545 41219 21603 41225
rect 23474 41216 23480 41268
rect 23532 41256 23538 41268
rect 23569 41259 23627 41265
rect 23569 41256 23581 41259
rect 23532 41228 23581 41256
rect 23532 41216 23538 41228
rect 23569 41225 23581 41228
rect 23615 41225 23627 41259
rect 25314 41256 25320 41268
rect 23569 41219 23627 41225
rect 24136 41228 25320 41256
rect 16040 41188 16068 41216
rect 15580 41160 16068 41188
rect 17310 41148 17316 41200
rect 17368 41188 17374 41200
rect 18322 41188 18328 41200
rect 17368 41160 18328 41188
rect 17368 41148 17374 41160
rect 18322 41148 18328 41160
rect 18380 41188 18386 41200
rect 18380 41160 20300 41188
rect 18380 41148 18386 41160
rect 14644 41123 14702 41129
rect 14644 41089 14656 41123
rect 14690 41089 14702 41123
rect 14644 41083 14702 41089
rect 14734 41080 14740 41132
rect 14792 41080 14798 41132
rect 15013 41123 15071 41129
rect 15013 41089 15025 41123
rect 15059 41120 15071 41123
rect 15059 41092 15424 41120
rect 15059 41089 15071 41092
rect 15013 41083 15071 41089
rect 14093 40987 14151 40993
rect 14093 40953 14105 40987
rect 14139 40984 14151 40987
rect 14642 40984 14648 40996
rect 14139 40956 14648 40984
rect 14139 40953 14151 40956
rect 14093 40947 14151 40953
rect 14642 40944 14648 40956
rect 14700 40944 14706 40996
rect 15396 40993 15424 41092
rect 15838 41012 15844 41064
rect 15896 41012 15902 41064
rect 16025 41055 16083 41061
rect 16025 41021 16037 41055
rect 16071 41052 16083 41055
rect 17328 41052 17356 41148
rect 18690 41080 18696 41132
rect 18748 41080 18754 41132
rect 20272 41129 20300 41160
rect 20438 41148 20444 41200
rect 20496 41188 20502 41200
rect 20533 41191 20591 41197
rect 20533 41188 20545 41191
rect 20496 41160 20545 41188
rect 20496 41148 20502 41160
rect 20533 41157 20545 41160
rect 20579 41157 20591 41191
rect 21192 41188 21220 41216
rect 22186 41188 22192 41200
rect 21192 41160 21496 41188
rect 20533 41151 20591 41157
rect 21468 41129 21496 41160
rect 21652 41160 22192 41188
rect 21652 41129 21680 41160
rect 22186 41148 22192 41160
rect 22244 41148 22250 41200
rect 23290 41188 23296 41200
rect 23032 41160 23296 41188
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41120 20315 41123
rect 21177 41123 21235 41129
rect 20303 41092 20576 41120
rect 20303 41089 20315 41092
rect 20257 41083 20315 41089
rect 16071 41024 17356 41052
rect 16071 41021 16083 41024
rect 16025 41015 16083 41021
rect 15381 40987 15439 40993
rect 15381 40953 15393 40987
rect 15427 40953 15439 40987
rect 15381 40947 15439 40953
rect 3510 40876 3516 40928
rect 3568 40916 3574 40928
rect 3789 40919 3847 40925
rect 3789 40916 3801 40919
rect 3568 40888 3801 40916
rect 3568 40876 3574 40888
rect 3789 40885 3801 40888
rect 3835 40885 3847 40919
rect 3789 40879 3847 40885
rect 4246 40876 4252 40928
rect 4304 40916 4310 40928
rect 5442 40916 5448 40928
rect 4304 40888 5448 40916
rect 4304 40876 4310 40888
rect 5442 40876 5448 40888
rect 5500 40876 5506 40928
rect 7466 40876 7472 40928
rect 7524 40876 7530 40928
rect 13630 40876 13636 40928
rect 13688 40916 13694 40928
rect 16040 40916 16068 41015
rect 20548 40928 20576 41092
rect 21177 41089 21189 41123
rect 21223 41089 21235 41123
rect 21177 41083 21235 41089
rect 21453 41123 21511 41129
rect 21453 41089 21465 41123
rect 21499 41089 21511 41123
rect 21453 41083 21511 41089
rect 21637 41123 21695 41129
rect 21637 41089 21649 41123
rect 21683 41089 21695 41123
rect 21637 41083 21695 41089
rect 22005 41123 22063 41129
rect 22005 41089 22017 41123
rect 22051 41120 22063 41123
rect 22373 41123 22431 41129
rect 22373 41120 22385 41123
rect 22051 41092 22385 41120
rect 22051 41089 22063 41092
rect 22005 41083 22063 41089
rect 22373 41089 22385 41092
rect 22419 41120 22431 41123
rect 22419 41092 22784 41120
rect 22419 41089 22431 41092
rect 22373 41083 22431 41089
rect 21192 41052 21220 41083
rect 21821 41055 21879 41061
rect 21821 41052 21833 41055
rect 21192 41024 21833 41052
rect 21821 41021 21833 41024
rect 21867 41021 21879 41055
rect 21821 41015 21879 41021
rect 22189 41055 22247 41061
rect 22189 41021 22201 41055
rect 22235 41052 22247 41055
rect 22554 41052 22560 41064
rect 22235 41024 22560 41052
rect 22235 41021 22247 41024
rect 22189 41015 22247 41021
rect 22554 41012 22560 41024
rect 22612 41012 22618 41064
rect 22756 41052 22784 41092
rect 22830 41080 22836 41132
rect 22888 41080 22894 41132
rect 23032 41129 23060 41160
rect 23290 41148 23296 41160
rect 23348 41148 23354 41200
rect 24136 41197 24164 41228
rect 25314 41216 25320 41228
rect 25372 41216 25378 41268
rect 28077 41259 28135 41265
rect 28077 41225 28089 41259
rect 28123 41256 28135 41259
rect 28258 41256 28264 41268
rect 28123 41228 28264 41256
rect 28123 41225 28135 41228
rect 28077 41219 28135 41225
rect 28258 41216 28264 41228
rect 28316 41216 28322 41268
rect 30193 41259 30251 41265
rect 30193 41225 30205 41259
rect 30239 41256 30251 41259
rect 30282 41256 30288 41268
rect 30239 41228 30288 41256
rect 30239 41225 30251 41228
rect 30193 41219 30251 41225
rect 30282 41216 30288 41228
rect 30340 41216 30346 41268
rect 30469 41259 30527 41265
rect 30469 41225 30481 41259
rect 30515 41225 30527 41259
rect 30469 41219 30527 41225
rect 30561 41259 30619 41265
rect 30561 41225 30573 41259
rect 30607 41256 30619 41259
rect 30834 41256 30840 41268
rect 30607 41228 30840 41256
rect 30607 41225 30619 41228
rect 30561 41219 30619 41225
rect 24121 41191 24179 41197
rect 24121 41157 24133 41191
rect 24167 41157 24179 41191
rect 24121 41151 24179 41157
rect 25222 41148 25228 41200
rect 25280 41148 25286 41200
rect 26786 41148 26792 41200
rect 26844 41188 26850 41200
rect 28629 41191 28687 41197
rect 26844 41160 28120 41188
rect 26844 41148 26850 41160
rect 23017 41123 23075 41129
rect 23017 41089 23029 41123
rect 23063 41089 23075 41123
rect 23017 41083 23075 41089
rect 23198 41080 23204 41132
rect 23256 41080 23262 41132
rect 23385 41123 23443 41129
rect 23385 41089 23397 41123
rect 23431 41120 23443 41123
rect 23474 41120 23480 41132
rect 23431 41092 23480 41120
rect 23431 41089 23443 41092
rect 23385 41083 23443 41089
rect 23474 41080 23480 41092
rect 23532 41080 23538 41132
rect 23746 41123 23804 41129
rect 23746 41120 23758 41123
rect 23676 41092 23758 41120
rect 23216 41052 23244 41080
rect 23676 41064 23704 41092
rect 23746 41089 23758 41092
rect 23792 41089 23804 41123
rect 23746 41083 23804 41089
rect 23845 41123 23903 41129
rect 23845 41089 23857 41123
rect 23891 41089 23903 41123
rect 23845 41083 23903 41089
rect 22756 41024 23244 41052
rect 23216 40984 23244 41024
rect 23293 41055 23351 41061
rect 23293 41021 23305 41055
rect 23339 41052 23351 41055
rect 23658 41052 23664 41064
rect 23339 41024 23664 41052
rect 23339 41021 23351 41024
rect 23293 41015 23351 41021
rect 23658 41012 23664 41024
rect 23716 41012 23722 41064
rect 23860 40984 23888 41083
rect 26326 41080 26332 41132
rect 26384 41120 26390 41132
rect 27246 41120 27252 41132
rect 26384 41092 27252 41120
rect 26384 41080 26390 41092
rect 27246 41080 27252 41092
rect 27304 41080 27310 41132
rect 28092 41130 28120 41160
rect 28399 41157 28457 41163
rect 28092 41129 28212 41130
rect 27893 41123 27951 41129
rect 27893 41120 27905 41123
rect 27540 41092 27905 41120
rect 24394 41012 24400 41064
rect 24452 41012 24458 41064
rect 24670 41012 24676 41064
rect 24728 41012 24734 41064
rect 27540 41061 27568 41092
rect 27893 41089 27905 41092
rect 27939 41089 27951 41123
rect 28092 41123 28227 41129
rect 28092 41102 28181 41123
rect 27893 41083 27951 41089
rect 28169 41089 28181 41102
rect 28215 41118 28227 41123
rect 28399 41123 28411 41157
rect 28445 41123 28457 41157
rect 28629 41157 28641 41191
rect 28675 41157 28687 41191
rect 28629 41151 28687 41157
rect 28399 41120 28457 41123
rect 28276 41118 28457 41120
rect 28215 41117 28457 41118
rect 28215 41092 28456 41117
rect 28215 41090 28304 41092
rect 28215 41089 28227 41090
rect 28169 41083 28227 41089
rect 26145 41055 26203 41061
rect 26145 41021 26157 41055
rect 26191 41052 26203 41055
rect 27525 41055 27583 41061
rect 27525 41052 27537 41055
rect 26191 41024 27537 41052
rect 26191 41021 26203 41024
rect 26145 41015 26203 41021
rect 27525 41021 27537 41024
rect 27571 41021 27583 41055
rect 27525 41015 27583 41021
rect 23216 40956 23888 40984
rect 27908 40984 27936 41083
rect 28644 41052 28672 41151
rect 28810 41148 28816 41200
rect 28868 41148 28874 41200
rect 30484 41188 30512 41219
rect 30834 41216 30840 41228
rect 30892 41216 30898 41268
rect 31662 41216 31668 41268
rect 31720 41256 31726 41268
rect 31720 41228 32260 41256
rect 31720 41216 31726 41228
rect 30484 41160 30880 41188
rect 30193 41123 30251 41129
rect 30193 41120 30205 41123
rect 28460 41024 28672 41052
rect 28736 41092 30205 41120
rect 28460 40984 28488 41024
rect 28736 40984 28764 41092
rect 30193 41089 30205 41092
rect 30239 41089 30251 41123
rect 30193 41083 30251 41089
rect 30653 41123 30711 41129
rect 30653 41089 30665 41123
rect 30699 41089 30711 41123
rect 30653 41083 30711 41089
rect 30745 41123 30803 41129
rect 30745 41089 30757 41123
rect 30791 41089 30803 41123
rect 30852 41120 30880 41160
rect 30926 41148 30932 41200
rect 30984 41148 30990 41200
rect 31570 41148 31576 41200
rect 31628 41148 31634 41200
rect 31202 41120 31208 41132
rect 30852 41092 31208 41120
rect 30745 41083 30803 41089
rect 29089 41055 29147 41061
rect 29089 41021 29101 41055
rect 29135 41052 29147 41055
rect 30558 41052 30564 41064
rect 29135 41024 30564 41052
rect 29135 41021 29147 41024
rect 29089 41015 29147 41021
rect 30558 41012 30564 41024
rect 30616 41012 30622 41064
rect 27908 40956 28488 40984
rect 28552 40956 28764 40984
rect 30668 40984 30696 41083
rect 30760 41052 30788 41083
rect 31202 41080 31208 41092
rect 31260 41080 31266 41132
rect 31481 41123 31539 41129
rect 31481 41089 31493 41123
rect 31527 41120 31539 41123
rect 31588 41120 31616 41148
rect 31527 41092 31616 41120
rect 31665 41123 31723 41129
rect 31527 41089 31539 41092
rect 31481 41083 31539 41089
rect 31665 41089 31677 41123
rect 31711 41120 31723 41123
rect 31846 41120 31852 41132
rect 31711 41092 31852 41120
rect 31711 41089 31723 41092
rect 31665 41083 31723 41089
rect 31846 41080 31852 41092
rect 31904 41080 31910 41132
rect 32122 41080 32128 41132
rect 32180 41080 32186 41132
rect 32232 41120 32260 41228
rect 33686 41216 33692 41268
rect 33744 41256 33750 41268
rect 34149 41259 34207 41265
rect 34149 41256 34161 41259
rect 33744 41228 34161 41256
rect 33744 41216 33750 41228
rect 34149 41225 34161 41228
rect 34195 41225 34207 41259
rect 34149 41219 34207 41225
rect 34238 41216 34244 41268
rect 34296 41256 34302 41268
rect 34517 41259 34575 41265
rect 34517 41256 34529 41259
rect 34296 41228 34529 41256
rect 34296 41216 34302 41228
rect 34517 41225 34529 41228
rect 34563 41256 34575 41259
rect 34790 41256 34796 41268
rect 34563 41228 34796 41256
rect 34563 41225 34575 41228
rect 34517 41219 34575 41225
rect 34790 41216 34796 41228
rect 34848 41216 34854 41268
rect 35066 41216 35072 41268
rect 35124 41256 35130 41268
rect 35526 41256 35532 41268
rect 35124 41228 35532 41256
rect 35124 41216 35130 41228
rect 35526 41216 35532 41228
rect 35584 41256 35590 41268
rect 35584 41228 35664 41256
rect 35584 41216 35590 41228
rect 32490 41148 32496 41200
rect 32548 41188 32554 41200
rect 33042 41188 33048 41200
rect 32548 41160 33048 41188
rect 32548 41148 32554 41160
rect 32300 41123 32358 41129
rect 32300 41120 32312 41123
rect 32232 41092 32312 41120
rect 32300 41089 32312 41092
rect 32346 41089 32358 41123
rect 32300 41083 32358 41089
rect 32398 41080 32404 41132
rect 32456 41080 32462 41132
rect 32600 41129 32628 41160
rect 33042 41148 33048 41160
rect 33100 41148 33106 41200
rect 34057 41191 34115 41197
rect 33612 41160 34008 41188
rect 33612 41132 33640 41160
rect 32585 41123 32643 41129
rect 32585 41089 32597 41123
rect 32631 41089 32643 41123
rect 32585 41083 32643 41089
rect 33594 41080 33600 41132
rect 33652 41080 33658 41132
rect 33689 41123 33747 41129
rect 33689 41089 33701 41123
rect 33735 41089 33747 41123
rect 33689 41083 33747 41089
rect 30926 41052 30932 41064
rect 30760 41024 30932 41052
rect 30926 41012 30932 41024
rect 30984 41012 30990 41064
rect 31110 41012 31116 41064
rect 31168 41012 31174 41064
rect 31389 41055 31447 41061
rect 31389 41021 31401 41055
rect 31435 41021 31447 41055
rect 31389 41015 31447 41021
rect 31404 40984 31432 41015
rect 31570 41012 31576 41064
rect 31628 41012 31634 41064
rect 31938 41012 31944 41064
rect 31996 41052 32002 41064
rect 32217 41055 32275 41061
rect 32217 41052 32229 41055
rect 31996 41024 32229 41052
rect 31996 41012 32002 41024
rect 32217 41021 32229 41024
rect 32263 41021 32275 41055
rect 32217 41015 32275 41021
rect 31754 40984 31760 40996
rect 30668 40956 31340 40984
rect 31404 40956 31760 40984
rect 28552 40928 28580 40956
rect 13688 40888 16068 40916
rect 13688 40876 13694 40888
rect 20530 40876 20536 40928
rect 20588 40916 20594 40928
rect 20901 40919 20959 40925
rect 20901 40916 20913 40919
rect 20588 40888 20913 40916
rect 20588 40876 20594 40888
rect 20901 40885 20913 40888
rect 20947 40885 20959 40919
rect 20901 40879 20959 40885
rect 22646 40876 22652 40928
rect 22704 40876 22710 40928
rect 22925 40919 22983 40925
rect 22925 40885 22937 40919
rect 22971 40916 22983 40919
rect 24486 40916 24492 40928
rect 22971 40888 24492 40916
rect 22971 40885 22983 40888
rect 22925 40879 22983 40885
rect 24486 40876 24492 40888
rect 24544 40876 24550 40928
rect 26510 40876 26516 40928
rect 26568 40916 26574 40928
rect 26973 40919 27031 40925
rect 26973 40916 26985 40919
rect 26568 40888 26985 40916
rect 26568 40876 26574 40888
rect 26973 40885 26985 40888
rect 27019 40885 27031 40919
rect 26973 40879 27031 40885
rect 27154 40876 27160 40928
rect 27212 40916 27218 40928
rect 27709 40919 27767 40925
rect 27709 40916 27721 40919
rect 27212 40888 27721 40916
rect 27212 40876 27218 40888
rect 27709 40885 27721 40888
rect 27755 40885 27767 40919
rect 27709 40879 27767 40885
rect 28258 40876 28264 40928
rect 28316 40876 28322 40928
rect 28350 40876 28356 40928
rect 28408 40916 28414 40928
rect 28445 40919 28503 40925
rect 28445 40916 28457 40919
rect 28408 40888 28457 40916
rect 28408 40876 28414 40888
rect 28445 40885 28457 40888
rect 28491 40885 28503 40919
rect 28445 40879 28503 40885
rect 28534 40876 28540 40928
rect 28592 40876 28598 40928
rect 30282 40876 30288 40928
rect 30340 40876 30346 40928
rect 31202 40876 31208 40928
rect 31260 40876 31266 40928
rect 31312 40916 31340 40956
rect 31754 40944 31760 40956
rect 31812 40944 31818 40996
rect 32140 40956 32536 40984
rect 31386 40916 31392 40928
rect 31312 40888 31392 40916
rect 31386 40876 31392 40888
rect 31444 40916 31450 40928
rect 32140 40916 32168 40956
rect 32508 40925 32536 40956
rect 31444 40888 32168 40916
rect 32493 40919 32551 40925
rect 31444 40876 31450 40888
rect 32493 40885 32505 40919
rect 32539 40885 32551 40919
rect 33704 40916 33732 41083
rect 33778 41080 33784 41132
rect 33836 41120 33842 41132
rect 33873 41123 33931 41129
rect 33873 41120 33885 41123
rect 33836 41092 33885 41120
rect 33836 41080 33842 41092
rect 33873 41089 33885 41092
rect 33919 41089 33931 41123
rect 33980 41120 34008 41160
rect 34057 41157 34069 41191
rect 34103 41188 34115 41191
rect 34698 41188 34704 41200
rect 34103 41160 34704 41188
rect 34103 41157 34115 41160
rect 34057 41151 34115 41157
rect 34698 41148 34704 41160
rect 34756 41148 34762 41200
rect 35636 41197 35664 41228
rect 35621 41191 35679 41197
rect 35621 41157 35633 41191
rect 35667 41157 35679 41191
rect 35621 41151 35679 41157
rect 34149 41123 34207 41129
rect 34149 41120 34161 41123
rect 33980 41092 34161 41120
rect 33873 41083 33931 41089
rect 34149 41089 34161 41092
rect 34195 41089 34207 41123
rect 34149 41083 34207 41089
rect 33888 40984 33916 41083
rect 34330 41080 34336 41132
rect 34388 41080 34394 41132
rect 34425 41123 34483 41129
rect 34425 41089 34437 41123
rect 34471 41089 34483 41123
rect 34425 41083 34483 41089
rect 34440 41052 34468 41083
rect 34514 41080 34520 41132
rect 34572 41120 34578 41132
rect 34609 41123 34667 41129
rect 34609 41120 34621 41123
rect 34572 41092 34621 41120
rect 34572 41080 34578 41092
rect 34609 41089 34621 41092
rect 34655 41089 34667 41123
rect 34609 41083 34667 41089
rect 34440 41024 35940 41052
rect 34440 40984 34468 41024
rect 33888 40956 34468 40984
rect 35912 40928 35940 41024
rect 34422 40916 34428 40928
rect 33704 40888 34428 40916
rect 32493 40879 32551 40885
rect 34422 40876 34428 40888
rect 34480 40876 34486 40928
rect 35529 40919 35587 40925
rect 35529 40885 35541 40919
rect 35575 40916 35587 40919
rect 35802 40916 35808 40928
rect 35575 40888 35808 40916
rect 35575 40885 35587 40888
rect 35529 40879 35587 40885
rect 35802 40876 35808 40888
rect 35860 40876 35866 40928
rect 35894 40876 35900 40928
rect 35952 40876 35958 40928
rect 1104 40826 45172 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 45172 40826
rect 1104 40752 45172 40774
rect 4614 40672 4620 40724
rect 4672 40712 4678 40724
rect 4801 40715 4859 40721
rect 4801 40712 4813 40715
rect 4672 40684 4813 40712
rect 4672 40672 4678 40684
rect 4801 40681 4813 40684
rect 4847 40681 4859 40715
rect 4801 40675 4859 40681
rect 6365 40715 6423 40721
rect 6365 40681 6377 40715
rect 6411 40712 6423 40715
rect 6730 40712 6736 40724
rect 6411 40684 6736 40712
rect 6411 40681 6423 40684
rect 6365 40675 6423 40681
rect 6730 40672 6736 40684
rect 6788 40672 6794 40724
rect 8754 40672 8760 40724
rect 8812 40712 8818 40724
rect 11790 40712 11796 40724
rect 8812 40684 11796 40712
rect 8812 40672 8818 40684
rect 11790 40672 11796 40684
rect 11848 40712 11854 40724
rect 16114 40712 16120 40724
rect 11848 40684 16120 40712
rect 11848 40672 11854 40684
rect 16114 40672 16120 40684
rect 16172 40712 16178 40724
rect 17862 40712 17868 40724
rect 16172 40684 17868 40712
rect 16172 40672 16178 40684
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 18690 40672 18696 40724
rect 18748 40712 18754 40724
rect 22646 40712 22652 40724
rect 18748 40684 22652 40712
rect 18748 40672 18754 40684
rect 22646 40672 22652 40684
rect 22704 40672 22710 40724
rect 24670 40672 24676 40724
rect 24728 40712 24734 40724
rect 25869 40715 25927 40721
rect 25869 40712 25881 40715
rect 24728 40684 25881 40712
rect 24728 40672 24734 40684
rect 25869 40681 25881 40684
rect 25915 40681 25927 40715
rect 28534 40712 28540 40724
rect 25869 40675 25927 40681
rect 26160 40684 28540 40712
rect 3329 40647 3387 40653
rect 3329 40613 3341 40647
rect 3375 40644 3387 40647
rect 12161 40647 12219 40653
rect 3375 40616 5396 40644
rect 3375 40613 3387 40616
rect 3329 40607 3387 40613
rect 1581 40579 1639 40585
rect 1581 40545 1593 40579
rect 1627 40576 1639 40579
rect 1854 40576 1860 40588
rect 1627 40548 1860 40576
rect 1627 40545 1639 40548
rect 1581 40539 1639 40545
rect 1854 40536 1860 40548
rect 1912 40576 1918 40588
rect 3602 40576 3608 40588
rect 1912 40548 3608 40576
rect 1912 40536 1918 40548
rect 3602 40536 3608 40548
rect 3660 40536 3666 40588
rect 4154 40536 4160 40588
rect 4212 40576 4218 40588
rect 4798 40576 4804 40588
rect 4212 40548 4804 40576
rect 4212 40536 4218 40548
rect 4798 40536 4804 40548
rect 4856 40536 4862 40588
rect 5368 40585 5396 40616
rect 12161 40613 12173 40647
rect 12207 40644 12219 40647
rect 12207 40616 12848 40644
rect 12207 40613 12219 40616
rect 12161 40607 12219 40613
rect 5353 40579 5411 40585
rect 5353 40545 5365 40579
rect 5399 40545 5411 40579
rect 5353 40539 5411 40545
rect 6178 40536 6184 40588
rect 6236 40576 6242 40588
rect 6457 40579 6515 40585
rect 6457 40576 6469 40579
rect 6236 40548 6469 40576
rect 6236 40536 6242 40548
rect 6457 40545 6469 40548
rect 6503 40545 6515 40579
rect 6457 40539 6515 40545
rect 6733 40579 6791 40585
rect 6733 40545 6745 40579
rect 6779 40576 6791 40579
rect 7466 40576 7472 40588
rect 6779 40548 7472 40576
rect 6779 40545 6791 40548
rect 6733 40539 6791 40545
rect 7466 40536 7472 40548
rect 7524 40536 7530 40588
rect 8205 40579 8263 40585
rect 8205 40545 8217 40579
rect 8251 40576 8263 40579
rect 8662 40576 8668 40588
rect 8251 40548 8668 40576
rect 8251 40545 8263 40548
rect 8205 40539 8263 40545
rect 8662 40536 8668 40548
rect 8720 40536 8726 40588
rect 12820 40585 12848 40616
rect 25314 40604 25320 40656
rect 25372 40644 25378 40656
rect 26160 40644 26188 40684
rect 28534 40672 28540 40684
rect 28592 40672 28598 40724
rect 31294 40672 31300 40724
rect 31352 40712 31358 40724
rect 31938 40712 31944 40724
rect 31352 40684 31944 40712
rect 31352 40672 31358 40684
rect 31938 40672 31944 40684
rect 31996 40672 32002 40724
rect 26878 40644 26884 40656
rect 25372 40616 26188 40644
rect 26252 40616 26884 40644
rect 25372 40604 25378 40616
rect 10965 40579 11023 40585
rect 10965 40545 10977 40579
rect 11011 40576 11023 40579
rect 12805 40579 12863 40585
rect 11011 40548 12756 40576
rect 11011 40545 11023 40548
rect 10965 40539 11023 40545
rect 4614 40468 4620 40520
rect 4672 40468 4678 40520
rect 5074 40468 5080 40520
rect 5132 40508 5138 40520
rect 5721 40511 5779 40517
rect 5721 40508 5733 40511
rect 5132 40480 5733 40508
rect 5132 40468 5138 40480
rect 5721 40477 5733 40480
rect 5767 40477 5779 40511
rect 8018 40508 8024 40520
rect 7866 40480 8024 40508
rect 5721 40471 5779 40477
rect 8018 40468 8024 40480
rect 8076 40468 8082 40520
rect 8481 40511 8539 40517
rect 8481 40477 8493 40511
rect 8527 40477 8539 40511
rect 8481 40471 8539 40477
rect 1854 40400 1860 40452
rect 1912 40400 1918 40452
rect 3326 40440 3332 40452
rect 3082 40412 3332 40440
rect 3326 40400 3332 40412
rect 3384 40440 3390 40452
rect 4338 40440 4344 40452
rect 3384 40412 4344 40440
rect 3384 40400 3390 40412
rect 4338 40400 4344 40412
rect 4396 40400 4402 40452
rect 8496 40440 8524 40471
rect 8570 40468 8576 40520
rect 8628 40508 8634 40520
rect 9493 40511 9551 40517
rect 9493 40508 9505 40511
rect 8628 40480 9505 40508
rect 8628 40468 8634 40480
rect 9493 40477 9505 40480
rect 9539 40477 9551 40511
rect 9493 40471 9551 40477
rect 9876 40502 11008 40508
rect 11146 40502 11152 40520
rect 9876 40480 11152 40502
rect 9876 40440 9904 40480
rect 10980 40474 11152 40480
rect 11146 40468 11152 40474
rect 11204 40468 11210 40520
rect 11333 40511 11391 40517
rect 11333 40477 11345 40511
rect 11379 40508 11391 40511
rect 11517 40511 11575 40517
rect 11517 40508 11529 40511
rect 11379 40480 11529 40508
rect 11379 40477 11391 40480
rect 11333 40471 11391 40477
rect 11517 40477 11529 40480
rect 11563 40477 11575 40511
rect 11517 40471 11575 40477
rect 11610 40511 11668 40517
rect 11610 40477 11622 40511
rect 11656 40477 11668 40511
rect 11610 40471 11668 40477
rect 11982 40511 12040 40517
rect 11982 40477 11994 40511
rect 12028 40477 12040 40511
rect 12728 40508 12756 40548
rect 12805 40545 12817 40579
rect 12851 40545 12863 40579
rect 15930 40576 15936 40588
rect 12805 40539 12863 40545
rect 13648 40548 15936 40576
rect 13648 40508 13676 40548
rect 15930 40536 15936 40548
rect 15988 40576 15994 40588
rect 16485 40579 16543 40585
rect 16485 40576 16497 40579
rect 15988 40548 16497 40576
rect 15988 40536 15994 40548
rect 16485 40545 16497 40548
rect 16531 40545 16543 40579
rect 17494 40576 17500 40588
rect 16485 40539 16543 40545
rect 16868 40548 17500 40576
rect 12728 40480 13676 40508
rect 11982 40471 12040 40477
rect 8220 40412 9904 40440
rect 8220 40384 8248 40412
rect 10042 40400 10048 40452
rect 10100 40440 10106 40452
rect 11624 40440 11652 40471
rect 10100 40412 11652 40440
rect 10100 40400 10106 40412
rect 11790 40400 11796 40452
rect 11848 40400 11854 40452
rect 11882 40400 11888 40452
rect 11940 40400 11946 40452
rect 11997 40440 12025 40471
rect 13722 40468 13728 40520
rect 13780 40468 13786 40520
rect 14458 40468 14464 40520
rect 14516 40508 14522 40520
rect 16868 40508 16896 40548
rect 17494 40536 17500 40548
rect 17552 40536 17558 40588
rect 18233 40579 18291 40585
rect 18233 40545 18245 40579
rect 18279 40576 18291 40579
rect 19150 40576 19156 40588
rect 18279 40548 19156 40576
rect 18279 40545 18291 40548
rect 18233 40539 18291 40545
rect 19150 40536 19156 40548
rect 19208 40536 19214 40588
rect 14516 40494 16896 40508
rect 18877 40511 18935 40517
rect 14516 40480 16882 40494
rect 14516 40468 14522 40480
rect 18877 40477 18889 40511
rect 18923 40477 18935 40511
rect 18877 40471 18935 40477
rect 17957 40443 18015 40449
rect 11997 40412 16068 40440
rect 4062 40332 4068 40384
rect 4120 40332 4126 40384
rect 8202 40332 8208 40384
rect 8260 40332 8266 40384
rect 8294 40332 8300 40384
rect 8352 40332 8358 40384
rect 8386 40332 8392 40384
rect 8444 40372 8450 40384
rect 8941 40375 8999 40381
rect 8941 40372 8953 40375
rect 8444 40344 8953 40372
rect 8444 40332 8450 40344
rect 8941 40341 8953 40344
rect 8987 40341 8999 40375
rect 8941 40335 8999 40341
rect 9214 40332 9220 40384
rect 9272 40372 9278 40384
rect 11997 40372 12025 40412
rect 16040 40384 16068 40412
rect 17957 40409 17969 40443
rect 18003 40440 18015 40443
rect 18325 40443 18383 40449
rect 18325 40440 18337 40443
rect 18003 40412 18337 40440
rect 18003 40409 18015 40412
rect 17957 40403 18015 40409
rect 18325 40409 18337 40412
rect 18371 40409 18383 40443
rect 18325 40403 18383 40409
rect 9272 40344 12025 40372
rect 9272 40332 9278 40344
rect 12250 40332 12256 40384
rect 12308 40332 12314 40384
rect 13906 40332 13912 40384
rect 13964 40332 13970 40384
rect 16022 40332 16028 40384
rect 16080 40332 16086 40384
rect 17678 40332 17684 40384
rect 17736 40372 17742 40384
rect 18892 40372 18920 40471
rect 20162 40468 20168 40520
rect 20220 40468 20226 40520
rect 23658 40468 23664 40520
rect 23716 40508 23722 40520
rect 23845 40511 23903 40517
rect 23845 40508 23857 40511
rect 23716 40480 23857 40508
rect 23716 40468 23722 40480
rect 23845 40477 23857 40480
rect 23891 40477 23903 40511
rect 23845 40471 23903 40477
rect 26053 40511 26111 40517
rect 26053 40477 26065 40511
rect 26099 40477 26111 40511
rect 26053 40471 26111 40477
rect 17736 40344 18920 40372
rect 20809 40375 20867 40381
rect 17736 40332 17742 40344
rect 20809 40341 20821 40375
rect 20855 40372 20867 40375
rect 20898 40372 20904 40384
rect 20855 40344 20904 40372
rect 20855 40341 20867 40344
rect 20809 40335 20867 40341
rect 20898 40332 20904 40344
rect 20956 40332 20962 40384
rect 24029 40375 24087 40381
rect 24029 40341 24041 40375
rect 24075 40372 24087 40375
rect 24118 40372 24124 40384
rect 24075 40344 24124 40372
rect 24075 40341 24087 40344
rect 24029 40335 24087 40341
rect 24118 40332 24124 40344
rect 24176 40332 24182 40384
rect 26068 40372 26096 40471
rect 26142 40468 26148 40520
rect 26200 40468 26206 40520
rect 26252 40517 26280 40616
rect 26878 40604 26884 40616
rect 26936 40604 26942 40656
rect 35805 40647 35863 40653
rect 35805 40613 35817 40647
rect 35851 40613 35863 40647
rect 35805 40607 35863 40613
rect 26510 40536 26516 40588
rect 26568 40536 26574 40588
rect 27798 40576 27804 40588
rect 27172 40548 27804 40576
rect 26237 40511 26295 40517
rect 26237 40477 26249 40511
rect 26283 40477 26295 40511
rect 26237 40471 26295 40477
rect 26881 40511 26939 40517
rect 26881 40477 26893 40511
rect 26927 40508 26939 40511
rect 27172 40508 27200 40548
rect 27798 40536 27804 40548
rect 27856 40536 27862 40588
rect 31570 40536 31576 40588
rect 31628 40576 31634 40588
rect 32398 40576 32404 40588
rect 31628 40548 32404 40576
rect 31628 40536 31634 40548
rect 32398 40536 32404 40548
rect 32456 40536 32462 40588
rect 35820 40576 35848 40607
rect 37369 40579 37427 40585
rect 37369 40576 37381 40579
rect 35820 40548 37381 40576
rect 37369 40545 37381 40548
rect 37415 40545 37427 40579
rect 37369 40539 37427 40545
rect 26927 40480 27200 40508
rect 27249 40511 27307 40517
rect 26927 40477 26939 40480
rect 26881 40471 26939 40477
rect 27249 40477 27261 40511
rect 27295 40508 27307 40511
rect 27338 40508 27344 40520
rect 27295 40480 27344 40508
rect 27295 40477 27307 40480
rect 27249 40471 27307 40477
rect 27338 40468 27344 40480
rect 27396 40468 27402 40520
rect 27525 40511 27583 40517
rect 27525 40477 27537 40511
rect 27571 40508 27583 40511
rect 28258 40508 28264 40520
rect 27571 40480 28264 40508
rect 27571 40477 27583 40480
rect 27525 40471 27583 40477
rect 28258 40468 28264 40480
rect 28316 40468 28322 40520
rect 35250 40468 35256 40520
rect 35308 40468 35314 40520
rect 35621 40511 35679 40517
rect 35621 40508 35633 40511
rect 35360 40480 35633 40508
rect 26326 40400 26332 40452
rect 26384 40449 26390 40452
rect 26384 40443 26413 40449
rect 26401 40409 26413 40443
rect 26384 40403 26413 40409
rect 26528 40412 27476 40440
rect 26384 40400 26390 40403
rect 26528 40372 26556 40412
rect 27448 40384 27476 40412
rect 30742 40400 30748 40452
rect 30800 40440 30806 40452
rect 35360 40440 35388 40480
rect 35621 40477 35633 40480
rect 35667 40508 35679 40511
rect 35986 40508 35992 40520
rect 35667 40480 35992 40508
rect 35667 40477 35679 40480
rect 35621 40471 35679 40477
rect 35986 40468 35992 40480
rect 36044 40468 36050 40520
rect 37645 40511 37703 40517
rect 37645 40477 37657 40511
rect 37691 40508 37703 40511
rect 38010 40508 38016 40520
rect 37691 40480 38016 40508
rect 37691 40477 37703 40480
rect 37645 40471 37703 40477
rect 38010 40468 38016 40480
rect 38068 40468 38074 40520
rect 30800 40412 35388 40440
rect 35437 40443 35495 40449
rect 30800 40400 30806 40412
rect 35437 40409 35449 40443
rect 35483 40409 35495 40443
rect 35437 40403 35495 40409
rect 26068 40344 26556 40372
rect 26697 40375 26755 40381
rect 26697 40341 26709 40375
rect 26743 40372 26755 40375
rect 26786 40372 26792 40384
rect 26743 40344 26792 40372
rect 26743 40341 26755 40344
rect 26697 40335 26755 40341
rect 26786 40332 26792 40344
rect 26844 40332 26850 40384
rect 26878 40332 26884 40384
rect 26936 40372 26942 40384
rect 27157 40375 27215 40381
rect 27157 40372 27169 40375
rect 26936 40344 27169 40372
rect 26936 40332 26942 40344
rect 27157 40341 27169 40344
rect 27203 40341 27215 40375
rect 27157 40335 27215 40341
rect 27430 40332 27436 40384
rect 27488 40332 27494 40384
rect 35452 40372 35480 40403
rect 35526 40400 35532 40452
rect 35584 40400 35590 40452
rect 35802 40400 35808 40452
rect 35860 40400 35866 40452
rect 36906 40400 36912 40452
rect 36964 40440 36970 40452
rect 36964 40412 37228 40440
rect 36964 40400 36970 40412
rect 35820 40372 35848 40400
rect 37200 40384 37228 40412
rect 35452 40344 35848 40372
rect 35894 40332 35900 40384
rect 35952 40332 35958 40384
rect 37182 40332 37188 40384
rect 37240 40332 37246 40384
rect 1104 40282 45172 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 45172 40282
rect 1104 40208 45172 40230
rect 1854 40128 1860 40180
rect 1912 40168 1918 40180
rect 2869 40171 2927 40177
rect 2869 40168 2881 40171
rect 1912 40140 2881 40168
rect 1912 40128 1918 40140
rect 2869 40137 2881 40140
rect 2915 40137 2927 40171
rect 4062 40168 4068 40180
rect 2869 40131 2927 40137
rect 3896 40140 4068 40168
rect 3896 40109 3924 40140
rect 4062 40128 4068 40140
rect 4120 40128 4126 40180
rect 8110 40128 8116 40180
rect 8168 40168 8174 40180
rect 8205 40171 8263 40177
rect 8205 40168 8217 40171
rect 8168 40140 8217 40168
rect 8168 40128 8174 40140
rect 8205 40137 8217 40140
rect 8251 40137 8263 40171
rect 8205 40131 8263 40137
rect 8570 40128 8576 40180
rect 8628 40128 8634 40180
rect 8662 40128 8668 40180
rect 8720 40128 8726 40180
rect 9766 40168 9772 40180
rect 8864 40140 9772 40168
rect 3881 40103 3939 40109
rect 3881 40069 3893 40103
rect 3927 40069 3939 40103
rect 3881 40063 3939 40069
rect 4338 40060 4344 40112
rect 4396 40060 4402 40112
rect 8018 40100 8024 40112
rect 7866 40072 8024 40100
rect 8018 40060 8024 40072
rect 8076 40060 8082 40112
rect 8588 40100 8616 40128
rect 8128 40072 8616 40100
rect 3602 39992 3608 40044
rect 3660 39992 3666 40044
rect 6178 39992 6184 40044
rect 6236 40032 6242 40044
rect 6365 40035 6423 40041
rect 6365 40032 6377 40035
rect 6236 40004 6377 40032
rect 6236 39992 6242 40004
rect 6365 40001 6377 40004
rect 6411 40001 6423 40035
rect 6365 39995 6423 40001
rect 3510 39924 3516 39976
rect 3568 39924 3574 39976
rect 3620 39964 3648 39992
rect 3970 39964 3976 39976
rect 3620 39936 3976 39964
rect 3970 39924 3976 39936
rect 4028 39924 4034 39976
rect 5353 39967 5411 39973
rect 5353 39933 5365 39967
rect 5399 39964 5411 39967
rect 5445 39967 5503 39973
rect 5445 39964 5457 39967
rect 5399 39936 5457 39964
rect 5399 39933 5411 39936
rect 5353 39927 5411 39933
rect 5445 39933 5457 39936
rect 5491 39933 5503 39967
rect 5445 39927 5503 39933
rect 6638 39924 6644 39976
rect 6696 39924 6702 39976
rect 8128 39973 8156 40072
rect 8384 40035 8442 40041
rect 8384 40032 8396 40035
rect 8312 40004 8396 40032
rect 8113 39967 8171 39973
rect 8113 39933 8125 39967
rect 8159 39933 8171 39967
rect 8113 39927 8171 39933
rect 8312 39964 8340 40004
rect 8384 40001 8396 40004
rect 8430 40001 8442 40035
rect 8384 39995 8442 40001
rect 8478 39992 8484 40044
rect 8536 39992 8542 40044
rect 8570 39992 8576 40044
rect 8628 39992 8634 40044
rect 8680 40041 8708 40128
rect 8864 40041 8892 40140
rect 9766 40128 9772 40140
rect 9824 40128 9830 40180
rect 10410 40128 10416 40180
rect 10468 40128 10474 40180
rect 11882 40128 11888 40180
rect 11940 40168 11946 40180
rect 11977 40171 12035 40177
rect 11977 40168 11989 40171
rect 11940 40140 11989 40168
rect 11940 40128 11946 40140
rect 11977 40137 11989 40140
rect 12023 40137 12035 40171
rect 11977 40131 12035 40137
rect 13449 40171 13507 40177
rect 13449 40137 13461 40171
rect 13495 40168 13507 40171
rect 13722 40168 13728 40180
rect 13495 40140 13728 40168
rect 13495 40137 13507 40140
rect 13449 40131 13507 40137
rect 13722 40128 13728 40140
rect 13780 40128 13786 40180
rect 14642 40168 14648 40180
rect 14200 40140 14648 40168
rect 10428 40100 10456 40128
rect 10350 40072 10456 40100
rect 10781 40103 10839 40109
rect 10781 40069 10793 40103
rect 10827 40100 10839 40103
rect 12250 40100 12256 40112
rect 10827 40072 12256 40100
rect 10827 40069 10839 40072
rect 10781 40063 10839 40069
rect 12250 40060 12256 40072
rect 12308 40060 12314 40112
rect 13081 40103 13139 40109
rect 13081 40069 13093 40103
rect 13127 40100 13139 40103
rect 14200 40100 14228 40140
rect 14642 40128 14648 40140
rect 14700 40168 14706 40180
rect 15289 40171 15347 40177
rect 15289 40168 15301 40171
rect 14700 40140 15301 40168
rect 14700 40128 14706 40140
rect 15289 40137 15301 40140
rect 15335 40137 15347 40171
rect 15289 40131 15347 40137
rect 16485 40171 16543 40177
rect 16485 40137 16497 40171
rect 16531 40168 16543 40171
rect 17678 40168 17684 40180
rect 16531 40140 17684 40168
rect 16531 40137 16543 40140
rect 16485 40131 16543 40137
rect 17678 40128 17684 40140
rect 17736 40128 17742 40180
rect 21174 40168 21180 40180
rect 17788 40140 21180 40168
rect 13127 40072 14228 40100
rect 13127 40069 13139 40072
rect 13081 40063 13139 40069
rect 14458 40060 14464 40112
rect 14516 40060 14522 40112
rect 16942 40060 16948 40112
rect 17000 40100 17006 40112
rect 17788 40100 17816 40140
rect 21174 40128 21180 40140
rect 21232 40128 21238 40180
rect 22738 40128 22744 40180
rect 22796 40168 22802 40180
rect 23201 40171 23259 40177
rect 23201 40168 23213 40171
rect 22796 40140 23213 40168
rect 22796 40128 22802 40140
rect 23201 40137 23213 40140
rect 23247 40168 23259 40171
rect 26234 40168 26240 40180
rect 23247 40140 26240 40168
rect 23247 40137 23259 40140
rect 23201 40131 23259 40137
rect 26234 40128 26240 40140
rect 26292 40128 26298 40180
rect 27430 40128 27436 40180
rect 27488 40128 27494 40180
rect 27985 40171 28043 40177
rect 27985 40137 27997 40171
rect 28031 40168 28043 40171
rect 28166 40168 28172 40180
rect 28031 40140 28172 40168
rect 28031 40137 28043 40140
rect 27985 40131 28043 40137
rect 28166 40128 28172 40140
rect 28224 40128 28230 40180
rect 28258 40128 28264 40180
rect 28316 40128 28322 40180
rect 35250 40128 35256 40180
rect 35308 40128 35314 40180
rect 35526 40128 35532 40180
rect 35584 40168 35590 40180
rect 35713 40171 35771 40177
rect 35713 40168 35725 40171
rect 35584 40140 35725 40168
rect 35584 40128 35590 40140
rect 35713 40137 35725 40140
rect 35759 40137 35771 40171
rect 40589 40171 40647 40177
rect 40589 40168 40601 40171
rect 35713 40131 35771 40137
rect 40512 40140 40601 40168
rect 20622 40100 20628 40112
rect 17000 40072 17816 40100
rect 19826 40072 20628 40100
rect 17000 40060 17006 40072
rect 20622 40060 20628 40072
rect 20680 40060 20686 40112
rect 20898 40100 20904 40112
rect 20824 40072 20904 40100
rect 8680 40035 8759 40041
rect 8680 40004 8713 40035
rect 8701 40001 8713 40004
rect 8747 40001 8759 40035
rect 8701 39995 8759 40001
rect 8849 40035 8907 40041
rect 8849 40001 8861 40035
rect 8895 40001 8907 40035
rect 8849 39995 8907 40001
rect 11146 39992 11152 40044
rect 11204 39992 11210 40044
rect 15841 40035 15899 40041
rect 15841 40001 15853 40035
rect 15887 40001 15899 40035
rect 15841 39995 15899 40001
rect 9214 39964 9220 39976
rect 8312 39936 9220 39964
rect 8312 39896 8340 39936
rect 9214 39924 9220 39936
rect 9272 39924 9278 39976
rect 9309 39967 9367 39973
rect 9309 39933 9321 39967
rect 9355 39964 9367 39967
rect 10042 39964 10048 39976
rect 9355 39936 10048 39964
rect 9355 39933 9367 39936
rect 9309 39927 9367 39933
rect 10042 39924 10048 39936
rect 10100 39924 10106 39976
rect 11054 39924 11060 39976
rect 11112 39924 11118 39976
rect 8128 39868 8340 39896
rect 8128 39840 8156 39868
rect 6086 39788 6092 39840
rect 6144 39788 6150 39840
rect 8110 39788 8116 39840
rect 8168 39788 8174 39840
rect 10778 39788 10784 39840
rect 10836 39828 10842 39840
rect 11072 39828 11100 39924
rect 10836 39800 11100 39828
rect 11164 39828 11192 39992
rect 12434 39924 12440 39976
rect 12492 39964 12498 39976
rect 12529 39967 12587 39973
rect 12529 39964 12541 39967
rect 12492 39936 12541 39964
rect 12492 39924 12498 39936
rect 12529 39933 12541 39936
rect 12575 39933 12587 39967
rect 12529 39927 12587 39933
rect 12802 39924 12808 39976
rect 12860 39924 12866 39976
rect 12986 39924 12992 39976
rect 13044 39924 13050 39976
rect 13541 39967 13599 39973
rect 13541 39933 13553 39967
rect 13587 39964 13599 39967
rect 13817 39967 13875 39973
rect 13587 39936 13676 39964
rect 13587 39933 13599 39936
rect 13541 39927 13599 39933
rect 13648 39840 13676 39936
rect 13817 39933 13829 39967
rect 13863 39964 13875 39967
rect 13906 39964 13912 39976
rect 13863 39936 13912 39964
rect 13863 39933 13875 39936
rect 13817 39927 13875 39933
rect 13906 39924 13912 39936
rect 13964 39924 13970 39976
rect 15378 39964 15384 39976
rect 14844 39936 15384 39964
rect 13538 39828 13544 39840
rect 11164 39800 13544 39828
rect 10836 39788 10842 39800
rect 13538 39788 13544 39800
rect 13596 39788 13602 39840
rect 13630 39788 13636 39840
rect 13688 39828 13694 39840
rect 14844 39828 14872 39936
rect 15378 39924 15384 39936
rect 15436 39924 15442 39976
rect 15856 39964 15884 39995
rect 15930 39992 15936 40044
rect 15988 40032 15994 40044
rect 15988 40004 16033 40032
rect 15988 39992 15994 40004
rect 16114 39992 16120 40044
rect 16172 39992 16178 40044
rect 16206 39992 16212 40044
rect 16264 39992 16270 40044
rect 16306 40035 16364 40041
rect 16306 40001 16318 40035
rect 16352 40001 16364 40035
rect 16306 39995 16364 40001
rect 17037 40035 17095 40041
rect 17037 40001 17049 40035
rect 17083 40030 17095 40035
rect 17126 40030 17132 40044
rect 17083 40002 17132 40030
rect 17083 40001 17095 40002
rect 17037 39995 17095 40001
rect 15856 39936 15967 39964
rect 13688 39800 14872 39828
rect 15939 39828 15967 39936
rect 16022 39924 16028 39976
rect 16080 39964 16086 39976
rect 16321 39964 16349 39995
rect 17126 39992 17132 40002
rect 17184 39992 17190 40044
rect 18325 40035 18383 40041
rect 18325 40032 18337 40035
rect 17236 40004 18337 40032
rect 16080 39936 16349 39964
rect 16080 39924 16086 39936
rect 16321 39896 16349 39936
rect 16942 39896 16948 39908
rect 16321 39868 16948 39896
rect 16942 39856 16948 39868
rect 17000 39856 17006 39908
rect 17236 39828 17264 40004
rect 18325 40001 18337 40004
rect 18371 40001 18383 40035
rect 18325 39995 18383 40001
rect 18509 40035 18567 40041
rect 18509 40001 18521 40035
rect 18555 40001 18567 40035
rect 18509 39995 18567 40001
rect 20533 40035 20591 40041
rect 20533 40001 20545 40035
rect 20579 40032 20591 40035
rect 20714 40032 20720 40044
rect 20579 40004 20720 40032
rect 20579 40001 20591 40004
rect 20533 39995 20591 40001
rect 18524 39964 18552 39995
rect 20714 39992 20720 40004
rect 20772 39992 20778 40044
rect 18340 39936 18552 39964
rect 18693 39967 18751 39973
rect 18340 39840 18368 39936
rect 18693 39933 18705 39967
rect 18739 39964 18751 39967
rect 20257 39967 20315 39973
rect 18739 39936 18828 39964
rect 18739 39933 18751 39936
rect 18693 39927 18751 39933
rect 18800 39840 18828 39936
rect 20257 39933 20269 39967
rect 20303 39964 20315 39967
rect 20824 39964 20852 40072
rect 20898 40060 20904 40072
rect 20956 40060 20962 40112
rect 22373 40103 22431 40109
rect 22373 40069 22385 40103
rect 22419 40100 22431 40103
rect 23293 40103 23351 40109
rect 23293 40100 23305 40103
rect 22419 40072 23305 40100
rect 22419 40069 22431 40072
rect 22373 40063 22431 40069
rect 23293 40069 23305 40072
rect 23339 40100 23351 40103
rect 23845 40103 23903 40109
rect 23845 40100 23857 40103
rect 23339 40072 23857 40100
rect 23339 40069 23351 40072
rect 23293 40063 23351 40069
rect 23845 40069 23857 40072
rect 23891 40100 23903 40103
rect 24029 40103 24087 40109
rect 24029 40100 24041 40103
rect 23891 40072 24041 40100
rect 23891 40069 23903 40072
rect 23845 40063 23903 40069
rect 24029 40069 24041 40072
rect 24075 40069 24087 40103
rect 27448 40100 27476 40128
rect 24029 40063 24087 40069
rect 26804 40072 27476 40100
rect 23474 39992 23480 40044
rect 23532 40032 23538 40044
rect 26804 40041 26832 40072
rect 27614 40060 27620 40112
rect 27672 40060 27678 40112
rect 28276 40100 28304 40128
rect 40512 40112 40540 40140
rect 40589 40137 40601 40140
rect 40635 40137 40647 40171
rect 40589 40131 40647 40137
rect 28092 40072 28304 40100
rect 24213 40035 24271 40041
rect 24213 40032 24225 40035
rect 23532 40004 24225 40032
rect 23532 39992 23538 40004
rect 24213 40001 24225 40004
rect 24259 40001 24271 40035
rect 24213 39995 24271 40001
rect 26789 40035 26847 40041
rect 26789 40001 26801 40035
rect 26835 40001 26847 40035
rect 26789 39995 26847 40001
rect 20303 39936 20852 39964
rect 20303 39933 20315 39936
rect 20257 39927 20315 39933
rect 20898 39924 20904 39976
rect 20956 39924 20962 39976
rect 22097 39899 22155 39905
rect 22097 39896 22109 39899
rect 21100 39868 22109 39896
rect 21100 39840 21128 39868
rect 22097 39865 22109 39868
rect 22143 39865 22155 39899
rect 24228 39896 24256 39995
rect 27154 39992 27160 40044
rect 27212 39992 27218 40044
rect 27338 39992 27344 40044
rect 27396 40032 27402 40044
rect 27801 40035 27859 40041
rect 27801 40032 27813 40035
rect 27396 40004 27813 40032
rect 27396 39992 27402 40004
rect 27801 40001 27813 40004
rect 27847 40032 27859 40035
rect 27890 40032 27896 40044
rect 27847 40004 27896 40032
rect 27847 40001 27859 40004
rect 27801 39995 27859 40001
rect 27890 39992 27896 40004
rect 27948 39992 27954 40044
rect 28092 40041 28120 40072
rect 30926 40060 30932 40112
rect 30984 40100 30990 40112
rect 34054 40100 34060 40112
rect 30984 40072 33272 40100
rect 30984 40060 30990 40072
rect 28077 40035 28135 40041
rect 28077 40001 28089 40035
rect 28123 40001 28135 40035
rect 28077 39995 28135 40001
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39964 24455 39967
rect 24578 39964 24584 39976
rect 24443 39936 24584 39964
rect 24443 39933 24455 39936
rect 24397 39927 24455 39933
rect 24578 39924 24584 39936
rect 24636 39924 24642 39976
rect 26697 39967 26755 39973
rect 26697 39933 26709 39967
rect 26743 39964 26755 39967
rect 26878 39964 26884 39976
rect 26743 39936 26884 39964
rect 26743 39933 26755 39936
rect 26697 39927 26755 39933
rect 26878 39924 26884 39936
rect 26936 39924 26942 39976
rect 27249 39967 27307 39973
rect 27249 39933 27261 39967
rect 27295 39933 27307 39967
rect 27249 39927 27307 39933
rect 27433 39967 27491 39973
rect 27433 39933 27445 39967
rect 27479 39964 27491 39967
rect 28258 39964 28264 39976
rect 27479 39936 28264 39964
rect 27479 39933 27491 39936
rect 27433 39927 27491 39933
rect 27264 39896 27292 39927
rect 28258 39924 28264 39936
rect 28316 39924 28322 39976
rect 33244 39964 33272 40072
rect 33336 40072 34060 40100
rect 33336 40041 33364 40072
rect 34054 40060 34060 40072
rect 34112 40100 34118 40112
rect 34112 40072 34928 40100
rect 34112 40060 34118 40072
rect 33321 40035 33379 40041
rect 33321 40001 33333 40035
rect 33367 40001 33379 40035
rect 33321 39995 33379 40001
rect 34149 40035 34207 40041
rect 34149 40001 34161 40035
rect 34195 40032 34207 40035
rect 34330 40032 34336 40044
rect 34195 40004 34336 40032
rect 34195 40001 34207 40004
rect 34149 39995 34207 40001
rect 34330 39992 34336 40004
rect 34388 39992 34394 40044
rect 34900 40041 34928 40072
rect 40494 40060 40500 40112
rect 40552 40060 40558 40112
rect 34885 40035 34943 40041
rect 34885 40001 34897 40035
rect 34931 40001 34943 40035
rect 34885 39995 34943 40001
rect 35894 39992 35900 40044
rect 35952 40032 35958 40044
rect 36265 40035 36323 40041
rect 36265 40032 36277 40035
rect 35952 40004 36277 40032
rect 35952 39992 35958 40004
rect 36265 40001 36277 40004
rect 36311 40001 36323 40035
rect 40678 40032 40684 40044
rect 40250 40004 40684 40032
rect 36265 39995 36323 40001
rect 40678 39992 40684 40004
rect 40736 39992 40742 40044
rect 34241 39967 34299 39973
rect 34241 39964 34253 39967
rect 33244 39936 34253 39964
rect 34241 39933 34253 39936
rect 34287 39964 34299 39967
rect 34422 39964 34428 39976
rect 34287 39936 34428 39964
rect 34287 39933 34299 39936
rect 34241 39927 34299 39933
rect 34422 39924 34428 39936
rect 34480 39924 34486 39976
rect 34977 39967 35035 39973
rect 34977 39933 34989 39967
rect 35023 39964 35035 39967
rect 35434 39964 35440 39976
rect 35023 39936 35440 39964
rect 35023 39933 35035 39936
rect 34977 39927 35035 39933
rect 35434 39924 35440 39936
rect 35492 39924 35498 39976
rect 38010 39924 38016 39976
rect 38068 39964 38074 39976
rect 38841 39967 38899 39973
rect 38841 39964 38853 39967
rect 38068 39936 38853 39964
rect 38068 39924 38074 39936
rect 38841 39933 38853 39936
rect 38887 39933 38899 39967
rect 38841 39927 38899 39933
rect 39114 39924 39120 39976
rect 39172 39924 39178 39976
rect 27522 39896 27528 39908
rect 24228 39868 26832 39896
rect 27264 39868 27528 39896
rect 22097 39859 22155 39865
rect 15939 39800 17264 39828
rect 13688 39788 13694 39800
rect 17586 39788 17592 39840
rect 17644 39788 17650 39840
rect 18322 39788 18328 39840
rect 18380 39788 18386 39840
rect 18782 39788 18788 39840
rect 18840 39788 18846 39840
rect 21082 39788 21088 39840
rect 21140 39788 21146 39840
rect 21542 39788 21548 39840
rect 21600 39788 21606 39840
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 23753 39831 23811 39837
rect 23753 39828 23765 39831
rect 23716 39800 23765 39828
rect 23716 39788 23722 39800
rect 23753 39797 23765 39800
rect 23799 39828 23811 39831
rect 26326 39828 26332 39840
rect 23799 39800 26332 39828
rect 23799 39797 23811 39800
rect 23753 39791 23811 39797
rect 26326 39788 26332 39800
rect 26384 39788 26390 39840
rect 26421 39831 26479 39837
rect 26421 39797 26433 39831
rect 26467 39828 26479 39831
rect 26510 39828 26516 39840
rect 26467 39800 26516 39828
rect 26467 39797 26479 39800
rect 26421 39791 26479 39797
rect 26510 39788 26516 39800
rect 26568 39788 26574 39840
rect 26804 39837 26832 39868
rect 27522 39856 27528 39868
rect 27580 39856 27586 39908
rect 26789 39831 26847 39837
rect 26789 39797 26801 39831
rect 26835 39828 26847 39831
rect 26973 39831 27031 39837
rect 26973 39828 26985 39831
rect 26835 39800 26985 39828
rect 26835 39797 26847 39800
rect 26789 39791 26847 39797
rect 26973 39797 26985 39800
rect 27019 39828 27031 39831
rect 30282 39828 30288 39840
rect 27019 39800 30288 39828
rect 27019 39797 27031 39800
rect 26973 39791 27031 39797
rect 30282 39788 30288 39800
rect 30340 39788 30346 39840
rect 1104 39738 45172 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 45172 39738
rect 1104 39664 45172 39686
rect 3970 39584 3976 39636
rect 4028 39624 4034 39636
rect 4249 39627 4307 39633
rect 4249 39624 4261 39627
rect 4028 39596 4261 39624
rect 4028 39584 4034 39596
rect 4249 39593 4261 39596
rect 4295 39624 4307 39627
rect 6178 39624 6184 39636
rect 4295 39596 6184 39624
rect 4295 39593 4307 39596
rect 4249 39587 4307 39593
rect 6178 39584 6184 39596
rect 6236 39584 6242 39636
rect 6638 39584 6644 39636
rect 6696 39624 6702 39636
rect 6917 39627 6975 39633
rect 6917 39624 6929 39627
rect 6696 39596 6929 39624
rect 6696 39584 6702 39596
rect 6917 39593 6929 39596
rect 6963 39593 6975 39627
rect 6917 39587 6975 39593
rect 8018 39584 8024 39636
rect 8076 39624 8082 39636
rect 8570 39624 8576 39636
rect 8076 39596 8576 39624
rect 8076 39584 8082 39596
rect 8570 39584 8576 39596
rect 8628 39584 8634 39636
rect 9677 39627 9735 39633
rect 9677 39593 9689 39627
rect 9723 39624 9735 39627
rect 9766 39624 9772 39636
rect 9723 39596 9772 39624
rect 9723 39593 9735 39596
rect 9677 39587 9735 39593
rect 9766 39584 9772 39596
rect 9824 39584 9830 39636
rect 12345 39627 12403 39633
rect 12345 39593 12357 39627
rect 12391 39624 12403 39627
rect 12434 39624 12440 39636
rect 12391 39596 12440 39624
rect 12391 39593 12403 39596
rect 12345 39587 12403 39593
rect 12434 39584 12440 39596
rect 12492 39584 12498 39636
rect 13538 39584 13544 39636
rect 13596 39624 13602 39636
rect 16761 39627 16819 39633
rect 13596 39596 16712 39624
rect 13596 39584 13602 39596
rect 4522 39516 4528 39568
rect 4580 39556 4586 39568
rect 4798 39556 4804 39568
rect 4580 39528 4804 39556
rect 4580 39516 4586 39528
rect 4798 39516 4804 39528
rect 4856 39556 4862 39568
rect 8036 39556 8064 39584
rect 4856 39528 8064 39556
rect 4856 39516 4862 39528
rect 8202 39516 8208 39568
rect 8260 39556 8266 39568
rect 16684 39556 16712 39596
rect 16761 39593 16773 39627
rect 16807 39624 16819 39627
rect 17126 39624 17132 39636
rect 16807 39596 17132 39624
rect 16807 39593 16819 39596
rect 16761 39587 16819 39593
rect 17126 39584 17132 39596
rect 17184 39584 17190 39636
rect 20533 39627 20591 39633
rect 20533 39593 20545 39627
rect 20579 39624 20591 39627
rect 20898 39624 20904 39636
rect 20579 39596 20904 39624
rect 20579 39593 20591 39596
rect 20533 39587 20591 39593
rect 20898 39584 20904 39596
rect 20956 39584 20962 39636
rect 26145 39627 26203 39633
rect 26145 39593 26157 39627
rect 26191 39624 26203 39627
rect 27522 39624 27528 39636
rect 26191 39596 27528 39624
rect 26191 39593 26203 39596
rect 26145 39587 26203 39593
rect 27522 39584 27528 39596
rect 27580 39584 27586 39636
rect 27890 39584 27896 39636
rect 27948 39624 27954 39636
rect 28261 39627 28319 39633
rect 28261 39624 28273 39627
rect 27948 39596 28273 39624
rect 27948 39584 27954 39596
rect 28261 39593 28273 39596
rect 28307 39593 28319 39627
rect 28261 39587 28319 39593
rect 18322 39556 18328 39568
rect 8260 39528 9904 39556
rect 16684 39528 18328 39556
rect 8260 39516 8266 39528
rect 6362 39488 6368 39500
rect 5552 39460 6368 39488
rect 2590 39380 2596 39432
rect 2648 39420 2654 39432
rect 5552 39429 5580 39460
rect 6362 39448 6368 39460
rect 6420 39488 6426 39500
rect 6420 39460 9076 39488
rect 6420 39448 6426 39460
rect 9048 39432 9076 39460
rect 3053 39423 3111 39429
rect 3053 39420 3065 39423
rect 2648 39392 3065 39420
rect 2648 39380 2654 39392
rect 3053 39389 3065 39392
rect 3099 39389 3111 39423
rect 3053 39383 3111 39389
rect 5537 39423 5595 39429
rect 5537 39389 5549 39423
rect 5583 39389 5595 39423
rect 5537 39383 5595 39389
rect 7561 39423 7619 39429
rect 7561 39389 7573 39423
rect 7607 39420 7619 39423
rect 7832 39423 7890 39429
rect 7607 39392 7696 39420
rect 7607 39389 7619 39392
rect 7561 39383 7619 39389
rect 2498 39244 2504 39296
rect 2556 39244 2562 39296
rect 3142 39244 3148 39296
rect 3200 39284 3206 39296
rect 5902 39284 5908 39296
rect 3200 39256 5908 39284
rect 3200 39244 3206 39256
rect 5902 39244 5908 39256
rect 5960 39244 5966 39296
rect 7668 39293 7696 39392
rect 7832 39389 7844 39423
rect 7878 39420 7890 39423
rect 8110 39420 8116 39432
rect 7878 39392 8116 39420
rect 7878 39389 7890 39392
rect 7832 39383 7890 39389
rect 8110 39380 8116 39392
rect 8168 39380 8174 39432
rect 8204 39423 8262 39429
rect 8204 39389 8216 39423
rect 8250 39389 8262 39423
rect 8204 39383 8262 39389
rect 7929 39355 7987 39361
rect 7929 39321 7941 39355
rect 7975 39321 7987 39355
rect 7929 39315 7987 39321
rect 7653 39287 7711 39293
rect 7653 39253 7665 39287
rect 7699 39253 7711 39287
rect 7944 39284 7972 39315
rect 8018 39312 8024 39364
rect 8076 39312 8082 39364
rect 8220 39352 8248 39383
rect 8294 39380 8300 39432
rect 8352 39380 8358 39432
rect 8386 39380 8392 39432
rect 8444 39380 8450 39432
rect 8938 39380 8944 39432
rect 8996 39380 9002 39432
rect 9030 39380 9036 39432
rect 9088 39380 9094 39432
rect 9876 39429 9904 39528
rect 18322 39516 18328 39528
rect 18380 39556 18386 39568
rect 20346 39556 20352 39568
rect 18380 39528 20352 39556
rect 18380 39516 18386 39528
rect 20346 39516 20352 39528
rect 20404 39516 20410 39568
rect 30193 39559 30251 39565
rect 30193 39556 30205 39559
rect 29656 39528 30205 39556
rect 10042 39448 10048 39500
rect 10100 39448 10106 39500
rect 13630 39448 13636 39500
rect 13688 39448 13694 39500
rect 15378 39448 15384 39500
rect 15436 39448 15442 39500
rect 20364 39488 20392 39516
rect 21634 39488 21640 39500
rect 20364 39460 21640 39488
rect 21634 39448 21640 39460
rect 21692 39448 21698 39500
rect 24394 39448 24400 39500
rect 24452 39488 24458 39500
rect 26513 39491 26571 39497
rect 26513 39488 26525 39491
rect 24452 39460 26525 39488
rect 24452 39448 24458 39460
rect 26513 39457 26525 39460
rect 26559 39457 26571 39491
rect 26513 39451 26571 39457
rect 26786 39448 26792 39500
rect 26844 39448 26850 39500
rect 29656 39497 29684 39528
rect 30193 39525 30205 39528
rect 30239 39556 30251 39559
rect 30282 39556 30288 39568
rect 30239 39528 30288 39556
rect 30239 39525 30251 39528
rect 30193 39519 30251 39525
rect 30282 39516 30288 39528
rect 30340 39516 30346 39568
rect 36173 39559 36231 39565
rect 36173 39525 36185 39559
rect 36219 39525 36231 39559
rect 36173 39519 36231 39525
rect 29641 39491 29699 39497
rect 29641 39457 29653 39491
rect 29687 39457 29699 39491
rect 29641 39451 29699 39457
rect 30006 39448 30012 39500
rect 30064 39488 30070 39500
rect 30374 39488 30380 39500
rect 30064 39460 30380 39488
rect 30064 39448 30070 39460
rect 9861 39423 9919 39429
rect 9861 39389 9873 39423
rect 9907 39389 9919 39423
rect 9861 39383 9919 39389
rect 10778 39380 10784 39432
rect 10836 39420 10842 39432
rect 10965 39423 11023 39429
rect 10965 39420 10977 39423
rect 10836 39392 10977 39420
rect 10836 39380 10842 39392
rect 10965 39389 10977 39392
rect 11011 39389 11023 39423
rect 10965 39383 11023 39389
rect 12437 39423 12495 39429
rect 12437 39389 12449 39423
rect 12483 39420 12495 39423
rect 13648 39420 13676 39448
rect 12483 39392 13676 39420
rect 12483 39389 12495 39392
rect 12437 39383 12495 39389
rect 15102 39380 15108 39432
rect 15160 39380 15166 39432
rect 17678 39380 17684 39432
rect 17736 39380 17742 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 19613 39423 19671 39429
rect 19613 39420 19625 39423
rect 19484 39392 19625 39420
rect 19484 39380 19490 39392
rect 19613 39389 19625 39392
rect 19659 39389 19671 39423
rect 19613 39383 19671 39389
rect 22278 39380 22284 39432
rect 22336 39380 22342 39432
rect 26418 39380 26424 39432
rect 26476 39380 26482 39432
rect 29822 39380 29828 39432
rect 29880 39380 29886 39432
rect 30116 39429 30144 39460
rect 30374 39448 30380 39460
rect 30432 39448 30438 39500
rect 32214 39448 32220 39500
rect 32272 39448 32278 39500
rect 36188 39488 36216 39519
rect 37737 39491 37795 39497
rect 37737 39488 37749 39491
rect 36188 39460 37749 39488
rect 37737 39457 37749 39460
rect 37783 39457 37795 39491
rect 37737 39451 37795 39457
rect 39298 39448 39304 39500
rect 39356 39488 39362 39500
rect 41601 39491 41659 39497
rect 39356 39460 39528 39488
rect 39356 39448 39362 39460
rect 30101 39423 30159 39429
rect 30101 39389 30113 39423
rect 30147 39389 30159 39423
rect 30101 39383 30159 39389
rect 30190 39380 30196 39432
rect 30248 39420 30254 39432
rect 30285 39423 30343 39429
rect 30285 39420 30297 39423
rect 30248 39392 30297 39420
rect 30248 39380 30254 39392
rect 30285 39389 30297 39392
rect 30331 39389 30343 39423
rect 30285 39383 30343 39389
rect 8404 39352 8432 39380
rect 8220 39324 8432 39352
rect 11232 39355 11290 39361
rect 11232 39321 11244 39355
rect 11278 39352 11290 39355
rect 11514 39352 11520 39364
rect 11278 39324 11520 39352
rect 11278 39321 11290 39324
rect 11232 39315 11290 39321
rect 11514 39312 11520 39324
rect 11572 39312 11578 39364
rect 12704 39355 12762 39361
rect 12704 39321 12716 39355
rect 12750 39352 12762 39355
rect 14182 39352 14188 39364
rect 12750 39324 14188 39352
rect 12750 39321 12762 39324
rect 12704 39315 12762 39321
rect 14182 39312 14188 39324
rect 14240 39312 14246 39364
rect 15626 39355 15684 39361
rect 15626 39352 15638 39355
rect 15304 39324 15638 39352
rect 8110 39284 8116 39296
rect 7944 39256 8116 39284
rect 7653 39247 7711 39253
rect 8110 39244 8116 39256
rect 8168 39244 8174 39296
rect 8478 39244 8484 39296
rect 8536 39284 8542 39296
rect 9030 39284 9036 39296
rect 8536 39256 9036 39284
rect 8536 39244 8542 39256
rect 9030 39244 9036 39256
rect 9088 39284 9094 39296
rect 9585 39287 9643 39293
rect 9585 39284 9597 39287
rect 9088 39256 9597 39284
rect 9088 39244 9094 39256
rect 9585 39253 9597 39256
rect 9631 39253 9643 39287
rect 9585 39247 9643 39253
rect 13814 39244 13820 39296
rect 13872 39244 13878 39296
rect 15304 39293 15332 39324
rect 15626 39321 15638 39324
rect 15672 39321 15684 39355
rect 15626 39315 15684 39321
rect 19978 39312 19984 39364
rect 20036 39352 20042 39364
rect 20036 39324 20668 39352
rect 20036 39312 20042 39324
rect 15289 39287 15347 39293
rect 15289 39253 15301 39287
rect 15335 39253 15347 39287
rect 15289 39247 15347 39253
rect 17034 39244 17040 39296
rect 17092 39284 17098 39296
rect 17129 39287 17187 39293
rect 17129 39284 17141 39287
rect 17092 39256 17141 39284
rect 17092 39244 17098 39256
rect 17129 39253 17141 39256
rect 17175 39253 17187 39287
rect 17129 39247 17187 39253
rect 19150 39244 19156 39296
rect 19208 39284 19214 39296
rect 20254 39284 20260 39296
rect 19208 39256 20260 39284
rect 19208 39244 19214 39256
rect 20254 39244 20260 39256
rect 20312 39244 20318 39296
rect 20640 39284 20668 39324
rect 20714 39312 20720 39364
rect 20772 39352 20778 39364
rect 20772 39324 20838 39352
rect 20772 39312 20778 39324
rect 22002 39312 22008 39364
rect 22060 39312 22066 39364
rect 22465 39355 22523 39361
rect 22465 39321 22477 39355
rect 22511 39352 22523 39355
rect 22646 39352 22652 39364
rect 22511 39324 22652 39352
rect 22511 39321 22523 39324
rect 22465 39315 22523 39321
rect 22646 39312 22652 39324
rect 22704 39312 22710 39364
rect 24670 39312 24676 39364
rect 24728 39312 24734 39364
rect 30392 39352 30420 39448
rect 35618 39380 35624 39432
rect 35676 39380 35682 39432
rect 35986 39380 35992 39432
rect 36044 39380 36050 39432
rect 38010 39380 38016 39432
rect 38068 39380 38074 39432
rect 38286 39380 38292 39432
rect 38344 39420 38350 39432
rect 39500 39429 39528 39460
rect 41601 39457 41613 39491
rect 41647 39488 41659 39491
rect 42058 39488 42064 39500
rect 41647 39460 42064 39488
rect 41647 39457 41659 39460
rect 41601 39451 41659 39457
rect 42058 39448 42064 39460
rect 42116 39448 42122 39500
rect 39117 39423 39175 39429
rect 39117 39420 39129 39423
rect 38344 39392 39129 39420
rect 38344 39380 38350 39392
rect 39117 39389 39129 39392
rect 39163 39389 39175 39423
rect 39393 39423 39451 39429
rect 39393 39420 39405 39423
rect 39117 39383 39175 39389
rect 39224 39392 39405 39420
rect 25898 39324 27278 39352
rect 30392 39324 30604 39352
rect 21082 39284 21088 39296
rect 20640 39256 21088 39284
rect 21082 39244 21088 39256
rect 21140 39244 21146 39296
rect 21174 39244 21180 39296
rect 21232 39284 21238 39296
rect 22741 39287 22799 39293
rect 22741 39284 22753 39287
rect 21232 39256 22753 39284
rect 21232 39244 21238 39256
rect 22741 39253 22753 39256
rect 22787 39284 22799 39287
rect 23382 39284 23388 39296
rect 22787 39256 23388 39284
rect 22787 39253 22799 39256
rect 22741 39247 22799 39253
rect 23382 39244 23388 39256
rect 23440 39244 23446 39296
rect 25682 39244 25688 39296
rect 25740 39284 25746 39296
rect 25976 39284 26004 39324
rect 25740 39256 26004 39284
rect 25740 39244 25746 39256
rect 26326 39244 26332 39296
rect 26384 39244 26390 39296
rect 30006 39244 30012 39296
rect 30064 39244 30070 39296
rect 30466 39244 30472 39296
rect 30524 39244 30530 39296
rect 30576 39284 30604 39324
rect 31478 39312 31484 39364
rect 31536 39312 31542 39364
rect 31941 39355 31999 39361
rect 31941 39321 31953 39355
rect 31987 39352 31999 39355
rect 35802 39352 35808 39364
rect 31987 39324 35808 39352
rect 31987 39321 31999 39324
rect 31941 39315 31999 39321
rect 35802 39312 35808 39324
rect 35860 39312 35866 39364
rect 35894 39312 35900 39364
rect 35952 39312 35958 39364
rect 37182 39312 37188 39364
rect 37240 39312 37246 39364
rect 38746 39312 38752 39364
rect 38804 39352 38810 39364
rect 39224 39352 39252 39392
rect 39393 39389 39405 39392
rect 39439 39389 39451 39423
rect 39393 39383 39451 39389
rect 39485 39423 39543 39429
rect 39485 39389 39497 39423
rect 39531 39389 39543 39423
rect 39485 39383 39543 39389
rect 39850 39380 39856 39432
rect 39908 39380 39914 39432
rect 41782 39380 41788 39432
rect 41840 39420 41846 39432
rect 42245 39423 42303 39429
rect 42245 39420 42257 39423
rect 41840 39392 42257 39420
rect 41840 39380 41846 39392
rect 42245 39389 42257 39392
rect 42291 39389 42303 39423
rect 42245 39383 42303 39389
rect 38804 39324 39252 39352
rect 39301 39355 39359 39361
rect 38804 39312 38810 39324
rect 39301 39321 39313 39355
rect 39347 39352 39359 39355
rect 39347 39324 39528 39352
rect 39347 39321 39359 39324
rect 39301 39315 39359 39321
rect 39500 39296 39528 39324
rect 40126 39312 40132 39364
rect 40184 39312 40190 39364
rect 40678 39312 40684 39364
rect 40736 39312 40742 39364
rect 34146 39284 34152 39296
rect 30576 39256 34152 39284
rect 34146 39244 34152 39256
rect 34204 39244 34210 39296
rect 34330 39244 34336 39296
rect 34388 39284 34394 39296
rect 36262 39284 36268 39296
rect 34388 39256 36268 39284
rect 34388 39244 34394 39256
rect 36262 39244 36268 39256
rect 36320 39244 36326 39296
rect 39482 39244 39488 39296
rect 39540 39244 39546 39296
rect 39669 39287 39727 39293
rect 39669 39253 39681 39287
rect 39715 39284 39727 39287
rect 40034 39284 40040 39296
rect 39715 39256 40040 39284
rect 39715 39253 39727 39256
rect 39669 39247 39727 39253
rect 40034 39244 40040 39256
rect 40092 39244 40098 39296
rect 41690 39244 41696 39296
rect 41748 39244 41754 39296
rect 1104 39194 45172 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 45172 39194
rect 1104 39120 45172 39142
rect 2590 39040 2596 39092
rect 2648 39040 2654 39092
rect 4157 39083 4215 39089
rect 4157 39049 4169 39083
rect 4203 39080 4215 39083
rect 4614 39080 4620 39092
rect 4203 39052 4620 39080
rect 4203 39049 4215 39052
rect 4157 39043 4215 39049
rect 4614 39040 4620 39052
rect 4672 39040 4678 39092
rect 8478 39040 8484 39092
rect 8536 39080 8542 39092
rect 8665 39083 8723 39089
rect 8665 39080 8677 39083
rect 8536 39052 8677 39080
rect 8536 39040 8542 39052
rect 8665 39049 8677 39052
rect 8711 39049 8723 39083
rect 8665 39043 8723 39049
rect 11514 39040 11520 39092
rect 11572 39040 11578 39092
rect 11882 39040 11888 39092
rect 11940 39080 11946 39092
rect 12161 39083 12219 39089
rect 12161 39080 12173 39083
rect 11940 39052 12173 39080
rect 11940 39040 11946 39052
rect 12161 39049 12173 39052
rect 12207 39080 12219 39083
rect 12897 39083 12955 39089
rect 12897 39080 12909 39083
rect 12207 39052 12909 39080
rect 12207 39049 12219 39052
rect 12161 39043 12219 39049
rect 12897 39049 12909 39052
rect 12943 39049 12955 39083
rect 12897 39043 12955 39049
rect 12986 39040 12992 39092
rect 13044 39080 13050 39092
rect 13449 39083 13507 39089
rect 13449 39080 13461 39083
rect 13044 39052 13461 39080
rect 13044 39040 13050 39052
rect 13449 39049 13461 39052
rect 13495 39049 13507 39083
rect 13449 39043 13507 39049
rect 13814 39040 13820 39092
rect 13872 39040 13878 39092
rect 14182 39040 14188 39092
rect 14240 39040 14246 39092
rect 15102 39040 15108 39092
rect 15160 39080 15166 39092
rect 15565 39083 15623 39089
rect 15565 39080 15577 39083
rect 15160 39052 15577 39080
rect 15160 39040 15166 39052
rect 15565 39049 15577 39052
rect 15611 39049 15623 39083
rect 15565 39043 15623 39049
rect 15933 39083 15991 39089
rect 15933 39049 15945 39083
rect 15979 39080 15991 39083
rect 16206 39080 16212 39092
rect 15979 39052 16212 39080
rect 15979 39049 15991 39052
rect 15933 39043 15991 39049
rect 16206 39040 16212 39052
rect 16264 39080 16270 39092
rect 17129 39083 17187 39089
rect 17129 39080 17141 39083
rect 16264 39052 17141 39080
rect 16264 39040 16270 39052
rect 17129 39049 17141 39052
rect 17175 39080 17187 39083
rect 17586 39080 17592 39092
rect 17175 39052 17592 39080
rect 17175 39049 17187 39052
rect 17129 39043 17187 39049
rect 17586 39040 17592 39052
rect 17644 39040 17650 39092
rect 19978 39080 19984 39092
rect 17880 39052 19984 39080
rect 6086 39012 6092 39024
rect 4356 38984 4660 39012
rect 2866 38904 2872 38956
rect 2924 38944 2930 38956
rect 4356 38953 4384 38984
rect 2961 38947 3019 38953
rect 2961 38944 2973 38947
rect 2924 38916 2973 38944
rect 2924 38904 2930 38916
rect 2961 38913 2973 38916
rect 3007 38944 3019 38947
rect 3421 38947 3479 38953
rect 3421 38944 3433 38947
rect 3007 38916 3433 38944
rect 3007 38913 3019 38916
rect 2961 38907 3019 38913
rect 3421 38913 3433 38916
rect 3467 38913 3479 38947
rect 3421 38907 3479 38913
rect 4336 38947 4394 38953
rect 4336 38913 4348 38947
rect 4382 38913 4394 38947
rect 4336 38907 4394 38913
rect 4433 38947 4491 38953
rect 4433 38913 4445 38947
rect 4479 38913 4491 38947
rect 4433 38907 4491 38913
rect 3053 38879 3111 38885
rect 3053 38845 3065 38879
rect 3099 38845 3111 38879
rect 3053 38839 3111 38845
rect 3068 38808 3096 38839
rect 3142 38836 3148 38888
rect 3200 38836 3206 38888
rect 3970 38836 3976 38888
rect 4028 38836 4034 38888
rect 4448 38808 4476 38907
rect 4522 38904 4528 38956
rect 4580 38904 4586 38956
rect 4632 38876 4660 38984
rect 4724 38984 6092 39012
rect 4724 38953 4752 38984
rect 6086 38972 6092 38984
rect 6144 38972 6150 39024
rect 8202 39012 8208 39024
rect 7392 38984 8208 39012
rect 7392 38953 7420 38984
rect 8202 38972 8208 38984
rect 8260 38972 8266 39024
rect 12253 39015 12311 39021
rect 12253 38981 12265 39015
rect 12299 39012 12311 39015
rect 12342 39012 12348 39024
rect 12299 38984 12348 39012
rect 12299 38981 12311 38984
rect 12253 38975 12311 38981
rect 12342 38972 12348 38984
rect 12400 38972 12406 39024
rect 4708 38947 4766 38953
rect 4708 38913 4720 38947
rect 4754 38913 4766 38947
rect 4708 38907 4766 38913
rect 4801 38947 4859 38953
rect 4801 38913 4813 38947
rect 4847 38944 4859 38947
rect 7193 38947 7251 38953
rect 7193 38944 7205 38947
rect 4847 38916 7205 38944
rect 4847 38913 4859 38916
rect 4801 38907 4859 38913
rect 7193 38913 7205 38916
rect 7239 38913 7251 38947
rect 7193 38907 7251 38913
rect 7377 38947 7435 38953
rect 7377 38913 7389 38947
rect 7423 38913 7435 38947
rect 7377 38907 7435 38913
rect 7561 38947 7619 38953
rect 7561 38913 7573 38947
rect 7607 38944 7619 38947
rect 8386 38944 8392 38956
rect 7607 38916 8392 38944
rect 7607 38913 7619 38916
rect 7561 38907 7619 38913
rect 8386 38904 8392 38916
rect 8444 38904 8450 38956
rect 8573 38947 8631 38953
rect 8573 38913 8585 38947
rect 8619 38944 8631 38947
rect 10042 38944 10048 38956
rect 8619 38916 10048 38944
rect 8619 38913 8631 38916
rect 8573 38907 8631 38913
rect 10042 38904 10048 38916
rect 10100 38904 10106 38956
rect 11701 38947 11759 38953
rect 11701 38913 11713 38947
rect 11747 38944 11759 38947
rect 13832 38944 13860 39040
rect 17880 39024 17908 39052
rect 15949 38984 17540 39012
rect 14001 38947 14059 38953
rect 14001 38944 14013 38947
rect 11747 38916 11836 38944
rect 13832 38916 14013 38944
rect 11747 38913 11759 38916
rect 11701 38907 11759 38913
rect 4982 38876 4988 38888
rect 4632 38848 4988 38876
rect 4982 38836 4988 38848
rect 5040 38836 5046 38888
rect 8849 38879 8907 38885
rect 8849 38845 8861 38879
rect 8895 38845 8907 38879
rect 8849 38839 8907 38845
rect 4706 38808 4712 38820
rect 3068 38780 3188 38808
rect 4448 38780 4712 38808
rect 3160 38740 3188 38780
rect 4706 38768 4712 38780
rect 4764 38768 4770 38820
rect 5902 38768 5908 38820
rect 5960 38808 5966 38820
rect 8864 38808 8892 38839
rect 9398 38836 9404 38888
rect 9456 38836 9462 38888
rect 11808 38817 11836 38916
rect 14001 38913 14013 38916
rect 14047 38913 14059 38947
rect 14001 38907 14059 38913
rect 14369 38947 14427 38953
rect 14369 38913 14381 38947
rect 14415 38913 14427 38947
rect 14369 38907 14427 38913
rect 12158 38836 12164 38888
rect 12216 38876 12222 38888
rect 12345 38879 12403 38885
rect 12345 38876 12357 38879
rect 12216 38848 12357 38876
rect 12216 38836 12222 38848
rect 12345 38845 12357 38848
rect 12391 38845 12403 38879
rect 12345 38839 12403 38845
rect 12713 38879 12771 38885
rect 12713 38845 12725 38879
rect 12759 38845 12771 38879
rect 14384 38876 14412 38907
rect 12713 38839 12771 38845
rect 13372 38848 14412 38876
rect 15949 38876 15977 38984
rect 16025 38947 16083 38953
rect 16025 38913 16037 38947
rect 16071 38944 16083 38947
rect 16390 38944 16396 38956
rect 16071 38916 16396 38944
rect 16071 38913 16083 38916
rect 16025 38907 16083 38913
rect 16390 38904 16396 38916
rect 16448 38904 16454 38956
rect 17034 38904 17040 38956
rect 17092 38904 17098 38956
rect 16117 38879 16175 38885
rect 16117 38876 16129 38879
rect 15949 38848 16129 38876
rect 5960 38780 8892 38808
rect 5960 38768 5966 38780
rect 5258 38740 5264 38752
rect 3160 38712 5264 38740
rect 5258 38700 5264 38712
rect 5316 38700 5322 38752
rect 8202 38700 8208 38752
rect 8260 38700 8266 38752
rect 8864 38740 8892 38780
rect 11793 38811 11851 38817
rect 11793 38777 11805 38811
rect 11839 38777 11851 38811
rect 11793 38771 11851 38777
rect 12719 38740 12747 38839
rect 13372 38817 13400 38848
rect 16117 38845 16129 38848
rect 16163 38845 16175 38879
rect 17221 38879 17279 38885
rect 17221 38876 17233 38879
rect 16117 38839 16175 38845
rect 16224 38848 17233 38876
rect 13357 38811 13415 38817
rect 13357 38777 13369 38811
rect 13403 38777 13415 38811
rect 13357 38771 13415 38777
rect 16224 38740 16252 38848
rect 17221 38845 17233 38848
rect 17267 38876 17279 38879
rect 17402 38876 17408 38888
rect 17267 38848 17408 38876
rect 17267 38845 17279 38848
rect 17221 38839 17279 38845
rect 17402 38836 17408 38848
rect 17460 38836 17466 38888
rect 8864 38712 16252 38740
rect 16574 38700 16580 38752
rect 16632 38740 16638 38752
rect 16669 38743 16727 38749
rect 16669 38740 16681 38743
rect 16632 38712 16681 38740
rect 16632 38700 16638 38712
rect 16669 38709 16681 38712
rect 16715 38709 16727 38743
rect 17512 38740 17540 38984
rect 17862 38972 17868 39024
rect 17920 38972 17926 39024
rect 18782 38972 18788 39024
rect 18840 39012 18846 39024
rect 19812 39021 19840 39052
rect 19978 39040 19984 39052
rect 20036 39040 20042 39092
rect 20162 39040 20168 39092
rect 20220 39040 20226 39092
rect 20254 39040 20260 39092
rect 20312 39040 20318 39092
rect 20346 39040 20352 39092
rect 20404 39080 20410 39092
rect 20404 39052 20576 39080
rect 20404 39040 20410 39052
rect 19797 39015 19855 39021
rect 18840 38984 19656 39012
rect 18840 38972 18846 38984
rect 18049 38947 18107 38953
rect 18049 38913 18061 38947
rect 18095 38913 18107 38947
rect 18049 38907 18107 38913
rect 18316 38947 18374 38953
rect 18316 38913 18328 38947
rect 18362 38944 18374 38947
rect 18598 38944 18604 38956
rect 18362 38916 18604 38944
rect 18362 38913 18374 38916
rect 18316 38907 18374 38913
rect 17586 38768 17592 38820
rect 17644 38808 17650 38820
rect 18064 38808 18092 38907
rect 18598 38904 18604 38916
rect 18656 38904 18662 38956
rect 19426 38904 19432 38956
rect 19484 38904 19490 38956
rect 19628 38953 19656 38984
rect 19797 38981 19809 39015
rect 19843 38981 19855 39015
rect 19797 38975 19855 38981
rect 19889 39015 19947 39021
rect 19889 38981 19901 39015
rect 19935 39012 19947 39015
rect 20272 39012 20300 39040
rect 19935 38984 20300 39012
rect 19935 38981 19947 38984
rect 19889 38975 19947 38981
rect 19521 38947 19579 38953
rect 19521 38913 19533 38947
rect 19567 38913 19579 38947
rect 19521 38907 19579 38913
rect 19614 38947 19672 38953
rect 19614 38913 19626 38947
rect 19660 38913 19672 38947
rect 19614 38907 19672 38913
rect 20027 38947 20085 38953
rect 20027 38913 20039 38947
rect 20073 38944 20085 38947
rect 20441 38947 20499 38953
rect 20073 38916 20392 38944
rect 20073 38913 20085 38916
rect 20027 38907 20085 38913
rect 19444 38817 19472 38904
rect 19536 38876 19564 38907
rect 20257 38879 20315 38885
rect 20257 38876 20269 38879
rect 19536 38848 20269 38876
rect 20257 38845 20269 38848
rect 20303 38845 20315 38879
rect 20364 38876 20392 38916
rect 20441 38913 20453 38947
rect 20487 38944 20499 38947
rect 20548 38944 20576 39052
rect 20898 39040 20904 39092
rect 20956 39040 20962 39092
rect 21082 39040 21088 39092
rect 21140 39040 21146 39092
rect 21542 39040 21548 39092
rect 21600 39040 21606 39092
rect 21634 39040 21640 39092
rect 21692 39040 21698 39092
rect 22002 39040 22008 39092
rect 22060 39080 22066 39092
rect 22465 39083 22523 39089
rect 22465 39080 22477 39083
rect 22060 39052 22477 39080
rect 22060 39040 22066 39052
rect 22465 39049 22477 39052
rect 22511 39049 22523 39083
rect 22465 39043 22523 39049
rect 24670 39040 24676 39092
rect 24728 39080 24734 39092
rect 24863 39083 24921 39089
rect 24863 39080 24875 39083
rect 24728 39052 24875 39080
rect 24728 39040 24734 39052
rect 24863 39049 24875 39052
rect 24909 39049 24921 39083
rect 24863 39043 24921 39049
rect 24949 39083 25007 39089
rect 24949 39049 24961 39083
rect 24995 39080 25007 39083
rect 26326 39080 26332 39092
rect 24995 39052 26332 39080
rect 24995 39049 25007 39052
rect 24949 39043 25007 39049
rect 26326 39040 26332 39052
rect 26384 39040 26390 39092
rect 26418 39040 26424 39092
rect 26476 39080 26482 39092
rect 26973 39083 27031 39089
rect 26973 39080 26985 39083
rect 26476 39052 26985 39080
rect 26476 39040 26482 39052
rect 26973 39049 26985 39052
rect 27019 39049 27031 39083
rect 26973 39043 27031 39049
rect 27614 39040 27620 39092
rect 27672 39080 27678 39092
rect 27867 39083 27925 39089
rect 27867 39080 27879 39083
rect 27672 39052 27879 39080
rect 27672 39040 27678 39052
rect 27867 39049 27879 39052
rect 27913 39049 27925 39083
rect 27867 39043 27925 39049
rect 28258 39040 28264 39092
rect 28316 39040 28322 39092
rect 29549 39083 29607 39089
rect 29549 39049 29561 39083
rect 29595 39080 29607 39083
rect 29822 39080 29828 39092
rect 29595 39052 29828 39080
rect 29595 39049 29607 39052
rect 29549 39043 29607 39049
rect 29822 39040 29828 39052
rect 29880 39040 29886 39092
rect 30006 39040 30012 39092
rect 30064 39040 30070 39092
rect 30466 39040 30472 39092
rect 30524 39040 30530 39092
rect 30558 39040 30564 39092
rect 30616 39080 30622 39092
rect 31589 39083 31647 39089
rect 31589 39080 31601 39083
rect 30616 39052 31601 39080
rect 30616 39040 30622 39052
rect 31589 39049 31601 39052
rect 31635 39049 31647 39083
rect 31589 39043 31647 39049
rect 32398 39040 32404 39092
rect 32456 39040 32462 39092
rect 34149 39083 34207 39089
rect 34149 39080 34161 39083
rect 33152 39052 34161 39080
rect 20916 39012 20944 39040
rect 20640 38984 20944 39012
rect 20640 38953 20668 38984
rect 20898 38953 20904 38956
rect 20487 38916 20576 38944
rect 20625 38947 20683 38953
rect 20487 38913 20499 38916
rect 20441 38907 20499 38913
rect 20625 38913 20637 38947
rect 20671 38913 20683 38947
rect 20896 38944 20904 38953
rect 20859 38916 20904 38944
rect 20625 38907 20683 38913
rect 20896 38907 20904 38916
rect 20898 38904 20904 38907
rect 20956 38904 20962 38956
rect 20990 38904 20996 38956
rect 21048 38904 21054 38956
rect 21100 38953 21128 39040
rect 21560 39012 21588 39040
rect 21284 38984 21588 39012
rect 21652 39012 21680 39040
rect 21652 38984 22784 39012
rect 21284 38953 21312 38984
rect 22756 38953 22784 38984
rect 24578 38972 24584 39024
rect 24636 39012 24642 39024
rect 28077 39015 28135 39021
rect 28077 39012 28089 39015
rect 24636 38984 28089 39012
rect 24636 38972 24642 38984
rect 28077 38981 28089 38984
rect 28123 38981 28135 39015
rect 28077 38975 28135 38981
rect 21085 38947 21143 38953
rect 21085 38913 21097 38947
rect 21131 38913 21143 38947
rect 21085 38907 21143 38913
rect 21268 38947 21326 38953
rect 21268 38913 21280 38947
rect 21314 38913 21326 38947
rect 21268 38907 21326 38913
rect 21361 38947 21419 38953
rect 21361 38913 21373 38947
rect 21407 38944 21419 38947
rect 22557 38947 22615 38953
rect 22557 38944 22569 38947
rect 21407 38916 22569 38944
rect 21407 38913 21419 38916
rect 21361 38907 21419 38913
rect 22557 38913 22569 38916
rect 22603 38913 22615 38947
rect 22557 38907 22615 38913
rect 22741 38947 22799 38953
rect 22741 38913 22753 38947
rect 22787 38944 22799 38947
rect 22787 38916 23704 38944
rect 22787 38913 22799 38916
rect 22741 38907 22799 38913
rect 21821 38879 21879 38885
rect 21821 38876 21833 38879
rect 20364 38848 20484 38876
rect 20257 38839 20315 38845
rect 17644 38780 18092 38808
rect 19429 38811 19487 38817
rect 17644 38768 17650 38780
rect 19429 38777 19441 38811
rect 19475 38777 19487 38811
rect 19429 38771 19487 38777
rect 20346 38768 20352 38820
rect 20404 38768 20410 38820
rect 20364 38740 20392 38768
rect 17512 38712 20392 38740
rect 20456 38740 20484 38848
rect 21100 38848 21833 38876
rect 20717 38811 20775 38817
rect 20717 38777 20729 38811
rect 20763 38808 20775 38811
rect 21100 38808 21128 38848
rect 21821 38845 21833 38848
rect 21867 38845 21879 38879
rect 21821 38839 21879 38845
rect 22925 38879 22983 38885
rect 22925 38845 22937 38879
rect 22971 38876 22983 38879
rect 23474 38876 23480 38888
rect 22971 38848 23480 38876
rect 22971 38845 22983 38848
rect 22925 38839 22983 38845
rect 23474 38836 23480 38848
rect 23532 38836 23538 38888
rect 23566 38836 23572 38888
rect 23624 38836 23630 38888
rect 23676 38876 23704 38916
rect 23750 38904 23756 38956
rect 23808 38944 23814 38956
rect 24029 38947 24087 38953
rect 24029 38944 24041 38947
rect 23808 38916 24041 38944
rect 23808 38904 23814 38916
rect 24029 38913 24041 38916
rect 24075 38913 24087 38947
rect 24029 38907 24087 38913
rect 24765 38947 24823 38953
rect 24765 38913 24777 38947
rect 24811 38913 24823 38947
rect 24765 38907 24823 38913
rect 25041 38947 25099 38953
rect 25041 38913 25053 38947
rect 25087 38944 25099 38947
rect 25087 38916 26556 38944
rect 25087 38913 25099 38916
rect 25041 38907 25099 38913
rect 24118 38876 24124 38888
rect 23676 38848 24124 38876
rect 24118 38836 24124 38848
rect 24176 38836 24182 38888
rect 24780 38820 24808 38907
rect 26528 38820 26556 38916
rect 27522 38904 27528 38956
rect 27580 38904 27586 38956
rect 20763 38780 21128 38808
rect 20763 38777 20775 38780
rect 20717 38771 20775 38777
rect 21174 38768 21180 38820
rect 21232 38768 21238 38820
rect 23382 38768 23388 38820
rect 23440 38808 23446 38820
rect 24762 38808 24768 38820
rect 23440 38780 24768 38808
rect 23440 38768 23446 38780
rect 24762 38768 24768 38780
rect 24820 38768 24826 38820
rect 26510 38768 26516 38820
rect 26568 38808 26574 38820
rect 28092 38808 28120 38975
rect 29914 38972 29920 39024
rect 29972 38972 29978 39024
rect 30024 39012 30052 39040
rect 30377 39015 30435 39021
rect 30377 39012 30389 39015
rect 30024 38984 30389 39012
rect 30377 38981 30389 38984
rect 30423 38981 30435 39015
rect 30484 39012 30512 39040
rect 31389 39015 31447 39021
rect 31389 39012 31401 39015
rect 30484 38984 31401 39012
rect 30377 38975 30435 38981
rect 31389 38981 31401 38984
rect 31435 38981 31447 39015
rect 33152 39012 33180 39052
rect 34149 39049 34161 39052
rect 34195 39049 34207 39083
rect 34149 39043 34207 39049
rect 35434 39040 35440 39092
rect 35492 39040 35498 39092
rect 35894 39040 35900 39092
rect 35952 39080 35958 39092
rect 36081 39083 36139 39089
rect 36081 39080 36093 39083
rect 35952 39052 36093 39080
rect 35952 39040 35958 39052
rect 36081 39049 36093 39052
rect 36127 39049 36139 39083
rect 36081 39043 36139 39049
rect 31389 38975 31447 38981
rect 32600 38984 33180 39012
rect 28166 38904 28172 38956
rect 28224 38944 28230 38956
rect 28353 38947 28411 38953
rect 28353 38944 28365 38947
rect 28224 38916 28365 38944
rect 28224 38904 28230 38916
rect 28353 38913 28365 38916
rect 28399 38944 28411 38947
rect 28902 38944 28908 38956
rect 28399 38916 28908 38944
rect 28399 38913 28411 38916
rect 28353 38907 28411 38913
rect 28902 38904 28908 38916
rect 28960 38904 28966 38956
rect 29733 38947 29791 38953
rect 29733 38913 29745 38947
rect 29779 38913 29791 38947
rect 29733 38907 29791 38913
rect 29748 38876 29776 38907
rect 30098 38904 30104 38956
rect 30156 38904 30162 38956
rect 30193 38947 30251 38953
rect 30193 38913 30205 38947
rect 30239 38913 30251 38947
rect 30392 38944 30420 38975
rect 30469 38947 30527 38953
rect 30469 38944 30481 38947
rect 30392 38916 30481 38944
rect 30193 38907 30251 38913
rect 30469 38913 30481 38916
rect 30515 38913 30527 38947
rect 30469 38907 30527 38913
rect 30653 38947 30711 38953
rect 30653 38913 30665 38947
rect 30699 38944 30711 38947
rect 31202 38944 31208 38956
rect 30699 38916 31208 38944
rect 30699 38913 30711 38916
rect 30653 38907 30711 38913
rect 30116 38876 30144 38904
rect 29748 38848 30144 38876
rect 30208 38876 30236 38907
rect 30668 38876 30696 38907
rect 31202 38904 31208 38916
rect 31260 38904 31266 38956
rect 32600 38953 32628 38984
rect 32585 38947 32643 38953
rect 32585 38913 32597 38947
rect 32631 38913 32643 38947
rect 32585 38907 32643 38913
rect 32858 38904 32864 38956
rect 32916 38904 32922 38956
rect 32953 38947 33011 38953
rect 32953 38913 32965 38947
rect 32999 38944 33011 38947
rect 33042 38944 33048 38956
rect 32999 38916 33048 38944
rect 32999 38913 33011 38916
rect 32953 38907 33011 38913
rect 33042 38904 33048 38916
rect 33100 38904 33106 38956
rect 33152 38953 33180 38984
rect 33594 38972 33600 39024
rect 33652 38972 33658 39024
rect 33870 38972 33876 39024
rect 33928 39012 33934 39024
rect 37277 39015 37335 39021
rect 37277 39012 37289 39015
rect 33928 38984 37289 39012
rect 33928 38972 33934 38984
rect 37277 38981 37289 38984
rect 37323 39012 37335 39015
rect 39390 39012 39396 39024
rect 37323 38984 39396 39012
rect 37323 38981 37335 38984
rect 37277 38975 37335 38981
rect 39390 38972 39396 38984
rect 39448 38972 39454 39024
rect 40678 38972 40684 39024
rect 40736 38972 40742 39024
rect 33137 38947 33195 38953
rect 33137 38913 33149 38947
rect 33183 38913 33195 38947
rect 33137 38907 33195 38913
rect 33229 38947 33287 38953
rect 33229 38913 33241 38947
rect 33275 38913 33287 38947
rect 33229 38907 33287 38913
rect 33321 38947 33379 38953
rect 33321 38913 33333 38947
rect 33367 38944 33379 38947
rect 33410 38944 33416 38956
rect 33367 38916 33416 38944
rect 33367 38913 33379 38916
rect 33321 38907 33379 38913
rect 30208 38848 30696 38876
rect 32493 38879 32551 38885
rect 32493 38845 32505 38879
rect 32539 38845 32551 38879
rect 32493 38839 32551 38845
rect 32769 38879 32827 38885
rect 32769 38845 32781 38879
rect 32815 38876 32827 38879
rect 33244 38876 33272 38907
rect 33410 38904 33416 38916
rect 33468 38904 33474 38956
rect 34054 38904 34060 38956
rect 34112 38904 34118 38956
rect 34330 38904 34336 38956
rect 34388 38944 34394 38956
rect 34425 38947 34483 38953
rect 34425 38944 34437 38947
rect 34388 38916 34437 38944
rect 34388 38904 34394 38916
rect 34425 38913 34437 38916
rect 34471 38913 34483 38947
rect 34977 38947 35035 38953
rect 34977 38944 34989 38947
rect 34425 38907 34483 38913
rect 34624 38916 34989 38944
rect 33965 38879 34023 38885
rect 32815 38848 33732 38876
rect 32815 38845 32827 38848
rect 32769 38839 32827 38845
rect 32508 38808 32536 38839
rect 33134 38808 33140 38820
rect 26568 38780 27936 38808
rect 28092 38780 31616 38808
rect 32508 38780 33140 38808
rect 26568 38768 26574 38780
rect 20898 38740 20904 38752
rect 20456 38712 20904 38740
rect 16669 38703 16727 38709
rect 20898 38700 20904 38712
rect 20956 38740 20962 38752
rect 21192 38740 21220 38768
rect 20956 38712 21220 38740
rect 20956 38700 20962 38712
rect 22830 38700 22836 38752
rect 22888 38740 22894 38752
rect 23017 38743 23075 38749
rect 23017 38740 23029 38743
rect 22888 38712 23029 38740
rect 22888 38700 22894 38712
rect 23017 38709 23029 38712
rect 23063 38709 23075 38743
rect 23017 38703 23075 38709
rect 24673 38743 24731 38749
rect 24673 38709 24685 38743
rect 24719 38740 24731 38743
rect 26234 38740 26240 38752
rect 24719 38712 26240 38740
rect 24719 38709 24731 38712
rect 24673 38703 24731 38709
rect 26234 38700 26240 38712
rect 26292 38700 26298 38752
rect 27709 38743 27767 38749
rect 27709 38709 27721 38743
rect 27755 38740 27767 38743
rect 27798 38740 27804 38752
rect 27755 38712 27804 38740
rect 27755 38709 27767 38712
rect 27709 38703 27767 38709
rect 27798 38700 27804 38712
rect 27856 38700 27862 38752
rect 27908 38749 27936 38780
rect 27893 38743 27951 38749
rect 27893 38709 27905 38743
rect 27939 38709 27951 38743
rect 27893 38703 27951 38709
rect 29730 38700 29736 38752
rect 29788 38740 29794 38752
rect 30009 38743 30067 38749
rect 30009 38740 30021 38743
rect 29788 38712 30021 38740
rect 29788 38700 29794 38712
rect 30009 38709 30021 38712
rect 30055 38709 30067 38743
rect 30009 38703 30067 38709
rect 30558 38700 30564 38752
rect 30616 38700 30622 38752
rect 31588 38749 31616 38780
rect 33134 38768 33140 38780
rect 33192 38768 33198 38820
rect 33318 38768 33324 38820
rect 33376 38808 33382 38820
rect 33704 38817 33732 38848
rect 33965 38845 33977 38879
rect 34011 38845 34023 38879
rect 33965 38839 34023 38845
rect 33689 38811 33747 38817
rect 33376 38780 33640 38808
rect 33376 38768 33382 38780
rect 31573 38743 31631 38749
rect 31573 38709 31585 38743
rect 31619 38709 31631 38743
rect 31573 38703 31631 38709
rect 31757 38743 31815 38749
rect 31757 38709 31769 38743
rect 31803 38740 31815 38743
rect 33502 38740 33508 38752
rect 31803 38712 33508 38740
rect 31803 38709 31815 38712
rect 31757 38703 31815 38709
rect 33502 38700 33508 38712
rect 33560 38700 33566 38752
rect 33612 38740 33640 38780
rect 33689 38777 33701 38811
rect 33735 38777 33747 38811
rect 33689 38771 33747 38777
rect 33980 38808 34008 38839
rect 34146 38836 34152 38888
rect 34204 38836 34210 38888
rect 34624 38808 34652 38916
rect 34977 38913 34989 38916
rect 35023 38944 35035 38947
rect 35250 38944 35256 38956
rect 35023 38916 35256 38944
rect 35023 38913 35035 38916
rect 34977 38907 35035 38913
rect 35250 38904 35256 38916
rect 35308 38904 35314 38956
rect 35618 38944 35624 38956
rect 35360 38916 35624 38944
rect 34698 38836 34704 38888
rect 34756 38876 34762 38888
rect 35360 38885 35388 38916
rect 35618 38904 35624 38916
rect 35676 38904 35682 38956
rect 35710 38904 35716 38956
rect 35768 38904 35774 38956
rect 36262 38904 36268 38956
rect 36320 38944 36326 38956
rect 36633 38947 36691 38953
rect 36633 38944 36645 38947
rect 36320 38916 36645 38944
rect 36320 38904 36326 38916
rect 36633 38913 36645 38916
rect 36679 38913 36691 38947
rect 36633 38907 36691 38913
rect 36998 38904 37004 38956
rect 37056 38944 37062 38956
rect 38654 38944 38660 38956
rect 37056 38916 38660 38944
rect 37056 38904 37062 38916
rect 38654 38904 38660 38916
rect 38712 38904 38718 38956
rect 39850 38904 39856 38956
rect 39908 38944 39914 38956
rect 39945 38947 40003 38953
rect 39945 38944 39957 38947
rect 39908 38916 39957 38944
rect 39908 38904 39914 38916
rect 39945 38913 39957 38916
rect 39991 38913 40003 38947
rect 39945 38907 40003 38913
rect 34885 38879 34943 38885
rect 34885 38876 34897 38879
rect 34756 38848 34897 38876
rect 34756 38836 34762 38848
rect 34885 38845 34897 38848
rect 34931 38845 34943 38879
rect 34885 38839 34943 38845
rect 35345 38879 35403 38885
rect 35345 38845 35357 38879
rect 35391 38845 35403 38879
rect 35345 38839 35403 38845
rect 35437 38879 35495 38885
rect 35437 38845 35449 38879
rect 35483 38876 35495 38879
rect 35526 38876 35532 38888
rect 35483 38848 35532 38876
rect 35483 38845 35495 38848
rect 35437 38839 35495 38845
rect 33980 38780 34652 38808
rect 34900 38808 34928 38839
rect 35526 38836 35532 38848
rect 35584 38836 35590 38888
rect 39758 38836 39764 38888
rect 39816 38836 39822 38888
rect 40218 38836 40224 38888
rect 40276 38836 40282 38888
rect 35621 38811 35679 38817
rect 35621 38808 35633 38811
rect 34900 38780 35633 38808
rect 33980 38740 34008 38780
rect 35621 38777 35633 38780
rect 35667 38777 35679 38811
rect 35621 38771 35679 38777
rect 38286 38768 38292 38820
rect 38344 38808 38350 38820
rect 39117 38811 39175 38817
rect 39117 38808 39129 38811
rect 38344 38780 39129 38808
rect 38344 38768 38350 38780
rect 39117 38777 39129 38780
rect 39163 38777 39175 38811
rect 39117 38771 39175 38777
rect 33612 38712 34008 38740
rect 34054 38700 34060 38752
rect 34112 38700 34118 38752
rect 34333 38743 34391 38749
rect 34333 38709 34345 38743
rect 34379 38740 34391 38743
rect 34790 38740 34796 38752
rect 34379 38712 34796 38740
rect 34379 38709 34391 38712
rect 34333 38703 34391 38709
rect 34790 38700 34796 38712
rect 34848 38700 34854 38752
rect 37274 38700 37280 38752
rect 37332 38740 37338 38752
rect 38010 38740 38016 38752
rect 37332 38712 38016 38740
rect 37332 38700 37338 38712
rect 38010 38700 38016 38712
rect 38068 38740 38074 38752
rect 38565 38743 38623 38749
rect 38565 38740 38577 38743
rect 38068 38712 38577 38740
rect 38068 38700 38074 38712
rect 38565 38709 38577 38712
rect 38611 38709 38623 38743
rect 38565 38703 38623 38709
rect 38746 38700 38752 38752
rect 38804 38740 38810 38752
rect 41693 38743 41751 38749
rect 41693 38740 41705 38743
rect 38804 38712 41705 38740
rect 38804 38700 38810 38712
rect 41693 38709 41705 38712
rect 41739 38740 41751 38743
rect 41782 38740 41788 38752
rect 41739 38712 41788 38740
rect 41739 38709 41751 38712
rect 41693 38703 41751 38709
rect 41782 38700 41788 38712
rect 41840 38700 41846 38752
rect 1104 38650 45172 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 45172 38650
rect 1104 38576 45172 38598
rect 2961 38539 3019 38545
rect 2961 38505 2973 38539
rect 3007 38536 3019 38539
rect 3970 38536 3976 38548
rect 3007 38508 3976 38536
rect 3007 38505 3019 38508
rect 2961 38499 3019 38505
rect 3970 38496 3976 38508
rect 4028 38496 4034 38548
rect 5074 38496 5080 38548
rect 5132 38496 5138 38548
rect 8757 38539 8815 38545
rect 8757 38505 8769 38539
rect 8803 38536 8815 38539
rect 9398 38536 9404 38548
rect 8803 38508 9404 38536
rect 8803 38505 8815 38508
rect 8757 38499 8815 38505
rect 9398 38496 9404 38508
rect 9456 38496 9462 38548
rect 17037 38539 17095 38545
rect 17037 38505 17049 38539
rect 17083 38536 17095 38539
rect 17678 38536 17684 38548
rect 17083 38508 17684 38536
rect 17083 38505 17095 38508
rect 17037 38499 17095 38505
rect 17678 38496 17684 38508
rect 17736 38496 17742 38548
rect 18598 38496 18604 38548
rect 18656 38496 18662 38548
rect 23474 38496 23480 38548
rect 23532 38536 23538 38548
rect 24213 38539 24271 38545
rect 24213 38536 24225 38539
rect 23532 38508 24225 38536
rect 23532 38496 23538 38508
rect 24213 38505 24225 38508
rect 24259 38505 24271 38539
rect 24213 38499 24271 38505
rect 4985 38403 5043 38409
rect 4985 38369 4997 38403
rect 5031 38400 5043 38403
rect 5258 38400 5264 38412
rect 5031 38372 5264 38400
rect 5031 38369 5043 38372
rect 4985 38363 5043 38369
rect 5258 38360 5264 38372
rect 5316 38360 5322 38412
rect 7377 38403 7435 38409
rect 7377 38400 7389 38403
rect 6932 38372 7389 38400
rect 6932 38344 6960 38372
rect 7377 38369 7389 38372
rect 7423 38369 7435 38403
rect 7377 38363 7435 38369
rect 9493 38403 9551 38409
rect 9493 38369 9505 38403
rect 9539 38400 9551 38403
rect 10778 38400 10784 38412
rect 9539 38372 10784 38400
rect 9539 38369 9551 38372
rect 9493 38363 9551 38369
rect 10778 38360 10784 38372
rect 10836 38360 10842 38412
rect 15378 38360 15384 38412
rect 15436 38400 15442 38412
rect 15657 38403 15715 38409
rect 15657 38400 15669 38403
rect 15436 38372 15669 38400
rect 15436 38360 15442 38372
rect 15657 38369 15669 38372
rect 15703 38369 15715 38403
rect 15657 38363 15715 38369
rect 17402 38360 17408 38412
rect 17460 38400 17466 38412
rect 18325 38403 18383 38409
rect 18325 38400 18337 38403
rect 17460 38372 18337 38400
rect 17460 38360 17466 38372
rect 18325 38369 18337 38372
rect 18371 38369 18383 38403
rect 19150 38400 19156 38412
rect 18325 38363 18383 38369
rect 18708 38372 19156 38400
rect 1486 38292 1492 38344
rect 1544 38332 1550 38344
rect 1581 38335 1639 38341
rect 1581 38332 1593 38335
rect 1544 38304 1593 38332
rect 1544 38292 1550 38304
rect 1581 38301 1593 38304
rect 1627 38301 1639 38335
rect 1581 38295 1639 38301
rect 6457 38335 6515 38341
rect 6457 38301 6469 38335
rect 6503 38332 6515 38335
rect 6914 38332 6920 38344
rect 6503 38304 6920 38332
rect 6503 38301 6515 38304
rect 6457 38295 6515 38301
rect 6914 38292 6920 38304
rect 6972 38292 6978 38344
rect 7101 38335 7159 38341
rect 7101 38301 7113 38335
rect 7147 38332 7159 38335
rect 8202 38332 8208 38344
rect 7147 38304 8208 38332
rect 7147 38301 7159 38304
rect 7101 38295 7159 38301
rect 8202 38292 8208 38304
rect 8260 38292 8266 38344
rect 9214 38292 9220 38344
rect 9272 38292 9278 38344
rect 17221 38335 17279 38341
rect 17221 38301 17233 38335
rect 17267 38332 17279 38335
rect 17310 38332 17316 38344
rect 17267 38304 17316 38332
rect 17267 38301 17279 38304
rect 17221 38295 17279 38301
rect 17310 38292 17316 38304
rect 17368 38292 17374 38344
rect 18230 38292 18236 38344
rect 18288 38332 18294 38344
rect 18708 38332 18736 38372
rect 19150 38360 19156 38372
rect 19208 38360 19214 38412
rect 22278 38400 22284 38412
rect 22066 38372 22284 38400
rect 18288 38304 18736 38332
rect 18288 38292 18294 38304
rect 18782 38292 18788 38344
rect 18840 38292 18846 38344
rect 19242 38292 19248 38344
rect 19300 38332 19306 38344
rect 19797 38335 19855 38341
rect 19797 38332 19809 38335
rect 19300 38304 19809 38332
rect 19300 38292 19306 38304
rect 19797 38301 19809 38304
rect 19843 38301 19855 38335
rect 19797 38295 19855 38301
rect 21450 38292 21456 38344
rect 21508 38332 21514 38344
rect 22066 38332 22094 38372
rect 22278 38360 22284 38372
rect 22336 38400 22342 38412
rect 22465 38403 22523 38409
rect 22465 38400 22477 38403
rect 22336 38372 22477 38400
rect 22336 38360 22342 38372
rect 22465 38369 22477 38372
rect 22511 38369 22523 38403
rect 22465 38363 22523 38369
rect 22741 38403 22799 38409
rect 22741 38369 22753 38403
rect 22787 38400 22799 38403
rect 22830 38400 22836 38412
rect 22787 38372 22836 38400
rect 22787 38369 22799 38372
rect 22741 38363 22799 38369
rect 22830 38360 22836 38372
rect 22888 38360 22894 38412
rect 24228 38400 24256 38499
rect 30374 38496 30380 38548
rect 30432 38536 30438 38548
rect 31205 38539 31263 38545
rect 31205 38536 31217 38539
rect 30432 38508 31217 38536
rect 30432 38496 30438 38508
rect 31205 38505 31217 38508
rect 31251 38505 31263 38539
rect 31205 38499 31263 38505
rect 33134 38496 33140 38548
rect 33192 38536 33198 38548
rect 33321 38539 33379 38545
rect 33321 38536 33333 38539
rect 33192 38508 33333 38536
rect 33192 38496 33198 38508
rect 33321 38505 33333 38508
rect 33367 38505 33379 38539
rect 33321 38499 33379 38505
rect 33962 38496 33968 38548
rect 34020 38496 34026 38548
rect 34057 38539 34115 38545
rect 34057 38505 34069 38539
rect 34103 38536 34115 38539
rect 34698 38536 34704 38548
rect 34103 38508 34704 38536
rect 34103 38505 34115 38508
rect 34057 38499 34115 38505
rect 34698 38496 34704 38508
rect 34756 38496 34762 38548
rect 35342 38496 35348 38548
rect 35400 38536 35406 38548
rect 35529 38539 35587 38545
rect 35529 38536 35541 38539
rect 35400 38508 35541 38536
rect 35400 38496 35406 38508
rect 35529 38505 35541 38508
rect 35575 38536 35587 38539
rect 35710 38536 35716 38548
rect 35575 38508 35716 38536
rect 35575 38505 35587 38508
rect 35529 38499 35587 38505
rect 35710 38496 35716 38508
rect 35768 38496 35774 38548
rect 35986 38496 35992 38548
rect 36044 38536 36050 38548
rect 36998 38536 37004 38548
rect 36044 38508 37004 38536
rect 36044 38496 36050 38508
rect 36998 38496 37004 38508
rect 37056 38496 37062 38548
rect 39114 38496 39120 38548
rect 39172 38496 39178 38548
rect 40218 38496 40224 38548
rect 40276 38536 40282 38548
rect 40681 38539 40739 38545
rect 40681 38536 40693 38539
rect 40276 38508 40693 38536
rect 40276 38496 40282 38508
rect 40681 38505 40693 38508
rect 40727 38505 40739 38539
rect 40681 38499 40739 38505
rect 33045 38471 33103 38477
rect 33045 38437 33057 38471
rect 33091 38468 33103 38471
rect 33980 38468 34008 38496
rect 39025 38471 39083 38477
rect 33091 38440 34008 38468
rect 34992 38440 35756 38468
rect 33091 38437 33103 38440
rect 33045 38431 33103 38437
rect 24949 38403 25007 38409
rect 24949 38400 24961 38403
rect 24228 38372 24961 38400
rect 24949 38369 24961 38372
rect 24995 38369 25007 38403
rect 25682 38400 25688 38412
rect 24949 38363 25007 38369
rect 25148 38372 25688 38400
rect 21508 38304 22094 38332
rect 21508 38292 21514 38304
rect 1848 38267 1906 38273
rect 1848 38233 1860 38267
rect 1894 38264 1906 38267
rect 2130 38264 2136 38276
rect 1894 38236 2136 38264
rect 1894 38233 1906 38236
rect 1848 38227 1906 38233
rect 2130 38224 2136 38236
rect 2188 38224 2194 38276
rect 6212 38267 6270 38273
rect 6212 38233 6224 38267
rect 6258 38264 6270 38267
rect 7006 38264 7012 38276
rect 6258 38236 7012 38264
rect 6258 38233 6270 38236
rect 6212 38227 6270 38233
rect 7006 38224 7012 38236
rect 7064 38224 7070 38276
rect 7622 38267 7680 38273
rect 7622 38264 7634 38267
rect 7300 38236 7634 38264
rect 4341 38199 4399 38205
rect 4341 38165 4353 38199
rect 4387 38196 4399 38199
rect 4614 38196 4620 38208
rect 4387 38168 4620 38196
rect 4387 38165 4399 38168
rect 4341 38159 4399 38165
rect 4614 38156 4620 38168
rect 4672 38156 4678 38208
rect 7300 38205 7328 38236
rect 7622 38233 7634 38236
rect 7668 38233 7680 38267
rect 9769 38267 9827 38273
rect 9769 38264 9781 38267
rect 7622 38227 7680 38233
rect 9416 38236 9781 38264
rect 9416 38205 9444 38236
rect 9769 38233 9781 38236
rect 9815 38233 9827 38267
rect 9769 38227 9827 38233
rect 10226 38224 10232 38276
rect 10284 38224 10290 38276
rect 15930 38273 15936 38276
rect 15924 38227 15936 38273
rect 15930 38224 15936 38227
rect 15988 38224 15994 38276
rect 25148 38273 25176 38372
rect 25682 38360 25688 38372
rect 25740 38400 25746 38412
rect 26050 38400 26056 38412
rect 25740 38372 26056 38400
rect 25740 38360 25746 38372
rect 26050 38360 26056 38372
rect 26108 38360 26114 38412
rect 32861 38403 32919 38409
rect 29840 38372 30604 38400
rect 25498 38292 25504 38344
rect 25556 38292 25562 38344
rect 29730 38292 29736 38344
rect 29788 38292 29794 38344
rect 29840 38341 29868 38372
rect 30576 38344 30604 38372
rect 32861 38369 32873 38403
rect 32907 38400 32919 38403
rect 33318 38400 33324 38412
rect 32907 38372 33324 38400
rect 32907 38369 32919 38372
rect 32861 38363 32919 38369
rect 33318 38360 33324 38372
rect 33376 38360 33382 38412
rect 34992 38400 35020 38440
rect 33520 38372 35020 38400
rect 35069 38403 35127 38409
rect 33520 38344 33548 38372
rect 35069 38369 35081 38403
rect 35115 38400 35127 38403
rect 35115 38372 35480 38400
rect 35115 38369 35127 38372
rect 35069 38363 35127 38369
rect 29825 38335 29883 38341
rect 29825 38301 29837 38335
rect 29871 38301 29883 38335
rect 29825 38295 29883 38301
rect 30006 38292 30012 38344
rect 30064 38341 30070 38344
rect 30064 38335 30113 38341
rect 30064 38301 30067 38335
rect 30101 38301 30113 38335
rect 30064 38295 30113 38301
rect 30193 38335 30251 38341
rect 30193 38301 30205 38335
rect 30239 38332 30251 38335
rect 30285 38335 30343 38341
rect 30285 38332 30297 38335
rect 30239 38304 30297 38332
rect 30239 38301 30251 38304
rect 30193 38295 30251 38301
rect 30285 38301 30297 38304
rect 30331 38301 30343 38335
rect 30285 38295 30343 38301
rect 30064 38292 30070 38295
rect 30558 38292 30564 38344
rect 30616 38292 30622 38344
rect 30834 38292 30840 38344
rect 30892 38292 30898 38344
rect 30926 38292 30932 38344
rect 30984 38332 30990 38344
rect 31021 38335 31079 38341
rect 31021 38332 31033 38335
rect 30984 38304 31033 38332
rect 30984 38292 30990 38304
rect 31021 38301 31033 38304
rect 31067 38301 31079 38335
rect 31021 38295 31079 38301
rect 32398 38292 32404 38344
rect 32456 38332 32462 38344
rect 32585 38335 32643 38341
rect 32585 38332 32597 38335
rect 32456 38304 32597 38332
rect 32456 38292 32462 38304
rect 32585 38301 32597 38304
rect 32631 38301 32643 38335
rect 32585 38295 32643 38301
rect 32953 38335 33011 38341
rect 32953 38301 32965 38335
rect 32999 38301 33011 38335
rect 32953 38295 33011 38301
rect 25133 38267 25191 38273
rect 25133 38264 25145 38267
rect 18156 38236 19288 38264
rect 23966 38236 25145 38264
rect 18156 38208 18184 38236
rect 7285 38199 7343 38205
rect 7285 38165 7297 38199
rect 7331 38165 7343 38199
rect 7285 38159 7343 38165
rect 9401 38199 9459 38205
rect 9401 38165 9413 38199
rect 9447 38165 9459 38199
rect 9401 38159 9459 38165
rect 11238 38156 11244 38208
rect 11296 38156 11302 38208
rect 17770 38156 17776 38208
rect 17828 38156 17834 38208
rect 18138 38156 18144 38208
rect 18196 38156 18202 38208
rect 19260 38205 19288 38236
rect 25133 38233 25145 38236
rect 25179 38233 25191 38267
rect 25961 38267 26019 38273
rect 25961 38264 25973 38267
rect 25133 38227 25191 38233
rect 25516 38236 25973 38264
rect 25516 38208 25544 38236
rect 25961 38233 25973 38236
rect 26007 38233 26019 38267
rect 25961 38227 26019 38233
rect 29362 38224 29368 38276
rect 29420 38264 29426 38276
rect 29638 38264 29644 38276
rect 29420 38236 29644 38264
rect 29420 38224 29426 38236
rect 29638 38224 29644 38236
rect 29696 38264 29702 38276
rect 29917 38267 29975 38273
rect 29917 38264 29929 38267
rect 29696 38236 29929 38264
rect 29696 38224 29702 38236
rect 29917 38233 29929 38236
rect 29963 38233 29975 38267
rect 32968 38264 32996 38295
rect 33410 38292 33416 38344
rect 33468 38292 33474 38344
rect 33502 38292 33508 38344
rect 33560 38292 33566 38344
rect 33597 38335 33655 38341
rect 33597 38301 33609 38335
rect 33643 38301 33655 38335
rect 33597 38295 33655 38301
rect 33428 38264 33456 38292
rect 33612 38264 33640 38295
rect 33686 38292 33692 38344
rect 33744 38332 33750 38344
rect 33873 38335 33931 38341
rect 33873 38332 33885 38335
rect 33744 38304 33885 38332
rect 33744 38292 33750 38304
rect 33873 38301 33885 38304
rect 33919 38301 33931 38335
rect 33873 38295 33931 38301
rect 34054 38292 34060 38344
rect 34112 38292 34118 38344
rect 34422 38292 34428 38344
rect 34480 38332 34486 38344
rect 34701 38335 34759 38341
rect 34701 38332 34713 38335
rect 34480 38304 34713 38332
rect 34480 38292 34486 38304
rect 34701 38301 34713 38304
rect 34747 38301 34759 38335
rect 34701 38295 34759 38301
rect 34072 38264 34100 38292
rect 32968 38236 33272 38264
rect 33428 38236 33548 38264
rect 33612 38236 34100 38264
rect 34716 38264 34744 38295
rect 34790 38292 34796 38344
rect 34848 38332 34854 38344
rect 34885 38335 34943 38341
rect 34885 38332 34897 38335
rect 34848 38304 34897 38332
rect 34848 38292 34854 38304
rect 34885 38301 34897 38304
rect 34931 38301 34943 38335
rect 35161 38335 35219 38341
rect 35161 38332 35173 38335
rect 34885 38295 34943 38301
rect 35084 38304 35173 38332
rect 35084 38264 35112 38304
rect 35161 38301 35173 38304
rect 35207 38301 35219 38335
rect 35161 38295 35219 38301
rect 35342 38292 35348 38344
rect 35400 38292 35406 38344
rect 35452 38341 35480 38372
rect 35437 38335 35495 38341
rect 35437 38301 35449 38335
rect 35483 38301 35495 38335
rect 35437 38295 35495 38301
rect 35621 38335 35679 38341
rect 35621 38301 35633 38335
rect 35667 38301 35679 38335
rect 35728 38332 35756 38440
rect 39025 38437 39037 38471
rect 39071 38468 39083 38471
rect 39758 38468 39764 38480
rect 39071 38440 39764 38468
rect 39071 38437 39083 38440
rect 39025 38431 39083 38437
rect 39758 38428 39764 38440
rect 39816 38428 39822 38480
rect 39868 38440 40724 38468
rect 38286 38400 38292 38412
rect 36924 38372 38292 38400
rect 36173 38335 36231 38341
rect 36173 38332 36185 38335
rect 35728 38304 36185 38332
rect 35621 38295 35679 38301
rect 36173 38301 36185 38304
rect 36219 38301 36231 38335
rect 36173 38295 36231 38301
rect 34716 38236 35112 38264
rect 35253 38267 35311 38273
rect 29917 38227 29975 38233
rect 33244 38208 33272 38236
rect 33520 38208 33548 38236
rect 35253 38233 35265 38267
rect 35299 38264 35311 38267
rect 35526 38264 35532 38276
rect 35299 38236 35532 38264
rect 35299 38233 35311 38236
rect 35253 38227 35311 38233
rect 35526 38224 35532 38236
rect 35584 38264 35590 38276
rect 35636 38264 35664 38295
rect 36538 38292 36544 38344
rect 36596 38332 36602 38344
rect 36924 38341 36952 38372
rect 38286 38360 38292 38372
rect 38344 38360 38350 38412
rect 39206 38400 39212 38412
rect 38672 38372 39212 38400
rect 36633 38335 36691 38341
rect 36633 38332 36645 38335
rect 36596 38304 36645 38332
rect 36596 38292 36602 38304
rect 36633 38301 36645 38304
rect 36679 38301 36691 38335
rect 36633 38295 36691 38301
rect 36909 38335 36967 38341
rect 36909 38301 36921 38335
rect 36955 38301 36967 38335
rect 36909 38295 36967 38301
rect 36998 38292 37004 38344
rect 37056 38341 37062 38344
rect 37056 38335 37083 38341
rect 37071 38301 37083 38335
rect 37056 38295 37083 38301
rect 37056 38292 37062 38295
rect 37274 38292 37280 38344
rect 37332 38292 37338 38344
rect 38672 38318 38700 38372
rect 39206 38360 39212 38372
rect 39264 38400 39270 38412
rect 39868 38400 39896 38440
rect 40696 38412 40724 38440
rect 39264 38372 39896 38400
rect 39264 38360 39270 38372
rect 40034 38360 40040 38412
rect 40092 38360 40098 38412
rect 40678 38360 40684 38412
rect 40736 38360 40742 38412
rect 39298 38292 39304 38344
rect 39356 38292 39362 38344
rect 39669 38335 39727 38341
rect 39669 38301 39681 38335
rect 39715 38301 39727 38335
rect 39669 38295 39727 38301
rect 35584 38236 35664 38264
rect 35584 38224 35590 38236
rect 36354 38224 36360 38276
rect 36412 38264 36418 38276
rect 36817 38267 36875 38273
rect 36817 38264 36829 38267
rect 36412 38236 36829 38264
rect 36412 38224 36418 38236
rect 36817 38233 36829 38236
rect 36863 38233 36875 38267
rect 37553 38267 37611 38273
rect 37553 38264 37565 38267
rect 36817 38227 36875 38233
rect 37200 38236 37565 38264
rect 19245 38199 19303 38205
rect 19245 38165 19257 38199
rect 19291 38165 19303 38199
rect 19245 38159 19303 38165
rect 24394 38156 24400 38208
rect 24452 38156 24458 38208
rect 25498 38156 25504 38208
rect 25556 38156 25562 38208
rect 26237 38199 26295 38205
rect 26237 38165 26249 38199
rect 26283 38196 26295 38199
rect 26418 38196 26424 38208
rect 26283 38168 26424 38196
rect 26283 38165 26295 38168
rect 26237 38159 26295 38165
rect 26418 38156 26424 38168
rect 26476 38196 26482 38208
rect 27522 38196 27528 38208
rect 26476 38168 27528 38196
rect 26476 38156 26482 38168
rect 27522 38156 27528 38168
rect 27580 38156 27586 38208
rect 29086 38156 29092 38208
rect 29144 38196 29150 38208
rect 29549 38199 29607 38205
rect 29549 38196 29561 38199
rect 29144 38168 29561 38196
rect 29144 38156 29150 38168
rect 29549 38165 29561 38168
rect 29595 38165 29607 38199
rect 29549 38159 29607 38165
rect 32677 38199 32735 38205
rect 32677 38165 32689 38199
rect 32723 38196 32735 38199
rect 32766 38196 32772 38208
rect 32723 38168 32772 38196
rect 32723 38165 32735 38168
rect 32677 38159 32735 38165
rect 32766 38156 32772 38168
rect 32824 38156 32830 38208
rect 33226 38156 33232 38208
rect 33284 38156 33290 38208
rect 33502 38156 33508 38208
rect 33560 38156 33566 38208
rect 34790 38156 34796 38208
rect 34848 38196 34854 38208
rect 35342 38196 35348 38208
rect 34848 38168 35348 38196
rect 34848 38156 34854 38168
rect 35342 38156 35348 38168
rect 35400 38156 35406 38208
rect 36446 38156 36452 38208
rect 36504 38156 36510 38208
rect 37200 38205 37228 38236
rect 37553 38233 37565 38236
rect 37599 38233 37611 38267
rect 37553 38227 37611 38233
rect 39393 38267 39451 38273
rect 39393 38233 39405 38267
rect 39439 38233 39451 38267
rect 39393 38227 39451 38233
rect 39485 38267 39543 38273
rect 39485 38233 39497 38267
rect 39531 38264 39543 38267
rect 39574 38264 39580 38276
rect 39531 38236 39580 38264
rect 39531 38233 39543 38236
rect 39485 38227 39543 38233
rect 37185 38199 37243 38205
rect 37185 38165 37197 38199
rect 37231 38165 37243 38199
rect 37185 38159 37243 38165
rect 38930 38156 38936 38208
rect 38988 38196 38994 38208
rect 39408 38196 39436 38227
rect 39574 38224 39580 38236
rect 39632 38224 39638 38276
rect 39684 38264 39712 38295
rect 40310 38292 40316 38344
rect 40368 38332 40374 38344
rect 40494 38332 40500 38344
rect 40368 38304 40500 38332
rect 40368 38292 40374 38304
rect 40494 38292 40500 38304
rect 40552 38332 40558 38344
rect 40773 38335 40831 38341
rect 40773 38332 40785 38335
rect 40552 38304 40785 38332
rect 40552 38292 40558 38304
rect 40773 38301 40785 38304
rect 40819 38301 40831 38335
rect 40773 38295 40831 38301
rect 42058 38292 42064 38344
rect 42116 38292 42122 38344
rect 40218 38264 40224 38276
rect 39684 38236 40224 38264
rect 40218 38224 40224 38236
rect 40276 38264 40282 38276
rect 41509 38267 41567 38273
rect 41509 38264 41521 38267
rect 40276 38236 41521 38264
rect 40276 38224 40282 38236
rect 41509 38233 41521 38236
rect 41555 38233 41567 38267
rect 41509 38227 41567 38233
rect 41322 38196 41328 38208
rect 38988 38168 41328 38196
rect 38988 38156 38994 38168
rect 41322 38156 41328 38168
rect 41380 38196 41386 38208
rect 41417 38199 41475 38205
rect 41417 38196 41429 38199
rect 41380 38168 41429 38196
rect 41380 38156 41386 38168
rect 41417 38165 41429 38168
rect 41463 38165 41475 38199
rect 41417 38159 41475 38165
rect 1104 38106 45172 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 45172 38106
rect 1104 38032 45172 38054
rect 2130 37952 2136 38004
rect 2188 37952 2194 38004
rect 2498 37952 2504 38004
rect 2556 37952 2562 38004
rect 4433 37995 4491 38001
rect 4433 37961 4445 37995
rect 4479 37992 4491 37995
rect 5258 37992 5264 38004
rect 4479 37964 5264 37992
rect 4479 37961 4491 37964
rect 4433 37955 4491 37961
rect 5258 37952 5264 37964
rect 5316 37952 5322 38004
rect 6730 37952 6736 38004
rect 6788 37952 6794 38004
rect 8573 37995 8631 38001
rect 8573 37961 8585 37995
rect 8619 37992 8631 37995
rect 8938 37992 8944 38004
rect 8619 37964 8944 37992
rect 8619 37961 8631 37964
rect 8573 37955 8631 37961
rect 8938 37952 8944 37964
rect 8996 37952 9002 38004
rect 9030 37952 9036 38004
rect 9088 37952 9094 38004
rect 9122 37952 9128 38004
rect 9180 37952 9186 38004
rect 9214 37952 9220 38004
rect 9272 37992 9278 38004
rect 9585 37995 9643 38001
rect 9585 37992 9597 37995
rect 9272 37964 9597 37992
rect 9272 37952 9278 37964
rect 9585 37961 9597 37964
rect 9631 37961 9643 37995
rect 9585 37955 9643 37961
rect 10042 37952 10048 38004
rect 10100 37952 10106 38004
rect 15194 37992 15200 38004
rect 11992 37964 15200 37992
rect 2317 37859 2375 37865
rect 2317 37825 2329 37859
rect 2363 37856 2375 37859
rect 2516 37856 2544 37952
rect 9140 37924 9168 37952
rect 3068 37896 3648 37924
rect 2363 37828 2544 37856
rect 2363 37825 2375 37828
rect 2317 37819 2375 37825
rect 2774 37816 2780 37868
rect 2832 37816 2838 37868
rect 3068 37865 3096 37896
rect 3620 37868 3648 37896
rect 6656 37896 9168 37924
rect 3053 37859 3111 37865
rect 3053 37856 3065 37859
rect 2976 37828 3065 37856
rect 1486 37748 1492 37800
rect 1544 37788 1550 37800
rect 2976 37788 3004 37828
rect 3053 37825 3065 37828
rect 3099 37825 3111 37859
rect 3309 37859 3367 37865
rect 3309 37856 3321 37859
rect 3053 37819 3111 37825
rect 3160 37828 3321 37856
rect 3160 37788 3188 37828
rect 3309 37825 3321 37828
rect 3355 37825 3367 37859
rect 3309 37819 3367 37825
rect 3602 37816 3608 37868
rect 3660 37816 3666 37868
rect 4890 37865 4896 37868
rect 4884 37819 4896 37865
rect 4890 37816 4896 37819
rect 4948 37816 4954 37868
rect 5442 37816 5448 37868
rect 5500 37856 5506 37868
rect 6656 37856 6684 37896
rect 7466 37865 7472 37868
rect 5500 37828 6684 37856
rect 5500 37816 5506 37828
rect 6564 37797 6592 37828
rect 7460 37819 7472 37865
rect 7466 37816 7472 37819
rect 7524 37816 7530 37868
rect 9140 37856 9168 37896
rect 9953 37927 10011 37933
rect 9953 37893 9965 37927
rect 9999 37924 10011 37927
rect 11238 37924 11244 37936
rect 9999 37896 11244 37924
rect 9999 37893 10011 37896
rect 9953 37887 10011 37893
rect 11238 37884 11244 37896
rect 11296 37884 11302 37936
rect 11992 37865 12020 37964
rect 12253 37927 12311 37933
rect 12253 37893 12265 37927
rect 12299 37924 12311 37927
rect 12526 37924 12532 37936
rect 12299 37896 12532 37924
rect 12299 37893 12311 37896
rect 12253 37887 12311 37893
rect 12526 37884 12532 37896
rect 12584 37884 12590 37936
rect 13924 37865 13952 37964
rect 15194 37952 15200 37964
rect 15252 37952 15258 38004
rect 15657 37995 15715 38001
rect 15657 37961 15669 37995
rect 15703 37992 15715 37995
rect 15838 37992 15844 38004
rect 15703 37964 15844 37992
rect 15703 37961 15715 37964
rect 15657 37955 15715 37961
rect 15838 37952 15844 37964
rect 15896 37952 15902 38004
rect 15930 37952 15936 38004
rect 15988 37952 15994 38004
rect 17313 37995 17371 38001
rect 17313 37961 17325 37995
rect 17359 37992 17371 37995
rect 17954 37992 17960 38004
rect 17359 37964 17960 37992
rect 17359 37961 17371 37964
rect 17313 37955 17371 37961
rect 17954 37952 17960 37964
rect 18012 37952 18018 38004
rect 18785 37995 18843 38001
rect 18785 37961 18797 37995
rect 18831 37992 18843 37995
rect 19242 37992 19248 38004
rect 18831 37964 19248 37992
rect 18831 37961 18843 37964
rect 18785 37955 18843 37961
rect 19242 37952 19248 37964
rect 19300 37952 19306 38004
rect 21177 37995 21235 38001
rect 21177 37961 21189 37995
rect 21223 37992 21235 37995
rect 21450 37992 21456 38004
rect 21223 37964 21456 37992
rect 21223 37961 21235 37964
rect 21177 37955 21235 37961
rect 21450 37952 21456 37964
rect 21508 37952 21514 38004
rect 23201 37995 23259 38001
rect 23201 37961 23213 37995
rect 23247 37992 23259 37995
rect 23566 37992 23572 38004
rect 23247 37964 23572 37992
rect 23247 37961 23259 37964
rect 23201 37955 23259 37961
rect 23566 37952 23572 37964
rect 23624 37952 23630 38004
rect 24394 37952 24400 38004
rect 24452 37952 24458 38004
rect 29086 37992 29092 38004
rect 28460 37964 29092 37992
rect 15470 37884 15476 37936
rect 15528 37924 15534 37936
rect 19705 37927 19763 37933
rect 19705 37924 19717 37927
rect 15528 37896 19717 37924
rect 15528 37884 15534 37896
rect 19705 37893 19717 37896
rect 19751 37924 19763 37927
rect 20806 37924 20812 37936
rect 19751 37896 20812 37924
rect 19751 37893 19763 37896
rect 19705 37887 19763 37893
rect 20806 37884 20812 37896
rect 20864 37884 20870 37936
rect 24412 37924 24440 37952
rect 28460 37933 28488 37964
rect 29086 37952 29092 37964
rect 29144 37952 29150 38004
rect 29917 37995 29975 38001
rect 29917 37961 29929 37995
rect 29963 37961 29975 37995
rect 29917 37955 29975 37961
rect 23768 37896 24440 37924
rect 28445 37927 28503 37933
rect 11977 37859 12035 37865
rect 9140 37828 9260 37856
rect 1544 37760 3004 37788
rect 3068 37760 3188 37788
rect 4617 37791 4675 37797
rect 1544 37748 1550 37760
rect 2961 37723 3019 37729
rect 2961 37689 2973 37723
rect 3007 37720 3019 37723
rect 3068 37720 3096 37760
rect 4617 37757 4629 37791
rect 4663 37757 4675 37791
rect 4617 37751 4675 37757
rect 6549 37791 6607 37797
rect 6549 37757 6561 37791
rect 6595 37757 6607 37791
rect 6549 37751 6607 37757
rect 6641 37791 6699 37797
rect 6641 37757 6653 37791
rect 6687 37788 6699 37791
rect 6822 37788 6828 37800
rect 6687 37760 6828 37788
rect 6687 37757 6699 37760
rect 6641 37751 6699 37757
rect 3007 37692 3096 37720
rect 3007 37689 3019 37692
rect 2961 37683 3019 37689
rect 4632 37652 4660 37751
rect 6822 37748 6828 37760
rect 6880 37748 6886 37800
rect 7193 37791 7251 37797
rect 7193 37757 7205 37791
rect 7239 37757 7251 37791
rect 7193 37751 7251 37757
rect 6914 37720 6920 37732
rect 5552 37692 6920 37720
rect 5552 37652 5580 37692
rect 6196 37664 6224 37692
rect 6914 37680 6920 37692
rect 6972 37720 6978 37732
rect 7208 37720 7236 37751
rect 9122 37748 9128 37800
rect 9180 37748 9186 37800
rect 9232 37797 9260 37828
rect 11977 37825 11989 37859
rect 12023 37825 12035 37859
rect 13909 37859 13967 37865
rect 13386 37828 13860 37856
rect 11977 37819 12035 37825
rect 9217 37791 9275 37797
rect 9217 37757 9229 37791
rect 9263 37757 9275 37791
rect 9217 37751 9275 37757
rect 9398 37748 9404 37800
rect 9456 37788 9462 37800
rect 10229 37791 10287 37797
rect 10229 37788 10241 37791
rect 9456 37760 10241 37788
rect 9456 37748 9462 37760
rect 10229 37757 10241 37760
rect 10275 37788 10287 37791
rect 12802 37788 12808 37800
rect 10275 37760 12808 37788
rect 10275 37757 10287 37760
rect 10229 37751 10287 37757
rect 12802 37748 12808 37760
rect 12860 37748 12866 37800
rect 6972 37692 7236 37720
rect 6972 37680 6978 37692
rect 4632 37624 5580 37652
rect 5994 37612 6000 37664
rect 6052 37612 6058 37664
rect 6178 37612 6184 37664
rect 6236 37612 6242 37664
rect 7098 37612 7104 37664
rect 7156 37612 7162 37664
rect 8662 37612 8668 37664
rect 8720 37612 8726 37664
rect 13354 37612 13360 37664
rect 13412 37652 13418 37664
rect 13725 37655 13783 37661
rect 13725 37652 13737 37655
rect 13412 37624 13737 37652
rect 13412 37612 13418 37624
rect 13725 37621 13737 37624
rect 13771 37621 13783 37655
rect 13832 37652 13860 37828
rect 13909 37825 13921 37859
rect 13955 37825 13967 37859
rect 13909 37819 13967 37825
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 15654 37856 15660 37868
rect 15252 37828 15660 37856
rect 15252 37816 15258 37828
rect 15654 37816 15660 37828
rect 15712 37816 15718 37868
rect 16117 37859 16175 37865
rect 16117 37825 16129 37859
rect 16163 37856 16175 37859
rect 16574 37856 16580 37868
rect 16163 37828 16580 37856
rect 16163 37825 16175 37828
rect 16117 37819 16175 37825
rect 16574 37816 16580 37828
rect 16632 37816 16638 37868
rect 17678 37865 17684 37868
rect 17405 37859 17463 37865
rect 17405 37825 17417 37859
rect 17451 37825 17463 37859
rect 17405 37819 17463 37825
rect 17672 37819 17684 37865
rect 14182 37748 14188 37800
rect 14240 37748 14246 37800
rect 14550 37748 14556 37800
rect 14608 37788 14614 37800
rect 16669 37791 16727 37797
rect 16669 37788 16681 37791
rect 14608 37760 16681 37788
rect 14608 37748 14614 37760
rect 16669 37757 16681 37760
rect 16715 37757 16727 37791
rect 16669 37751 16727 37757
rect 15194 37680 15200 37732
rect 15252 37680 15258 37732
rect 15212 37652 15240 37680
rect 13832 37624 15240 37652
rect 17420 37652 17448 37819
rect 17678 37816 17684 37819
rect 17736 37816 17742 37868
rect 23382 37865 23388 37868
rect 23380 37856 23388 37865
rect 23343 37828 23388 37856
rect 23380 37819 23388 37828
rect 23382 37816 23388 37819
rect 23440 37816 23446 37868
rect 23474 37816 23480 37868
rect 23532 37816 23538 37868
rect 23569 37859 23627 37865
rect 23569 37825 23581 37859
rect 23615 37856 23627 37859
rect 23658 37856 23664 37868
rect 23615 37828 23664 37856
rect 23615 37825 23627 37828
rect 23569 37819 23627 37825
rect 23658 37816 23664 37828
rect 23716 37816 23722 37868
rect 23768 37865 23796 37896
rect 28445 37893 28457 37927
rect 28491 37893 28503 37927
rect 29932 37924 29960 37955
rect 30834 37952 30840 38004
rect 30892 37952 30898 38004
rect 32762 37995 32820 38001
rect 32762 37961 32774 37995
rect 32808 37992 32820 37995
rect 33686 37992 33692 38004
rect 32808 37964 33692 37992
rect 32808 37961 32820 37964
rect 32762 37955 32820 37961
rect 33686 37952 33692 37964
rect 33744 37952 33750 38004
rect 39853 37995 39911 38001
rect 38304 37964 38654 37992
rect 30193 37927 30251 37933
rect 30193 37924 30205 37927
rect 29932 37896 30205 37924
rect 28445 37887 28503 37893
rect 30193 37893 30205 37896
rect 30239 37924 30251 37927
rect 30852 37924 30880 37952
rect 30239 37896 30880 37924
rect 30239 37893 30251 37896
rect 30193 37887 30251 37893
rect 23752 37859 23810 37865
rect 23752 37825 23764 37859
rect 23798 37825 23810 37859
rect 23752 37819 23810 37825
rect 23845 37859 23903 37865
rect 23845 37825 23857 37859
rect 23891 37856 23903 37859
rect 23937 37859 23995 37865
rect 23937 37856 23949 37859
rect 23891 37828 23949 37856
rect 23891 37825 23903 37828
rect 23845 37819 23903 37825
rect 23937 37825 23949 37828
rect 23983 37825 23995 37859
rect 23937 37819 23995 37825
rect 24118 37816 24124 37868
rect 24176 37856 24182 37868
rect 25498 37856 25504 37868
rect 24176 37828 25504 37856
rect 24176 37816 24182 37828
rect 25498 37816 25504 37828
rect 25556 37816 25562 37868
rect 24305 37791 24363 37797
rect 24305 37757 24317 37791
rect 24351 37788 24363 37791
rect 25038 37788 25044 37800
rect 24351 37760 25044 37788
rect 24351 37757 24363 37760
rect 24305 37751 24363 37757
rect 25038 37748 25044 37760
rect 25096 37748 25102 37800
rect 25130 37748 25136 37800
rect 25188 37748 25194 37800
rect 27798 37748 27804 37800
rect 27856 37788 27862 37800
rect 28169 37791 28227 37797
rect 28169 37788 28181 37791
rect 27856 37760 28181 37788
rect 27856 37748 27862 37760
rect 28169 37757 28181 37760
rect 28215 37757 28227 37791
rect 28169 37751 28227 37757
rect 29086 37748 29092 37800
rect 29144 37788 29150 37800
rect 29564 37788 29592 37842
rect 30374 37816 30380 37868
rect 30432 37816 30438 37868
rect 30484 37865 30512 37896
rect 38304 37868 38332 37964
rect 38626 37924 38654 37964
rect 39853 37961 39865 37995
rect 39899 37992 39911 37995
rect 40034 37992 40040 38004
rect 39899 37964 40040 37992
rect 39899 37961 39911 37964
rect 39853 37955 39911 37961
rect 40034 37952 40040 37964
rect 40092 37952 40098 38004
rect 41874 37952 41880 38004
rect 41932 37952 41938 38004
rect 39025 37927 39083 37933
rect 39025 37924 39037 37927
rect 38626 37896 39037 37924
rect 39025 37893 39037 37896
rect 39071 37924 39083 37927
rect 39574 37924 39580 37936
rect 39071 37896 39580 37924
rect 39071 37893 39083 37896
rect 39025 37887 39083 37893
rect 39574 37884 39580 37896
rect 39632 37924 39638 37936
rect 41892 37924 41920 37952
rect 39632 37896 40264 37924
rect 39632 37884 39638 37896
rect 30469 37859 30527 37865
rect 30469 37825 30481 37859
rect 30515 37825 30527 37859
rect 30469 37819 30527 37825
rect 30653 37859 30711 37865
rect 30653 37825 30665 37859
rect 30699 37825 30711 37859
rect 30653 37819 30711 37825
rect 29144 37760 29592 37788
rect 30392 37788 30420 37816
rect 30668 37788 30696 37819
rect 32398 37816 32404 37868
rect 32456 37856 32462 37868
rect 32585 37859 32643 37865
rect 32585 37856 32597 37859
rect 32456 37828 32597 37856
rect 32456 37816 32462 37828
rect 32585 37825 32597 37828
rect 32631 37825 32643 37859
rect 32585 37819 32643 37825
rect 32677 37859 32735 37865
rect 32677 37825 32689 37859
rect 32723 37856 32735 37859
rect 32766 37856 32772 37868
rect 32723 37828 32772 37856
rect 32723 37825 32735 37828
rect 32677 37819 32735 37825
rect 32766 37816 32772 37828
rect 32824 37816 32830 37868
rect 32861 37859 32919 37865
rect 32861 37825 32873 37859
rect 32907 37856 32919 37859
rect 32907 37828 33272 37856
rect 32907 37825 32919 37828
rect 32861 37819 32919 37825
rect 30392 37760 30696 37788
rect 29144 37748 29150 37760
rect 33244 37664 33272 37828
rect 38286 37816 38292 37868
rect 38344 37816 38350 37868
rect 38473 37859 38531 37865
rect 38473 37825 38485 37859
rect 38519 37825 38531 37859
rect 38473 37819 38531 37825
rect 38749 37859 38807 37865
rect 38749 37825 38761 37859
rect 38795 37825 38807 37859
rect 38749 37819 38807 37825
rect 38841 37859 38899 37865
rect 38841 37825 38853 37859
rect 38887 37856 38899 37859
rect 38930 37856 38936 37868
rect 38887 37828 38936 37856
rect 38887 37825 38899 37828
rect 38841 37819 38899 37825
rect 35526 37748 35532 37800
rect 35584 37788 35590 37800
rect 37274 37788 37280 37800
rect 35584 37760 37280 37788
rect 35584 37748 35590 37760
rect 37274 37748 37280 37760
rect 37332 37748 37338 37800
rect 37366 37748 37372 37800
rect 37424 37788 37430 37800
rect 37829 37791 37887 37797
rect 37829 37788 37841 37791
rect 37424 37760 37841 37788
rect 37424 37748 37430 37760
rect 37829 37757 37841 37760
rect 37875 37757 37887 37791
rect 37829 37751 37887 37757
rect 38488 37720 38516 37819
rect 38562 37748 38568 37800
rect 38620 37748 38626 37800
rect 38764 37788 38792 37819
rect 38930 37816 38936 37828
rect 38988 37816 38994 37868
rect 39114 37816 39120 37868
rect 39172 37816 39178 37868
rect 39209 37859 39267 37865
rect 39209 37825 39221 37859
rect 39255 37856 39267 37859
rect 39298 37856 39304 37868
rect 39255 37828 39304 37856
rect 39255 37825 39267 37828
rect 39209 37819 39267 37825
rect 39298 37816 39304 37828
rect 39356 37856 39362 37868
rect 39991 37859 40049 37865
rect 39991 37856 40003 37859
rect 39356 37828 40003 37856
rect 39356 37816 39362 37828
rect 39991 37825 40003 37828
rect 40037 37825 40049 37859
rect 39991 37819 40049 37825
rect 40126 37816 40132 37868
rect 40184 37816 40190 37868
rect 40236 37865 40264 37896
rect 41386 37896 41736 37924
rect 41892 37896 42012 37924
rect 40221 37859 40279 37865
rect 40221 37825 40233 37859
rect 40267 37825 40279 37859
rect 40221 37819 40279 37825
rect 40405 37859 40463 37865
rect 40405 37825 40417 37859
rect 40451 37856 40463 37859
rect 41386 37856 41414 37896
rect 41708 37868 41736 37896
rect 40451 37828 41414 37856
rect 41601 37859 41659 37865
rect 40451 37825 40463 37828
rect 40405 37819 40463 37825
rect 41601 37825 41613 37859
rect 41647 37825 41659 37859
rect 41601 37819 41659 37825
rect 40310 37788 40316 37800
rect 38764 37760 40316 37788
rect 40310 37748 40316 37760
rect 40368 37748 40374 37800
rect 41616 37788 41644 37819
rect 41690 37816 41696 37868
rect 41748 37816 41754 37868
rect 41782 37816 41788 37868
rect 41840 37856 41846 37868
rect 41984 37865 42012 37896
rect 41877 37859 41935 37865
rect 41877 37856 41889 37859
rect 41840 37828 41889 37856
rect 41840 37816 41846 37828
rect 41877 37825 41889 37828
rect 41923 37825 41935 37859
rect 41877 37819 41935 37825
rect 41969 37859 42027 37865
rect 41969 37825 41981 37859
rect 42015 37825 42027 37859
rect 43254 37856 43260 37868
rect 41969 37819 42027 37825
rect 42076 37828 43260 37856
rect 42076 37788 42104 37828
rect 43254 37816 43260 37828
rect 43312 37856 43318 37868
rect 43901 37859 43959 37865
rect 43901 37856 43913 37859
rect 43312 37828 43913 37856
rect 43312 37816 43318 37828
rect 43901 37825 43913 37828
rect 43947 37825 43959 37859
rect 43901 37819 43959 37825
rect 41616 37760 42104 37788
rect 42153 37791 42211 37797
rect 42153 37757 42165 37791
rect 42199 37788 42211 37791
rect 42429 37791 42487 37797
rect 42429 37788 42441 37791
rect 42199 37760 42441 37788
rect 42199 37757 42211 37760
rect 42153 37751 42211 37757
rect 42429 37757 42441 37760
rect 42475 37757 42487 37791
rect 42429 37751 42487 37757
rect 43809 37791 43867 37797
rect 43809 37757 43821 37791
rect 43855 37788 43867 37791
rect 44174 37788 44180 37800
rect 43855 37760 44180 37788
rect 43855 37757 43867 37760
rect 43809 37751 43867 37757
rect 44174 37748 44180 37760
rect 44232 37748 44238 37800
rect 44450 37748 44456 37800
rect 44508 37748 44514 37800
rect 42058 37720 42064 37732
rect 38488 37692 42064 37720
rect 42058 37680 42064 37692
rect 42116 37680 42122 37732
rect 42794 37680 42800 37732
rect 42852 37720 42858 37732
rect 43165 37723 43223 37729
rect 43165 37720 43177 37723
rect 42852 37692 43177 37720
rect 42852 37680 42858 37692
rect 43165 37689 43177 37692
rect 43211 37689 43223 37723
rect 43165 37683 43223 37689
rect 17586 37652 17592 37664
rect 17420 37624 17592 37652
rect 13725 37615 13783 37621
rect 17586 37612 17592 37624
rect 17644 37612 17650 37664
rect 25682 37612 25688 37664
rect 25740 37652 25746 37664
rect 25777 37655 25835 37661
rect 25777 37652 25789 37655
rect 25740 37624 25789 37652
rect 25740 37612 25746 37624
rect 25777 37621 25789 37624
rect 25823 37621 25835 37655
rect 25777 37615 25835 37621
rect 30006 37612 30012 37664
rect 30064 37612 30070 37664
rect 30558 37612 30564 37664
rect 30616 37612 30622 37664
rect 33226 37612 33232 37664
rect 33284 37612 33290 37664
rect 36538 37612 36544 37664
rect 36596 37652 36602 37664
rect 37277 37655 37335 37661
rect 37277 37652 37289 37655
rect 36596 37624 37289 37652
rect 36596 37612 36602 37624
rect 37277 37621 37289 37624
rect 37323 37621 37335 37655
rect 37277 37615 37335 37621
rect 37642 37612 37648 37664
rect 37700 37652 37706 37664
rect 38289 37655 38347 37661
rect 38289 37652 38301 37655
rect 37700 37624 38301 37652
rect 37700 37612 37706 37624
rect 38289 37621 38301 37624
rect 38335 37621 38347 37655
rect 38289 37615 38347 37621
rect 38746 37612 38752 37664
rect 38804 37612 38810 37664
rect 39393 37655 39451 37661
rect 39393 37621 39405 37655
rect 39439 37652 39451 37655
rect 39666 37652 39672 37664
rect 39439 37624 39672 37652
rect 39439 37621 39451 37624
rect 39393 37615 39451 37621
rect 39666 37612 39672 37624
rect 39724 37612 39730 37664
rect 41506 37612 41512 37664
rect 41564 37652 41570 37664
rect 41693 37655 41751 37661
rect 41693 37652 41705 37655
rect 41564 37624 41705 37652
rect 41564 37612 41570 37624
rect 41693 37621 41705 37624
rect 41739 37621 41751 37655
rect 41693 37615 41751 37621
rect 43070 37612 43076 37664
rect 43128 37612 43134 37664
rect 1104 37562 45172 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 45172 37562
rect 1104 37488 45172 37510
rect 2774 37408 2780 37460
rect 2832 37448 2838 37460
rect 3881 37451 3939 37457
rect 3881 37448 3893 37451
rect 2832 37420 3893 37448
rect 2832 37408 2838 37420
rect 3881 37417 3893 37420
rect 3927 37417 3939 37451
rect 3881 37411 3939 37417
rect 4890 37408 4896 37460
rect 4948 37448 4954 37460
rect 5077 37451 5135 37457
rect 5077 37448 5089 37451
rect 4948 37420 5089 37448
rect 4948 37408 4954 37420
rect 5077 37417 5089 37420
rect 5123 37417 5135 37451
rect 6270 37448 6276 37460
rect 5077 37411 5135 37417
rect 5184 37420 6276 37448
rect 5184 37380 5212 37420
rect 6270 37408 6276 37420
rect 6328 37408 6334 37460
rect 6730 37408 6736 37460
rect 6788 37408 6794 37460
rect 6917 37451 6975 37457
rect 6917 37417 6929 37451
rect 6963 37448 6975 37451
rect 7006 37448 7012 37460
rect 6963 37420 7012 37448
rect 6963 37417 6975 37420
rect 6917 37411 6975 37417
rect 7006 37408 7012 37420
rect 7064 37408 7070 37460
rect 7466 37408 7472 37460
rect 7524 37448 7530 37460
rect 7561 37451 7619 37457
rect 7561 37448 7573 37451
rect 7524 37420 7573 37448
rect 7524 37408 7530 37420
rect 7561 37417 7573 37420
rect 7607 37417 7619 37451
rect 7561 37411 7619 37417
rect 12437 37451 12495 37457
rect 12437 37417 12449 37451
rect 12483 37448 12495 37451
rect 12526 37448 12532 37460
rect 12483 37420 12532 37448
rect 12483 37417 12495 37420
rect 12437 37411 12495 37417
rect 12526 37408 12532 37420
rect 12584 37408 12590 37460
rect 17678 37408 17684 37460
rect 17736 37408 17742 37460
rect 18693 37451 18751 37457
rect 18693 37417 18705 37451
rect 18739 37448 18751 37451
rect 18782 37448 18788 37460
rect 18739 37420 18788 37448
rect 18739 37417 18751 37420
rect 18693 37411 18751 37417
rect 18782 37408 18788 37420
rect 18840 37408 18846 37460
rect 20438 37448 20444 37460
rect 19536 37420 20444 37448
rect 6748 37380 6776 37408
rect 3068 37352 5212 37380
rect 5828 37352 6776 37380
rect 2866 37272 2872 37324
rect 2924 37272 2930 37324
rect 3068 37321 3096 37352
rect 3053 37315 3111 37321
rect 3053 37281 3065 37315
rect 3099 37281 3111 37315
rect 3053 37275 3111 37281
rect 4525 37315 4583 37321
rect 4525 37281 4537 37315
rect 4571 37312 4583 37315
rect 4798 37312 4804 37324
rect 4571 37284 4804 37312
rect 4571 37281 4583 37284
rect 4525 37275 4583 37281
rect 4798 37272 4804 37284
rect 4856 37312 4862 37324
rect 5442 37312 5448 37324
rect 4856 37284 5448 37312
rect 4856 37272 4862 37284
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 5828 37321 5856 37352
rect 5813 37315 5871 37321
rect 5813 37281 5825 37315
rect 5859 37281 5871 37315
rect 5813 37275 5871 37281
rect 5902 37272 5908 37324
rect 5960 37272 5966 37324
rect 5994 37272 6000 37324
rect 6052 37312 6058 37324
rect 6733 37315 6791 37321
rect 6733 37312 6745 37315
rect 6052 37284 6745 37312
rect 6052 37272 6058 37284
rect 6733 37281 6745 37284
rect 6779 37281 6791 37315
rect 6733 37275 6791 37281
rect 18141 37315 18199 37321
rect 18141 37281 18153 37315
rect 18187 37312 18199 37315
rect 19536 37312 19564 37420
rect 20438 37408 20444 37420
rect 20496 37408 20502 37460
rect 27522 37408 27528 37460
rect 27580 37448 27586 37460
rect 27580 37420 28488 37448
rect 27580 37408 27586 37420
rect 28460 37380 28488 37420
rect 28902 37408 28908 37460
rect 28960 37408 28966 37460
rect 33226 37408 33232 37460
rect 33284 37408 33290 37460
rect 36354 37448 36360 37460
rect 35636 37420 36360 37448
rect 35636 37380 35664 37420
rect 36354 37408 36360 37420
rect 36412 37448 36418 37460
rect 36814 37448 36820 37460
rect 36412 37420 36820 37448
rect 36412 37408 36418 37420
rect 36814 37408 36820 37420
rect 36872 37448 36878 37460
rect 38286 37448 38292 37460
rect 36872 37420 38292 37448
rect 36872 37408 36878 37420
rect 38286 37408 38292 37420
rect 38344 37408 38350 37460
rect 38749 37451 38807 37457
rect 38749 37448 38761 37451
rect 38396 37420 38761 37448
rect 26988 37352 27292 37380
rect 28460 37352 35664 37380
rect 18187 37284 19564 37312
rect 18187 37281 18199 37284
rect 18141 37275 18199 37281
rect 21450 37272 21456 37324
rect 21508 37272 21514 37324
rect 25593 37315 25651 37321
rect 25593 37281 25605 37315
rect 25639 37312 25651 37315
rect 25682 37312 25688 37324
rect 25639 37284 25688 37312
rect 25639 37281 25651 37284
rect 25593 37275 25651 37281
rect 25682 37272 25688 37284
rect 25740 37272 25746 37324
rect 26050 37272 26056 37324
rect 26108 37312 26114 37324
rect 26988 37312 27016 37352
rect 26108 37284 27016 37312
rect 26108 37272 26114 37284
rect 27062 37272 27068 37324
rect 27120 37272 27126 37324
rect 27264 37312 27292 37352
rect 27264 37284 28580 37312
rect 934 37204 940 37256
rect 992 37244 998 37256
rect 1397 37247 1455 37253
rect 1397 37244 1409 37247
rect 992 37216 1409 37244
rect 992 37204 998 37216
rect 1397 37213 1409 37216
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 2133 37247 2191 37253
rect 2133 37213 2145 37247
rect 2179 37244 2191 37247
rect 4249 37247 4307 37253
rect 2179 37216 2452 37244
rect 2179 37213 2191 37216
rect 2133 37207 2191 37213
rect 1578 37068 1584 37120
rect 1636 37068 1642 37120
rect 1946 37068 1952 37120
rect 2004 37068 2010 37120
rect 2424 37117 2452 37216
rect 4249 37213 4261 37247
rect 4295 37244 4307 37247
rect 4614 37244 4620 37256
rect 4295 37216 4620 37244
rect 4295 37213 4307 37216
rect 4249 37207 4307 37213
rect 4614 37204 4620 37216
rect 4672 37204 4678 37256
rect 5261 37247 5319 37253
rect 5261 37213 5273 37247
rect 5307 37244 5319 37247
rect 5307 37216 5396 37244
rect 5307 37213 5319 37216
rect 5261 37207 5319 37213
rect 2409 37111 2467 37117
rect 2409 37077 2421 37111
rect 2455 37077 2467 37111
rect 2409 37071 2467 37077
rect 2774 37068 2780 37120
rect 2832 37068 2838 37120
rect 4341 37111 4399 37117
rect 4341 37077 4353 37111
rect 4387 37108 4399 37111
rect 4982 37108 4988 37120
rect 4387 37080 4988 37108
rect 4387 37077 4399 37080
rect 4341 37071 4399 37077
rect 4982 37068 4988 37080
rect 5040 37068 5046 37120
rect 5368 37117 5396 37216
rect 7098 37204 7104 37256
rect 7156 37204 7162 37256
rect 7745 37247 7803 37253
rect 7745 37213 7757 37247
rect 7791 37244 7803 37247
rect 8662 37244 8668 37256
rect 7791 37216 8668 37244
rect 7791 37213 7803 37216
rect 7745 37207 7803 37213
rect 8662 37204 8668 37216
rect 8720 37204 8726 37256
rect 12621 37247 12679 37253
rect 12621 37213 12633 37247
rect 12667 37244 12679 37247
rect 12802 37244 12808 37256
rect 12667 37216 12808 37244
rect 12667 37213 12679 37216
rect 12621 37207 12679 37213
rect 12802 37204 12808 37216
rect 12860 37204 12866 37256
rect 15013 37247 15071 37253
rect 15013 37213 15025 37247
rect 15059 37244 15071 37247
rect 15838 37244 15844 37256
rect 15059 37216 15844 37244
rect 15059 37213 15071 37216
rect 15013 37207 15071 37213
rect 15838 37204 15844 37216
rect 15896 37204 15902 37256
rect 17770 37204 17776 37256
rect 17828 37244 17834 37256
rect 17865 37247 17923 37253
rect 17865 37244 17877 37247
rect 17828 37216 17877 37244
rect 17828 37204 17834 37216
rect 17865 37213 17877 37216
rect 17911 37213 17923 37247
rect 17865 37207 17923 37213
rect 18233 37247 18291 37253
rect 18233 37213 18245 37247
rect 18279 37244 18291 37247
rect 18506 37244 18512 37256
rect 18279 37216 18512 37244
rect 18279 37213 18291 37216
rect 18233 37207 18291 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 19242 37204 19248 37256
rect 19300 37204 19306 37256
rect 19521 37247 19579 37253
rect 19521 37213 19533 37247
rect 19567 37244 19579 37247
rect 21468 37244 21496 37272
rect 23474 37244 23480 37256
rect 19567 37216 21496 37244
rect 22848 37216 23480 37244
rect 19567 37213 19579 37216
rect 19521 37207 19579 37213
rect 5721 37179 5779 37185
rect 5721 37145 5733 37179
rect 5767 37176 5779 37179
rect 5902 37176 5908 37188
rect 5767 37148 5908 37176
rect 5767 37145 5779 37148
rect 5721 37139 5779 37145
rect 5902 37136 5908 37148
rect 5960 37176 5966 37188
rect 6181 37179 6239 37185
rect 6181 37176 6193 37179
rect 5960 37148 6193 37176
rect 5960 37136 5966 37148
rect 6181 37145 6193 37148
rect 6227 37145 6239 37179
rect 19766 37179 19824 37185
rect 19766 37176 19778 37179
rect 6181 37139 6239 37145
rect 19444 37148 19778 37176
rect 5353 37111 5411 37117
rect 5353 37077 5365 37111
rect 5399 37077 5411 37111
rect 5353 37071 5411 37077
rect 13722 37068 13728 37120
rect 13780 37108 13786 37120
rect 14921 37111 14979 37117
rect 14921 37108 14933 37111
rect 13780 37080 14933 37108
rect 13780 37068 13786 37080
rect 14921 37077 14933 37080
rect 14967 37077 14979 37111
rect 14921 37071 14979 37077
rect 18230 37068 18236 37120
rect 18288 37108 18294 37120
rect 19444 37117 19472 37148
rect 19766 37145 19778 37148
rect 19812 37145 19824 37179
rect 19766 37139 19824 37145
rect 20806 37136 20812 37188
rect 20864 37176 20870 37188
rect 21698 37179 21756 37185
rect 21698 37176 21710 37179
rect 20864 37148 21710 37176
rect 20864 37136 20870 37148
rect 21698 37145 21710 37148
rect 21744 37145 21756 37179
rect 21698 37139 21756 37145
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18288 37080 18337 37108
rect 18288 37068 18294 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 19429 37111 19487 37117
rect 19429 37077 19441 37111
rect 19475 37077 19487 37111
rect 19429 37071 19487 37077
rect 20901 37111 20959 37117
rect 20901 37077 20913 37111
rect 20947 37108 20959 37111
rect 20990 37108 20996 37120
rect 20947 37080 20996 37108
rect 20947 37077 20959 37080
rect 20901 37071 20959 37077
rect 20990 37068 20996 37080
rect 21048 37108 21054 37120
rect 22278 37108 22284 37120
rect 21048 37080 22284 37108
rect 21048 37068 21054 37080
rect 22278 37068 22284 37080
rect 22336 37068 22342 37120
rect 22462 37068 22468 37120
rect 22520 37108 22526 37120
rect 22848 37117 22876 37216
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 24394 37204 24400 37256
rect 24452 37204 24458 37256
rect 25222 37204 25228 37256
rect 25280 37244 25286 37256
rect 25317 37247 25375 37253
rect 25317 37244 25329 37247
rect 25280 37216 25329 37244
rect 25280 37204 25286 37216
rect 25317 37213 25329 37216
rect 25363 37213 25375 37247
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 25317 37207 25375 37213
rect 26896 37216 27169 37244
rect 22833 37111 22891 37117
rect 22833 37108 22845 37111
rect 22520 37080 22845 37108
rect 22520 37068 22526 37080
rect 22833 37077 22845 37080
rect 22879 37077 22891 37111
rect 22833 37071 22891 37077
rect 22922 37068 22928 37120
rect 22980 37068 22986 37120
rect 24854 37068 24860 37120
rect 24912 37108 24918 37120
rect 25041 37111 25099 37117
rect 25041 37108 25053 37111
rect 24912 37080 25053 37108
rect 24912 37068 24918 37080
rect 25041 37077 25053 37080
rect 25087 37077 25099 37111
rect 25332 37108 25360 37207
rect 26050 37136 26056 37188
rect 26108 37136 26114 37188
rect 26896 37108 26924 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 28552 37244 28580 37284
rect 30558 37272 30564 37324
rect 30616 37272 30622 37324
rect 32861 37315 32919 37321
rect 32861 37312 32873 37315
rect 32416 37284 32873 37312
rect 29825 37247 29883 37253
rect 28552 37230 28994 37244
rect 28566 37216 28994 37230
rect 27157 37207 27215 37213
rect 27430 37136 27436 37188
rect 27488 37136 27494 37188
rect 28966 37176 28994 37216
rect 29825 37213 29837 37247
rect 29871 37213 29883 37247
rect 29825 37207 29883 37213
rect 29840 37176 29868 37207
rect 30006 37204 30012 37256
rect 30064 37204 30070 37256
rect 30576 37176 30604 37272
rect 32416 37256 32444 37284
rect 32861 37281 32873 37284
rect 32907 37281 32919 37315
rect 32861 37275 32919 37281
rect 35526 37272 35532 37324
rect 35584 37272 35590 37324
rect 35805 37315 35863 37321
rect 35805 37281 35817 37315
rect 35851 37312 35863 37315
rect 35894 37312 35900 37324
rect 35851 37284 35900 37312
rect 35851 37281 35863 37284
rect 35805 37275 35863 37281
rect 35894 37272 35900 37284
rect 35952 37272 35958 37324
rect 36446 37272 36452 37324
rect 36504 37312 36510 37324
rect 36998 37312 37004 37324
rect 36504 37284 37004 37312
rect 36504 37272 36510 37284
rect 36998 37272 37004 37284
rect 37056 37312 37062 37324
rect 37056 37284 37412 37312
rect 37056 37272 37062 37284
rect 32398 37204 32404 37256
rect 32456 37204 32462 37256
rect 32766 37204 32772 37256
rect 32824 37204 32830 37256
rect 33045 37247 33103 37253
rect 33045 37213 33057 37247
rect 33091 37244 33103 37247
rect 33134 37244 33140 37256
rect 33091 37216 33140 37244
rect 33091 37213 33103 37216
rect 33045 37207 33103 37213
rect 33134 37204 33140 37216
rect 33192 37204 33198 37256
rect 37384 37244 37412 37284
rect 38010 37244 38016 37256
rect 37384 37216 38016 37244
rect 38010 37204 38016 37216
rect 38068 37204 38074 37256
rect 38105 37247 38163 37253
rect 38105 37213 38117 37247
rect 38151 37244 38163 37247
rect 38396 37244 38424 37420
rect 38749 37417 38761 37420
rect 38795 37448 38807 37451
rect 39114 37448 39120 37460
rect 38795 37420 39120 37448
rect 38795 37417 38807 37420
rect 38749 37411 38807 37417
rect 39114 37408 39120 37420
rect 39172 37408 39178 37460
rect 39298 37408 39304 37460
rect 39356 37408 39362 37460
rect 44177 37451 44235 37457
rect 44177 37417 44189 37451
rect 44223 37448 44235 37451
rect 44450 37448 44456 37460
rect 44223 37420 44456 37448
rect 44223 37417 44235 37420
rect 44177 37411 44235 37417
rect 44450 37408 44456 37420
rect 44508 37408 44514 37460
rect 39316 37380 39344 37408
rect 38626 37352 39344 37380
rect 38151 37216 38424 37244
rect 38473 37247 38531 37253
rect 38151 37213 38163 37216
rect 38105 37207 38163 37213
rect 38473 37213 38485 37247
rect 38519 37244 38531 37247
rect 38626 37244 38654 37352
rect 42705 37315 42763 37321
rect 42705 37281 42717 37315
rect 42751 37312 42763 37315
rect 43070 37312 43076 37324
rect 42751 37284 43076 37312
rect 42751 37281 42763 37284
rect 42705 37275 42763 37281
rect 43070 37272 43076 37284
rect 43128 37272 43134 37324
rect 38519 37216 38654 37244
rect 39301 37247 39359 37253
rect 38519 37213 38531 37216
rect 38473 37207 38531 37213
rect 39301 37213 39313 37247
rect 39347 37213 39359 37247
rect 42426 37244 42432 37256
rect 39301 37207 39359 37213
rect 41892 37216 42432 37244
rect 28966 37148 29132 37176
rect 29840 37148 30604 37176
rect 37030 37148 37504 37176
rect 29104 37120 29132 37148
rect 25332 37080 26924 37108
rect 25041 37071 25099 37077
rect 29086 37068 29092 37120
rect 29144 37068 29150 37120
rect 29914 37068 29920 37120
rect 29972 37068 29978 37120
rect 30282 37068 30288 37120
rect 30340 37108 30346 37120
rect 30834 37108 30840 37120
rect 30340 37080 30840 37108
rect 30340 37068 30346 37080
rect 30834 37068 30840 37080
rect 30892 37068 30898 37120
rect 37274 37068 37280 37120
rect 37332 37068 37338 37120
rect 37476 37108 37504 37148
rect 38286 37136 38292 37188
rect 38344 37136 38350 37188
rect 38378 37136 38384 37188
rect 38436 37136 38442 37188
rect 39206 37176 39212 37188
rect 38488 37148 39212 37176
rect 38488 37108 38516 37148
rect 39206 37136 39212 37148
rect 39264 37136 39270 37188
rect 39316 37176 39344 37207
rect 39316 37148 39528 37176
rect 39500 37120 39528 37148
rect 39574 37136 39580 37188
rect 39632 37176 39638 37188
rect 39942 37176 39948 37188
rect 39632 37148 39948 37176
rect 39632 37136 39638 37148
rect 39942 37136 39948 37148
rect 40000 37176 40006 37188
rect 40589 37179 40647 37185
rect 40589 37176 40601 37179
rect 40000 37148 40601 37176
rect 40000 37136 40006 37148
rect 40589 37145 40601 37148
rect 40635 37145 40647 37179
rect 40589 37139 40647 37145
rect 37476 37080 38516 37108
rect 38654 37068 38660 37120
rect 38712 37068 38718 37120
rect 39482 37068 39488 37120
rect 39540 37068 39546 37120
rect 39850 37068 39856 37120
rect 39908 37108 39914 37120
rect 41892 37117 41920 37216
rect 42426 37204 42432 37216
rect 42484 37204 42490 37256
rect 41877 37111 41935 37117
rect 41877 37108 41889 37111
rect 39908 37080 41889 37108
rect 39908 37068 39914 37080
rect 41877 37077 41889 37080
rect 41923 37077 41935 37111
rect 41877 37071 41935 37077
rect 43714 37068 43720 37120
rect 43772 37108 43778 37120
rect 43824 37108 43852 37230
rect 43772 37080 43852 37108
rect 43772 37068 43778 37080
rect 1104 37018 45172 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 45172 37018
rect 1104 36944 45172 36966
rect 1946 36864 1952 36916
rect 2004 36864 2010 36916
rect 2774 36864 2780 36916
rect 2832 36904 2838 36916
rect 3329 36907 3387 36913
rect 3329 36904 3341 36907
rect 2832 36876 3341 36904
rect 2832 36864 2838 36876
rect 3329 36873 3341 36876
rect 3375 36873 3387 36907
rect 3329 36867 3387 36873
rect 12802 36864 12808 36916
rect 12860 36864 12866 36916
rect 14093 36907 14151 36913
rect 14093 36873 14105 36907
rect 14139 36904 14151 36907
rect 14182 36904 14188 36916
rect 14139 36876 14188 36904
rect 14139 36873 14151 36876
rect 14093 36867 14151 36873
rect 14182 36864 14188 36876
rect 14240 36864 14246 36916
rect 17034 36864 17040 36916
rect 17092 36904 17098 36916
rect 17129 36907 17187 36913
rect 17129 36904 17141 36907
rect 17092 36876 17141 36904
rect 17092 36864 17098 36876
rect 17129 36873 17141 36876
rect 17175 36873 17187 36907
rect 17129 36867 17187 36873
rect 19242 36864 19248 36916
rect 19300 36904 19306 36916
rect 19521 36907 19579 36913
rect 19521 36904 19533 36907
rect 19300 36876 19533 36904
rect 19300 36864 19306 36876
rect 19521 36873 19533 36876
rect 19567 36873 19579 36907
rect 19521 36867 19579 36873
rect 20806 36864 20812 36916
rect 20864 36864 20870 36916
rect 21269 36907 21327 36913
rect 21269 36873 21281 36907
rect 21315 36904 21327 36907
rect 22922 36904 22928 36916
rect 21315 36876 22928 36904
rect 21315 36873 21327 36876
rect 21269 36867 21327 36873
rect 22922 36864 22928 36876
rect 22980 36864 22986 36916
rect 23385 36907 23443 36913
rect 23385 36873 23397 36907
rect 23431 36904 23443 36907
rect 24394 36904 24400 36916
rect 23431 36876 24400 36904
rect 23431 36873 23443 36876
rect 23385 36867 23443 36873
rect 24394 36864 24400 36876
rect 24452 36864 24458 36916
rect 24581 36907 24639 36913
rect 24581 36873 24593 36907
rect 24627 36904 24639 36907
rect 25130 36904 25136 36916
rect 24627 36876 25136 36904
rect 24627 36873 24639 36876
rect 24581 36867 24639 36873
rect 25130 36864 25136 36876
rect 25188 36864 25194 36916
rect 26697 36907 26755 36913
rect 26697 36873 26709 36907
rect 26743 36904 26755 36907
rect 27430 36904 27436 36916
rect 26743 36876 27436 36904
rect 26743 36873 26755 36876
rect 26697 36867 26755 36873
rect 27430 36864 27436 36876
rect 27488 36864 27494 36916
rect 29270 36864 29276 36916
rect 29328 36904 29334 36916
rect 29822 36904 29828 36916
rect 29328 36876 29828 36904
rect 29328 36864 29334 36876
rect 29822 36864 29828 36876
rect 29880 36864 29886 36916
rect 29914 36864 29920 36916
rect 29972 36904 29978 36916
rect 29972 36876 30696 36904
rect 29972 36864 29978 36876
rect 1765 36839 1823 36845
rect 1765 36805 1777 36839
rect 1811 36836 1823 36839
rect 1964 36836 1992 36864
rect 5534 36836 5540 36848
rect 1811 36808 1992 36836
rect 2990 36808 5540 36836
rect 1811 36805 1823 36808
rect 1765 36799 1823 36805
rect 5534 36796 5540 36808
rect 5592 36796 5598 36848
rect 6362 36796 6368 36848
rect 6420 36796 6426 36848
rect 10520 36808 11284 36836
rect 1486 36728 1492 36780
rect 1544 36728 1550 36780
rect 9490 36728 9496 36780
rect 9548 36728 9554 36780
rect 10520 36777 10548 36808
rect 10505 36771 10563 36777
rect 10505 36737 10517 36771
rect 10551 36737 10563 36771
rect 10505 36731 10563 36737
rect 10686 36728 10692 36780
rect 10744 36728 10750 36780
rect 10781 36771 10839 36777
rect 10781 36737 10793 36771
rect 10827 36737 10839 36771
rect 10781 36731 10839 36737
rect 10873 36771 10931 36777
rect 10873 36737 10885 36771
rect 10919 36768 10931 36771
rect 11146 36768 11152 36780
rect 10919 36740 11152 36768
rect 10919 36737 10931 36740
rect 10873 36731 10931 36737
rect 3237 36703 3295 36709
rect 3237 36669 3249 36703
rect 3283 36700 3295 36703
rect 3786 36700 3792 36712
rect 3283 36672 3792 36700
rect 3283 36669 3295 36672
rect 3237 36663 3295 36669
rect 3786 36660 3792 36672
rect 3844 36700 3850 36712
rect 3881 36703 3939 36709
rect 3881 36700 3893 36703
rect 3844 36672 3893 36700
rect 3844 36660 3850 36672
rect 3881 36669 3893 36672
rect 3927 36669 3939 36703
rect 9508 36700 9536 36728
rect 10796 36700 10824 36731
rect 11146 36728 11152 36740
rect 11204 36728 11210 36780
rect 11256 36768 11284 36808
rect 12434 36796 12440 36848
rect 12492 36796 12498 36848
rect 12642 36839 12700 36845
rect 12642 36805 12654 36839
rect 12688 36836 12700 36839
rect 19981 36839 20039 36845
rect 12688 36808 14228 36836
rect 12688 36805 12700 36808
rect 12642 36799 12700 36805
rect 11256 36740 12756 36768
rect 9508 36672 10824 36700
rect 12728 36700 12756 36740
rect 12894 36728 12900 36780
rect 12952 36728 12958 36780
rect 13078 36728 13084 36780
rect 13136 36768 13142 36780
rect 13354 36768 13360 36780
rect 13136 36740 13360 36768
rect 13136 36728 13142 36740
rect 13354 36728 13360 36740
rect 13412 36728 13418 36780
rect 13449 36771 13507 36777
rect 13449 36737 13461 36771
rect 13495 36737 13507 36771
rect 13449 36731 13507 36737
rect 13464 36700 13492 36731
rect 13556 36712 13584 36808
rect 13740 36777 13768 36808
rect 13633 36771 13691 36777
rect 13633 36737 13645 36771
rect 13679 36737 13691 36771
rect 13633 36731 13691 36737
rect 13725 36771 13783 36777
rect 13725 36737 13737 36771
rect 13771 36737 13783 36771
rect 13725 36731 13783 36737
rect 12728 36672 13492 36700
rect 3881 36663 3939 36669
rect 13265 36635 13323 36641
rect 13265 36632 13277 36635
rect 12636 36604 13277 36632
rect 6178 36524 6184 36576
rect 6236 36564 6242 36576
rect 7653 36567 7711 36573
rect 7653 36564 7665 36567
rect 6236 36536 7665 36564
rect 6236 36524 6242 36536
rect 7653 36533 7665 36536
rect 7699 36564 7711 36567
rect 8294 36564 8300 36576
rect 7699 36536 8300 36564
rect 7699 36533 7711 36536
rect 7653 36527 7711 36533
rect 8294 36524 8300 36536
rect 8352 36524 8358 36576
rect 11054 36524 11060 36576
rect 11112 36564 11118 36576
rect 12636 36573 12664 36604
rect 13265 36601 13277 36604
rect 13311 36601 13323 36635
rect 13464 36632 13492 36672
rect 13538 36660 13544 36712
rect 13596 36660 13602 36712
rect 13648 36700 13676 36731
rect 13814 36728 13820 36780
rect 13872 36728 13878 36780
rect 14200 36777 14228 36808
rect 19981 36805 19993 36839
rect 20027 36836 20039 36839
rect 20070 36836 20076 36848
rect 20027 36808 20076 36836
rect 20027 36805 20039 36808
rect 19981 36799 20039 36805
rect 20070 36796 20076 36808
rect 20128 36796 20134 36848
rect 21450 36796 21456 36848
rect 21508 36796 21514 36848
rect 23658 36796 23664 36848
rect 23716 36836 23722 36848
rect 23716 36808 24992 36836
rect 23716 36796 23722 36808
rect 14185 36771 14243 36777
rect 14185 36737 14197 36771
rect 14231 36737 14243 36771
rect 14185 36731 14243 36737
rect 14369 36771 14427 36777
rect 14369 36737 14381 36771
rect 14415 36737 14427 36771
rect 14369 36731 14427 36737
rect 14277 36703 14335 36709
rect 14277 36700 14289 36703
rect 13648 36672 14289 36700
rect 14277 36669 14289 36672
rect 14323 36669 14335 36703
rect 14277 36663 14335 36669
rect 13464 36604 13676 36632
rect 13265 36595 13323 36601
rect 13648 36576 13676 36604
rect 13722 36592 13728 36644
rect 13780 36632 13786 36644
rect 14384 36632 14412 36731
rect 16022 36728 16028 36780
rect 16080 36768 16086 36780
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 16080 36740 17049 36768
rect 16080 36728 16086 36740
rect 17037 36737 17049 36740
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 19889 36771 19947 36777
rect 19889 36737 19901 36771
rect 19935 36768 19947 36771
rect 20346 36768 20352 36780
rect 19935 36740 20352 36768
rect 19935 36737 19947 36740
rect 19889 36731 19947 36737
rect 20346 36728 20352 36740
rect 20404 36728 20410 36780
rect 20625 36771 20683 36777
rect 20625 36737 20637 36771
rect 20671 36768 20683 36771
rect 21468 36768 21496 36796
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 20671 36740 20944 36768
rect 21468 36740 22017 36768
rect 20671 36737 20683 36740
rect 20625 36731 20683 36737
rect 17313 36703 17371 36709
rect 17313 36669 17325 36703
rect 17359 36700 17371 36703
rect 18414 36700 18420 36712
rect 17359 36672 18420 36700
rect 17359 36669 17371 36672
rect 17313 36663 17371 36669
rect 18414 36660 18420 36672
rect 18472 36660 18478 36712
rect 20165 36703 20223 36709
rect 20165 36669 20177 36703
rect 20211 36700 20223 36703
rect 20438 36700 20444 36712
rect 20211 36672 20444 36700
rect 20211 36669 20223 36672
rect 20165 36663 20223 36669
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 13780 36604 14412 36632
rect 13780 36592 13786 36604
rect 11149 36567 11207 36573
rect 11149 36564 11161 36567
rect 11112 36536 11161 36564
rect 11112 36524 11118 36536
rect 11149 36533 11161 36536
rect 11195 36533 11207 36567
rect 11149 36527 11207 36533
rect 12621 36567 12679 36573
rect 12621 36533 12633 36567
rect 12667 36533 12679 36567
rect 12621 36527 12679 36533
rect 13630 36524 13636 36576
rect 13688 36524 13694 36576
rect 16666 36524 16672 36576
rect 16724 36524 16730 36576
rect 20456 36564 20484 36660
rect 20916 36641 20944 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22272 36771 22330 36777
rect 22272 36737 22284 36771
rect 22318 36768 22330 36771
rect 23014 36768 23020 36780
rect 22318 36740 23020 36768
rect 22318 36737 22330 36740
rect 22272 36731 22330 36737
rect 23014 36728 23020 36740
rect 23072 36728 23078 36780
rect 24762 36777 24768 36780
rect 24760 36731 24768 36777
rect 24762 36728 24768 36731
rect 24820 36728 24826 36780
rect 24854 36728 24860 36780
rect 24912 36728 24918 36780
rect 24964 36777 24992 36808
rect 25038 36796 25044 36848
rect 25096 36836 25102 36848
rect 27062 36836 27068 36848
rect 25096 36808 27068 36836
rect 25096 36796 25102 36808
rect 25148 36777 25176 36808
rect 27062 36796 27068 36808
rect 27120 36796 27126 36848
rect 27157 36839 27215 36845
rect 27157 36805 27169 36839
rect 27203 36836 27215 36839
rect 27982 36836 27988 36848
rect 27203 36808 27988 36836
rect 27203 36805 27215 36808
rect 27157 36799 27215 36805
rect 27982 36796 27988 36808
rect 28040 36796 28046 36848
rect 30469 36839 30527 36845
rect 30469 36836 30481 36839
rect 29196 36808 30481 36836
rect 24949 36771 25007 36777
rect 24949 36737 24961 36771
rect 24995 36737 25007 36771
rect 24949 36731 25007 36737
rect 25132 36771 25190 36777
rect 25132 36737 25144 36771
rect 25178 36737 25190 36771
rect 25132 36731 25190 36737
rect 25225 36771 25283 36777
rect 25225 36737 25237 36771
rect 25271 36768 25283 36771
rect 25317 36771 25375 36777
rect 25317 36768 25329 36771
rect 25271 36740 25329 36768
rect 25271 36737 25283 36740
rect 25225 36731 25283 36737
rect 25317 36737 25329 36740
rect 25363 36737 25375 36771
rect 25317 36731 25375 36737
rect 21358 36660 21364 36712
rect 21416 36660 21422 36712
rect 21453 36703 21511 36709
rect 21453 36669 21465 36703
rect 21499 36669 21511 36703
rect 21453 36663 21511 36669
rect 20901 36635 20959 36641
rect 20901 36601 20913 36635
rect 20947 36601 20959 36635
rect 21468 36632 21496 36663
rect 20901 36595 20959 36601
rect 21376 36604 21496 36632
rect 24964 36632 24992 36731
rect 25498 36728 25504 36780
rect 25556 36728 25562 36780
rect 26789 36771 26847 36777
rect 26789 36737 26801 36771
rect 26835 36768 26847 36771
rect 27338 36768 27344 36780
rect 26835 36740 27344 36768
rect 26835 36737 26847 36740
rect 26789 36731 26847 36737
rect 27338 36728 27344 36740
rect 27396 36728 27402 36780
rect 29196 36777 29224 36808
rect 30469 36805 30481 36808
rect 30515 36805 30527 36839
rect 30469 36799 30527 36805
rect 30668 36836 30696 36876
rect 30834 36864 30840 36916
rect 30892 36904 30898 36916
rect 31018 36904 31024 36916
rect 30892 36876 31024 36904
rect 30892 36864 30898 36876
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 31665 36907 31723 36913
rect 31665 36873 31677 36907
rect 31711 36904 31723 36907
rect 31711 36876 35480 36904
rect 31711 36873 31723 36876
rect 31665 36867 31723 36873
rect 31297 36839 31355 36845
rect 31297 36836 31309 36839
rect 30668 36808 31309 36836
rect 29181 36771 29239 36777
rect 29181 36737 29193 36771
rect 29227 36737 29239 36771
rect 29181 36731 29239 36737
rect 29270 36728 29276 36780
rect 29328 36728 29334 36780
rect 29362 36728 29368 36780
rect 29420 36728 29426 36780
rect 29503 36771 29561 36777
rect 29503 36737 29515 36771
rect 29549 36768 29561 36771
rect 30098 36768 30104 36780
rect 29549 36740 30104 36768
rect 29549 36737 29561 36740
rect 29503 36731 29561 36737
rect 25685 36703 25743 36709
rect 25685 36669 25697 36703
rect 25731 36700 25743 36703
rect 26142 36700 26148 36712
rect 25731 36672 26148 36700
rect 25731 36669 25743 36672
rect 25685 36663 25743 36669
rect 26142 36660 26148 36672
rect 26200 36660 26206 36712
rect 29518 36700 29546 36731
rect 30098 36728 30104 36740
rect 30156 36768 30162 36780
rect 30374 36768 30380 36780
rect 30156 36740 30380 36768
rect 30156 36728 30162 36740
rect 30374 36728 30380 36740
rect 30432 36728 30438 36780
rect 30668 36777 30696 36808
rect 31297 36805 31309 36808
rect 31343 36836 31355 36839
rect 33137 36839 33195 36845
rect 31343 36808 31524 36836
rect 31343 36805 31355 36808
rect 31297 36799 31355 36805
rect 30653 36771 30711 36777
rect 30653 36737 30665 36771
rect 30699 36737 30711 36771
rect 30653 36731 30711 36737
rect 30742 36728 30748 36780
rect 30800 36768 30806 36780
rect 30929 36771 30987 36777
rect 30800 36766 30880 36768
rect 30929 36766 30941 36771
rect 30800 36740 30941 36766
rect 30800 36728 30806 36740
rect 30852 36738 30941 36740
rect 30929 36737 30941 36738
rect 30975 36737 30987 36771
rect 30929 36731 30987 36737
rect 31018 36728 31024 36780
rect 31076 36728 31082 36780
rect 31496 36777 31524 36808
rect 33137 36805 33149 36839
rect 33183 36805 33195 36839
rect 34149 36839 34207 36845
rect 34149 36836 34161 36839
rect 33137 36799 33195 36805
rect 33796 36808 34161 36836
rect 31113 36771 31171 36777
rect 31113 36737 31125 36771
rect 31159 36768 31171 36771
rect 31389 36771 31447 36777
rect 31389 36768 31401 36771
rect 31159 36740 31401 36768
rect 31159 36737 31171 36740
rect 31113 36731 31171 36737
rect 31389 36737 31401 36740
rect 31435 36737 31447 36771
rect 31389 36731 31447 36737
rect 31481 36771 31539 36777
rect 31481 36737 31493 36771
rect 31527 36737 31539 36771
rect 31481 36731 31539 36737
rect 32585 36771 32643 36777
rect 32585 36737 32597 36771
rect 32631 36768 32643 36771
rect 32766 36768 32772 36780
rect 32631 36740 32772 36768
rect 32631 36737 32643 36740
rect 32585 36731 32643 36737
rect 29380 36692 29546 36700
rect 29196 36672 29546 36692
rect 29641 36703 29699 36709
rect 29196 36664 29408 36672
rect 29641 36669 29653 36703
rect 29687 36700 29699 36703
rect 29733 36703 29791 36709
rect 29733 36700 29745 36703
rect 29687 36672 29745 36700
rect 29687 36669 29699 36672
rect 29196 36632 29224 36664
rect 29641 36663 29699 36669
rect 29733 36669 29745 36672
rect 29779 36669 29791 36703
rect 29733 36663 29791 36669
rect 29914 36660 29920 36712
rect 29972 36700 29978 36712
rect 30285 36703 30343 36709
rect 30285 36700 30297 36703
rect 29972 36672 30297 36700
rect 29972 36660 29978 36672
rect 30285 36669 30297 36672
rect 30331 36669 30343 36703
rect 30760 36700 30788 36728
rect 31128 36700 31156 36731
rect 32766 36728 32772 36740
rect 32824 36768 32830 36780
rect 33152 36768 33180 36799
rect 33796 36780 33824 36808
rect 34149 36805 34161 36808
rect 34195 36805 34207 36839
rect 34149 36799 34207 36805
rect 34241 36839 34299 36845
rect 34241 36805 34253 36839
rect 34287 36836 34299 36839
rect 34606 36836 34612 36848
rect 34287 36808 34612 36836
rect 34287 36805 34299 36808
rect 34241 36799 34299 36805
rect 32824 36740 33180 36768
rect 33229 36771 33287 36777
rect 32824 36728 32830 36740
rect 33229 36737 33241 36771
rect 33275 36737 33287 36771
rect 33229 36731 33287 36737
rect 30760 36672 31156 36700
rect 30285 36663 30343 36669
rect 31662 36660 31668 36712
rect 31720 36660 31726 36712
rect 32398 36660 32404 36712
rect 32456 36700 32462 36712
rect 32493 36703 32551 36709
rect 32493 36700 32505 36703
rect 32456 36672 32505 36700
rect 32456 36660 32462 36672
rect 32493 36669 32505 36672
rect 32539 36669 32551 36703
rect 33244 36700 33272 36731
rect 33778 36728 33784 36780
rect 33836 36728 33842 36780
rect 33962 36728 33968 36780
rect 34020 36728 34026 36780
rect 32493 36663 32551 36669
rect 32876 36672 33272 36700
rect 34164 36700 34192 36799
rect 34606 36796 34612 36808
rect 34664 36796 34670 36848
rect 34330 36728 34336 36780
rect 34388 36728 34394 36780
rect 35452 36777 35480 36876
rect 35894 36864 35900 36916
rect 35952 36904 35958 36916
rect 35989 36907 36047 36913
rect 35989 36904 36001 36907
rect 35952 36876 36001 36904
rect 35952 36864 35958 36876
rect 35989 36873 36001 36876
rect 36035 36873 36047 36907
rect 35989 36867 36047 36873
rect 37737 36907 37795 36913
rect 37737 36873 37749 36907
rect 37783 36904 37795 36907
rect 37783 36876 37872 36904
rect 37783 36873 37795 36876
rect 37737 36867 37795 36873
rect 35713 36839 35771 36845
rect 35713 36805 35725 36839
rect 35759 36836 35771 36839
rect 36538 36836 36544 36848
rect 35759 36808 36544 36836
rect 35759 36805 35771 36808
rect 35713 36799 35771 36805
rect 36538 36796 36544 36808
rect 36596 36796 36602 36848
rect 37277 36839 37335 36845
rect 37277 36805 37289 36839
rect 37323 36836 37335 36839
rect 37642 36836 37648 36848
rect 37323 36808 37648 36836
rect 37323 36805 37335 36808
rect 37277 36799 37335 36805
rect 37642 36796 37648 36808
rect 37700 36796 37706 36848
rect 35437 36771 35495 36777
rect 35437 36737 35449 36771
rect 35483 36737 35495 36771
rect 35437 36731 35495 36737
rect 35621 36771 35679 36777
rect 35621 36737 35633 36771
rect 35667 36737 35679 36771
rect 35621 36731 35679 36737
rect 35805 36771 35863 36777
rect 35805 36737 35817 36771
rect 35851 36768 35863 36771
rect 35986 36768 35992 36780
rect 35851 36740 35992 36768
rect 35851 36737 35863 36740
rect 35805 36731 35863 36737
rect 35636 36700 35664 36731
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 36170 36728 36176 36780
rect 36228 36728 36234 36780
rect 37844 36777 37872 36876
rect 38010 36864 38016 36916
rect 38068 36864 38074 36916
rect 38289 36907 38347 36913
rect 38289 36873 38301 36907
rect 38335 36904 38347 36907
rect 38470 36904 38476 36916
rect 38335 36876 38476 36904
rect 38335 36873 38347 36876
rect 38289 36867 38347 36873
rect 38470 36864 38476 36876
rect 38528 36904 38534 36916
rect 38528 36876 39528 36904
rect 38528 36864 38534 36876
rect 38028 36777 38056 36864
rect 39500 36848 39528 36876
rect 39850 36864 39856 36916
rect 39908 36864 39914 36916
rect 44174 36864 44180 36916
rect 44232 36864 44238 36916
rect 39206 36796 39212 36848
rect 39264 36796 39270 36848
rect 39482 36796 39488 36848
rect 39540 36796 39546 36848
rect 39666 36796 39672 36848
rect 39724 36836 39730 36848
rect 39761 36839 39819 36845
rect 39761 36836 39773 36839
rect 39724 36808 39773 36836
rect 39724 36796 39730 36808
rect 39761 36805 39773 36808
rect 39807 36805 39819 36839
rect 39868 36836 39896 36864
rect 42794 36836 42800 36848
rect 39868 36808 40080 36836
rect 39761 36799 39819 36805
rect 40052 36777 40080 36808
rect 42260 36808 42800 36836
rect 37553 36771 37611 36777
rect 36648 36740 37504 36768
rect 35710 36700 35716 36712
rect 34164 36672 35716 36700
rect 32876 36644 32904 36672
rect 35710 36660 35716 36672
rect 35768 36660 35774 36712
rect 36449 36703 36507 36709
rect 36449 36700 36461 36703
rect 36188 36672 36461 36700
rect 24964 36604 29224 36632
rect 21376 36564 21404 36604
rect 29822 36592 29828 36644
rect 29880 36632 29886 36644
rect 31021 36635 31079 36641
rect 31021 36632 31033 36635
rect 29880 36604 31033 36632
rect 29880 36592 29886 36604
rect 31021 36601 31033 36604
rect 31067 36601 31079 36635
rect 31021 36595 31079 36601
rect 32858 36592 32864 36644
rect 32916 36592 32922 36644
rect 32953 36635 33011 36641
rect 32953 36601 32965 36635
rect 32999 36632 33011 36635
rect 33410 36632 33416 36644
rect 32999 36604 33416 36632
rect 32999 36601 33011 36604
rect 32953 36595 33011 36601
rect 33410 36592 33416 36604
rect 33468 36592 33474 36644
rect 36188 36576 36216 36672
rect 36449 36669 36461 36672
rect 36495 36669 36507 36703
rect 36449 36663 36507 36669
rect 21542 36564 21548 36576
rect 20456 36536 21548 36564
rect 21542 36524 21548 36536
rect 21600 36524 21606 36576
rect 27798 36524 27804 36576
rect 27856 36564 27862 36576
rect 28445 36567 28503 36573
rect 28445 36564 28457 36567
rect 27856 36536 28457 36564
rect 27856 36524 27862 36536
rect 28445 36533 28457 36536
rect 28491 36533 28503 36567
rect 28445 36527 28503 36533
rect 28994 36524 29000 36576
rect 29052 36524 29058 36576
rect 29730 36524 29736 36576
rect 29788 36564 29794 36576
rect 30282 36564 30288 36576
rect 29788 36536 30288 36564
rect 29788 36524 29794 36536
rect 30282 36524 30288 36536
rect 30340 36524 30346 36576
rect 30374 36524 30380 36576
rect 30432 36564 30438 36576
rect 33042 36564 33048 36576
rect 30432 36536 33048 36564
rect 30432 36524 30438 36536
rect 33042 36524 33048 36536
rect 33100 36524 33106 36576
rect 34514 36524 34520 36576
rect 34572 36524 34578 36576
rect 36170 36524 36176 36576
rect 36228 36524 36234 36576
rect 36541 36567 36599 36573
rect 36541 36533 36553 36567
rect 36587 36564 36599 36567
rect 36648 36564 36676 36740
rect 37369 36703 37427 36709
rect 37369 36669 37381 36703
rect 37415 36669 37427 36703
rect 37369 36663 37427 36669
rect 36725 36635 36783 36641
rect 36725 36601 36737 36635
rect 36771 36632 36783 36635
rect 37384 36632 37412 36663
rect 36771 36604 37412 36632
rect 37476 36632 37504 36740
rect 37553 36737 37565 36771
rect 37599 36737 37611 36771
rect 37553 36731 37611 36737
rect 37829 36771 37887 36777
rect 37829 36737 37841 36771
rect 37875 36737 37887 36771
rect 37829 36731 37887 36737
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 40037 36771 40095 36777
rect 40037 36737 40049 36771
rect 40083 36737 40095 36771
rect 40037 36731 40095 36737
rect 41233 36771 41291 36777
rect 41233 36737 41245 36771
rect 41279 36737 41291 36771
rect 41233 36731 41291 36737
rect 37568 36700 37596 36731
rect 39758 36700 39764 36712
rect 37568 36672 39764 36700
rect 39758 36660 39764 36672
rect 39816 36660 39822 36712
rect 40957 36703 41015 36709
rect 40957 36669 40969 36703
rect 41003 36700 41015 36703
rect 41049 36703 41107 36709
rect 41049 36700 41061 36703
rect 41003 36672 41061 36700
rect 41003 36669 41015 36672
rect 40957 36663 41015 36669
rect 41049 36669 41061 36672
rect 41095 36669 41107 36703
rect 41248 36700 41276 36731
rect 41322 36728 41328 36780
rect 41380 36728 41386 36780
rect 41414 36728 41420 36780
rect 41472 36728 41478 36780
rect 41598 36728 41604 36780
rect 41656 36728 41662 36780
rect 41874 36728 41880 36780
rect 41932 36728 41938 36780
rect 41969 36771 42027 36777
rect 41969 36737 41981 36771
rect 42015 36768 42027 36771
rect 42058 36768 42064 36780
rect 42015 36740 42064 36768
rect 42015 36737 42027 36740
rect 41969 36731 42027 36737
rect 42058 36728 42064 36740
rect 42116 36728 42122 36780
rect 42260 36777 42288 36808
rect 42794 36796 42800 36808
rect 42852 36796 42858 36848
rect 43714 36796 43720 36848
rect 43772 36796 43778 36848
rect 42245 36771 42303 36777
rect 42245 36737 42257 36771
rect 42291 36737 42303 36771
rect 42245 36731 42303 36737
rect 42426 36728 42432 36780
rect 42484 36728 42490 36780
rect 41432 36700 41460 36728
rect 41892 36700 41920 36728
rect 41248 36672 41920 36700
rect 41049 36663 41107 36669
rect 42702 36660 42708 36712
rect 42760 36660 42766 36712
rect 42153 36635 42211 36641
rect 42153 36632 42165 36635
rect 37476 36604 37780 36632
rect 36771 36601 36783 36604
rect 36725 36595 36783 36601
rect 37752 36576 37780 36604
rect 39960 36604 41368 36632
rect 36587 36536 36676 36564
rect 36587 36533 36599 36536
rect 36541 36527 36599 36533
rect 37274 36524 37280 36576
rect 37332 36524 37338 36576
rect 37734 36524 37740 36576
rect 37792 36524 37798 36576
rect 37921 36567 37979 36573
rect 37921 36533 37933 36567
rect 37967 36564 37979 36567
rect 38286 36564 38292 36576
rect 37967 36536 38292 36564
rect 37967 36533 37979 36536
rect 37921 36527 37979 36533
rect 38286 36524 38292 36536
rect 38344 36564 38350 36576
rect 39960 36564 39988 36604
rect 41340 36576 41368 36604
rect 41524 36604 42165 36632
rect 41524 36576 41552 36604
rect 42153 36601 42165 36604
rect 42199 36601 42211 36635
rect 42153 36595 42211 36601
rect 38344 36536 39988 36564
rect 38344 36524 38350 36536
rect 40310 36524 40316 36576
rect 40368 36524 40374 36576
rect 41322 36524 41328 36576
rect 41380 36524 41386 36576
rect 41506 36524 41512 36576
rect 41564 36524 41570 36576
rect 41690 36524 41696 36576
rect 41748 36524 41754 36576
rect 1104 36474 45172 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 45172 36474
rect 1104 36400 45172 36422
rect 3786 36320 3792 36372
rect 3844 36320 3850 36372
rect 10505 36363 10563 36369
rect 10505 36329 10517 36363
rect 10551 36360 10563 36363
rect 10686 36360 10692 36372
rect 10551 36332 10692 36360
rect 10551 36329 10563 36332
rect 10505 36323 10563 36329
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 11974 36320 11980 36372
rect 12032 36360 12038 36372
rect 12437 36363 12495 36369
rect 12437 36360 12449 36363
rect 12032 36332 12449 36360
rect 12032 36320 12038 36332
rect 12437 36329 12449 36332
rect 12483 36329 12495 36363
rect 13722 36360 13728 36372
rect 12437 36323 12495 36329
rect 13372 36332 13728 36360
rect 3804 36165 3832 36320
rect 9766 36292 9772 36304
rect 8864 36264 9772 36292
rect 7006 36184 7012 36236
rect 7064 36224 7070 36236
rect 7742 36224 7748 36236
rect 7064 36196 7748 36224
rect 7064 36184 7070 36196
rect 7742 36184 7748 36196
rect 7800 36224 7806 36236
rect 8864 36224 8892 36264
rect 9766 36252 9772 36264
rect 9824 36252 9830 36304
rect 7800 36196 8892 36224
rect 7800 36184 7806 36196
rect 8938 36184 8944 36236
rect 8996 36224 9002 36236
rect 10689 36227 10747 36233
rect 10689 36224 10701 36227
rect 8996 36196 10701 36224
rect 8996 36184 9002 36196
rect 10689 36193 10701 36196
rect 10735 36193 10747 36227
rect 10689 36187 10747 36193
rect 10965 36227 11023 36233
rect 10965 36193 10977 36227
rect 11011 36224 11023 36227
rect 11054 36224 11060 36236
rect 11011 36196 11060 36224
rect 11011 36193 11023 36196
rect 10965 36187 11023 36193
rect 11054 36184 11060 36196
rect 11112 36184 11118 36236
rect 12894 36224 12900 36236
rect 12636 36196 12900 36224
rect 3789 36159 3847 36165
rect 3789 36125 3801 36159
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 5350 36116 5356 36168
rect 5408 36116 5414 36168
rect 6178 36116 6184 36168
rect 6236 36156 6242 36168
rect 6273 36159 6331 36165
rect 6273 36156 6285 36159
rect 6236 36128 6285 36156
rect 6236 36116 6242 36128
rect 6273 36125 6285 36128
rect 6319 36125 6331 36159
rect 9401 36159 9459 36165
rect 9401 36156 9413 36159
rect 6273 36119 6331 36125
rect 8956 36128 9413 36156
rect 6546 36048 6552 36100
rect 6604 36048 6610 36100
rect 7006 36088 7012 36100
rect 6840 36060 7012 36088
rect 3881 36023 3939 36029
rect 3881 35989 3893 36023
rect 3927 36020 3939 36023
rect 4062 36020 4068 36032
rect 3927 35992 4068 36020
rect 3927 35989 3939 35992
rect 3881 35983 3939 35989
rect 4062 35980 4068 35992
rect 4120 35980 4126 36032
rect 5074 35980 5080 36032
rect 5132 36020 5138 36032
rect 5169 36023 5227 36029
rect 5169 36020 5181 36023
rect 5132 35992 5181 36020
rect 5132 35980 5138 35992
rect 5169 35989 5181 35992
rect 5215 35989 5227 36023
rect 5169 35983 5227 35989
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 6840 36020 6868 36060
rect 7006 36048 7012 36060
rect 7064 36048 7070 36100
rect 8386 36048 8392 36100
rect 8444 36088 8450 36100
rect 8956 36097 8984 36128
rect 9401 36125 9413 36128
rect 9447 36125 9459 36159
rect 9582 36156 9588 36168
rect 9401 36119 9459 36125
rect 9508 36128 9588 36156
rect 8941 36091 8999 36097
rect 8941 36088 8953 36091
rect 8444 36060 8953 36088
rect 8444 36048 8450 36060
rect 8941 36057 8953 36060
rect 8987 36057 8999 36091
rect 8941 36051 8999 36057
rect 9125 36091 9183 36097
rect 9125 36057 9137 36091
rect 9171 36088 9183 36091
rect 9508 36088 9536 36128
rect 9582 36116 9588 36128
rect 9640 36116 9646 36168
rect 9858 36116 9864 36168
rect 9916 36116 9922 36168
rect 12636 36165 12664 36196
rect 12894 36184 12900 36196
rect 12952 36184 12958 36236
rect 10413 36159 10471 36165
rect 10413 36125 10425 36159
rect 10459 36125 10471 36159
rect 10413 36119 10471 36125
rect 10597 36159 10655 36165
rect 10597 36125 10609 36159
rect 10643 36125 10655 36159
rect 10597 36119 10655 36125
rect 12621 36159 12679 36165
rect 12621 36125 12633 36159
rect 12667 36125 12679 36159
rect 12621 36119 12679 36125
rect 10428 36088 10456 36119
rect 9171 36060 9536 36088
rect 9600 36060 10456 36088
rect 10612 36088 10640 36119
rect 12802 36116 12808 36168
rect 12860 36116 12866 36168
rect 12986 36116 12992 36168
rect 13044 36156 13050 36168
rect 13372 36165 13400 36332
rect 13722 36320 13728 36332
rect 13780 36320 13786 36372
rect 14185 36363 14243 36369
rect 14185 36329 14197 36363
rect 14231 36360 14243 36363
rect 14550 36360 14556 36372
rect 14231 36332 14556 36360
rect 14231 36329 14243 36332
rect 14185 36323 14243 36329
rect 14550 36320 14556 36332
rect 14608 36320 14614 36372
rect 16022 36320 16028 36372
rect 16080 36320 16086 36372
rect 20438 36320 20444 36372
rect 20496 36360 20502 36372
rect 22281 36363 22339 36369
rect 22281 36360 22293 36363
rect 20496 36332 22293 36360
rect 20496 36320 20502 36332
rect 22281 36329 22293 36332
rect 22327 36329 22339 36363
rect 22281 36323 22339 36329
rect 23014 36320 23020 36372
rect 23072 36320 23078 36372
rect 27696 36363 27754 36369
rect 27696 36329 27708 36363
rect 27742 36360 27754 36363
rect 28994 36360 29000 36372
rect 27742 36332 29000 36360
rect 27742 36329 27754 36332
rect 27696 36323 27754 36329
rect 28994 36320 29000 36332
rect 29052 36320 29058 36372
rect 30193 36363 30251 36369
rect 30193 36329 30205 36363
rect 30239 36360 30251 36363
rect 31662 36360 31668 36372
rect 30239 36332 31668 36360
rect 30239 36329 30251 36332
rect 30193 36323 30251 36329
rect 31662 36320 31668 36332
rect 31720 36320 31726 36372
rect 32493 36363 32551 36369
rect 32493 36329 32505 36363
rect 32539 36360 32551 36363
rect 32858 36360 32864 36372
rect 32539 36332 32864 36360
rect 32539 36329 32551 36332
rect 32493 36323 32551 36329
rect 32858 36320 32864 36332
rect 32916 36320 32922 36372
rect 34514 36320 34520 36372
rect 34572 36320 34578 36372
rect 35526 36320 35532 36372
rect 35584 36360 35590 36372
rect 39206 36360 39212 36372
rect 35584 36332 36492 36360
rect 35584 36320 35590 36332
rect 13541 36295 13599 36301
rect 13541 36261 13553 36295
rect 13587 36292 13599 36295
rect 13814 36292 13820 36304
rect 13587 36264 13820 36292
rect 13587 36261 13599 36264
rect 13541 36255 13599 36261
rect 13814 36252 13820 36264
rect 13872 36252 13878 36304
rect 21542 36252 21548 36304
rect 21600 36292 21606 36304
rect 22189 36295 22247 36301
rect 21600 36264 21680 36292
rect 21600 36252 21606 36264
rect 13630 36184 13636 36236
rect 13688 36184 13694 36236
rect 15933 36227 15991 36233
rect 15933 36193 15945 36227
rect 15979 36224 15991 36227
rect 16758 36224 16764 36236
rect 15979 36196 16764 36224
rect 15979 36193 15991 36196
rect 15933 36187 15991 36193
rect 16758 36184 16764 36196
rect 16816 36184 16822 36236
rect 16942 36184 16948 36236
rect 17000 36224 17006 36236
rect 17497 36227 17555 36233
rect 17497 36224 17509 36227
rect 17000 36196 17509 36224
rect 17000 36184 17006 36196
rect 17497 36193 17509 36196
rect 17543 36193 17555 36227
rect 17497 36187 17555 36193
rect 17770 36184 17776 36236
rect 17828 36224 17834 36236
rect 17828 36196 19564 36224
rect 17828 36184 17834 36196
rect 13357 36159 13415 36165
rect 13357 36156 13369 36159
rect 13044 36128 13369 36156
rect 13044 36116 13050 36128
rect 13357 36125 13369 36128
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 13538 36116 13544 36168
rect 13596 36116 13602 36168
rect 13906 36116 13912 36168
rect 13964 36116 13970 36168
rect 18046 36116 18052 36168
rect 18104 36116 18110 36168
rect 19245 36159 19303 36165
rect 19245 36125 19257 36159
rect 19291 36156 19303 36159
rect 19426 36156 19432 36168
rect 19291 36128 19432 36156
rect 19291 36125 19303 36128
rect 19245 36119 19303 36125
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 19536 36165 19564 36196
rect 21450 36184 21456 36236
rect 21508 36184 21514 36236
rect 21652 36233 21680 36264
rect 22189 36261 22201 36295
rect 22235 36292 22247 36295
rect 27249 36295 27307 36301
rect 22235 36264 23244 36292
rect 22235 36261 22247 36264
rect 22189 36255 22247 36261
rect 21637 36227 21695 36233
rect 21637 36193 21649 36227
rect 21683 36193 21695 36227
rect 21637 36187 21695 36193
rect 22278 36184 22284 36236
rect 22336 36224 22342 36236
rect 22833 36227 22891 36233
rect 22833 36224 22845 36227
rect 22336 36196 22845 36224
rect 22336 36184 22342 36196
rect 22833 36193 22845 36196
rect 22879 36193 22891 36227
rect 22833 36187 22891 36193
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36156 19579 36159
rect 21468 36156 21496 36184
rect 23216 36165 23244 36264
rect 27249 36261 27261 36295
rect 27295 36292 27307 36295
rect 27338 36292 27344 36304
rect 27295 36264 27344 36292
rect 27295 36261 27307 36264
rect 27249 36255 27307 36261
rect 27338 36252 27344 36264
rect 27396 36252 27402 36304
rect 29178 36252 29184 36304
rect 29236 36292 29242 36304
rect 29914 36292 29920 36304
rect 29236 36264 29920 36292
rect 29236 36252 29242 36264
rect 29914 36252 29920 36264
rect 29972 36252 29978 36304
rect 32876 36292 32904 36320
rect 32876 36264 33916 36292
rect 23290 36184 23296 36236
rect 23348 36224 23354 36236
rect 24949 36227 25007 36233
rect 24949 36224 24961 36227
rect 23348 36196 24961 36224
rect 23348 36184 23354 36196
rect 24949 36193 24961 36196
rect 24995 36193 25007 36227
rect 24949 36187 25007 36193
rect 25222 36184 25228 36236
rect 25280 36224 25286 36236
rect 27433 36227 27491 36233
rect 27433 36224 27445 36227
rect 25280 36196 27445 36224
rect 25280 36184 25286 36196
rect 27433 36193 27445 36196
rect 27479 36224 27491 36227
rect 27798 36224 27804 36236
rect 27479 36196 27804 36224
rect 27479 36193 27491 36196
rect 27433 36187 27491 36193
rect 27798 36184 27804 36196
rect 27856 36224 27862 36236
rect 33888 36233 33916 36264
rect 30745 36227 30803 36233
rect 30745 36224 30757 36227
rect 27856 36196 30757 36224
rect 27856 36184 27862 36196
rect 30745 36193 30757 36196
rect 30791 36193 30803 36227
rect 30745 36187 30803 36193
rect 31021 36227 31079 36233
rect 31021 36193 31033 36227
rect 31067 36224 31079 36227
rect 32585 36227 32643 36233
rect 32585 36224 32597 36227
rect 31067 36196 32597 36224
rect 31067 36193 31079 36196
rect 31021 36187 31079 36193
rect 32585 36193 32597 36196
rect 32631 36193 32643 36227
rect 33873 36227 33931 36233
rect 32585 36187 32643 36193
rect 32692 36196 32996 36224
rect 32692 36168 32720 36196
rect 19567 36128 21496 36156
rect 23201 36159 23259 36165
rect 19567 36125 19579 36128
rect 19521 36119 19579 36125
rect 23201 36125 23213 36159
rect 23247 36125 23259 36159
rect 24854 36156 24860 36168
rect 23201 36119 23259 36125
rect 24136 36128 24860 36156
rect 11054 36088 11060 36100
rect 10612 36060 11060 36088
rect 9171 36057 9183 36060
rect 9125 36051 9183 36057
rect 5592 35992 6868 36020
rect 5592 35980 5598 35992
rect 6914 35980 6920 36032
rect 6972 36020 6978 36032
rect 7834 36020 7840 36032
rect 6972 35992 7840 36020
rect 6972 35980 6978 35992
rect 7834 35980 7840 35992
rect 7892 36020 7898 36032
rect 8021 36023 8079 36029
rect 8021 36020 8033 36023
rect 7892 35992 8033 36020
rect 7892 35980 7898 35992
rect 8021 35989 8033 35992
rect 8067 35989 8079 36023
rect 8021 35983 8079 35989
rect 9306 35980 9312 36032
rect 9364 35980 9370 36032
rect 9490 35980 9496 36032
rect 9548 36020 9554 36032
rect 9600 36020 9628 36060
rect 11054 36048 11060 36060
rect 11112 36048 11118 36100
rect 12713 36091 12771 36097
rect 11348 36060 11454 36088
rect 9548 35992 9628 36020
rect 9548 35980 9554 35992
rect 9674 35980 9680 36032
rect 9732 35980 9738 36032
rect 9766 35980 9772 36032
rect 9824 36020 9830 36032
rect 10226 36020 10232 36032
rect 9824 35992 10232 36020
rect 9824 35980 9830 35992
rect 10226 35980 10232 35992
rect 10284 36020 10290 36032
rect 11348 36020 11376 36060
rect 12713 36057 12725 36091
rect 12759 36088 12771 36091
rect 13556 36088 13584 36116
rect 12759 36060 13584 36088
rect 12759 36057 12771 36060
rect 12713 36051 12771 36057
rect 15194 36048 15200 36100
rect 15252 36088 15258 36100
rect 15252 36060 15608 36088
rect 15252 36048 15258 36060
rect 10284 35992 11376 36020
rect 10284 35980 10290 35992
rect 12802 35980 12808 36032
rect 12860 36020 12866 36032
rect 13078 36020 13084 36032
rect 12860 35992 13084 36020
rect 12860 35980 12866 35992
rect 13078 35980 13084 35992
rect 13136 35980 13142 36032
rect 13633 36023 13691 36029
rect 13633 35989 13645 36023
rect 13679 36020 13691 36023
rect 13998 36020 14004 36032
rect 13679 35992 14004 36020
rect 13679 35989 13691 35992
rect 13633 35983 13691 35989
rect 13998 35980 14004 35992
rect 14056 35980 14062 36032
rect 15580 36020 15608 36060
rect 15654 36048 15660 36100
rect 15712 36048 15718 36100
rect 17954 36088 17960 36100
rect 17066 36060 17960 36088
rect 17144 36020 17172 36060
rect 17954 36048 17960 36060
rect 18012 36048 18018 36100
rect 19766 36091 19824 36097
rect 19766 36088 19778 36091
rect 19444 36060 19778 36088
rect 15580 35992 17172 36020
rect 17862 35980 17868 36032
rect 17920 35980 17926 36032
rect 19444 36029 19472 36060
rect 19766 36057 19778 36060
rect 19812 36057 19824 36091
rect 19766 36051 19824 36057
rect 21821 36091 21879 36097
rect 21821 36057 21833 36091
rect 21867 36088 21879 36091
rect 24136 36088 24164 36128
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 25774 36116 25780 36168
rect 25832 36116 25838 36168
rect 26326 36116 26332 36168
rect 26384 36156 26390 36168
rect 26973 36159 27031 36165
rect 26973 36156 26985 36159
rect 26384 36128 26985 36156
rect 26384 36116 26390 36128
rect 26973 36125 26985 36128
rect 27019 36125 27031 36159
rect 26973 36119 27031 36125
rect 29549 36159 29607 36165
rect 29549 36125 29561 36159
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 25225 36091 25283 36097
rect 25225 36088 25237 36091
rect 21867 36060 24164 36088
rect 24780 36060 25237 36088
rect 21867 36057 21879 36060
rect 21821 36051 21879 36057
rect 24780 36032 24808 36060
rect 25225 36057 25237 36060
rect 25271 36057 25283 36091
rect 26988 36088 27016 36119
rect 27614 36088 27620 36100
rect 26988 36060 27620 36088
rect 25225 36051 25283 36057
rect 27614 36048 27620 36060
rect 27672 36048 27678 36100
rect 29086 36088 29092 36100
rect 28934 36060 29092 36088
rect 29086 36048 29092 36060
rect 29144 36088 29150 36100
rect 29564 36088 29592 36119
rect 29730 36116 29736 36168
rect 29788 36116 29794 36168
rect 29822 36116 29828 36168
rect 29880 36116 29886 36168
rect 30006 36116 30012 36168
rect 30064 36116 30070 36168
rect 30558 36116 30564 36168
rect 30616 36116 30622 36168
rect 32674 36116 32680 36168
rect 32732 36116 32738 36168
rect 32766 36116 32772 36168
rect 32824 36116 32830 36168
rect 32968 36165 32996 36196
rect 33873 36193 33885 36227
rect 33919 36193 33931 36227
rect 34532 36224 34560 36320
rect 36464 36233 36492 36332
rect 36556 36332 39212 36360
rect 36173 36227 36231 36233
rect 36173 36224 36185 36227
rect 34532 36196 36185 36224
rect 33873 36187 33931 36193
rect 36173 36193 36185 36196
rect 36219 36193 36231 36227
rect 36173 36187 36231 36193
rect 36449 36227 36507 36233
rect 36449 36193 36461 36227
rect 36495 36193 36507 36227
rect 36449 36187 36507 36193
rect 32953 36159 33011 36165
rect 32953 36125 32965 36159
rect 32999 36125 33011 36159
rect 32953 36119 33011 36125
rect 33042 36116 33048 36168
rect 33100 36165 33106 36168
rect 33100 36159 33129 36165
rect 33117 36125 33129 36159
rect 33100 36119 33129 36125
rect 33229 36159 33287 36165
rect 33229 36125 33241 36159
rect 33275 36156 33287 36159
rect 33321 36159 33379 36165
rect 33321 36156 33333 36159
rect 33275 36128 33333 36156
rect 33275 36125 33287 36128
rect 33229 36119 33287 36125
rect 33321 36125 33333 36128
rect 33367 36125 33379 36159
rect 33321 36119 33379 36125
rect 33100 36116 33106 36119
rect 30576 36088 30604 36116
rect 29144 36060 29316 36088
rect 29564 36060 30604 36088
rect 30668 36060 31510 36088
rect 29144 36048 29150 36060
rect 19429 36023 19487 36029
rect 19429 35989 19441 36023
rect 19475 35989 19487 36023
rect 19429 35983 19487 35989
rect 20898 35980 20904 36032
rect 20956 35980 20962 36032
rect 21450 35980 21456 36032
rect 21508 36020 21514 36032
rect 21729 36023 21787 36029
rect 21729 36020 21741 36023
rect 21508 35992 21741 36020
rect 21508 35980 21514 35992
rect 21729 35989 21741 35992
rect 21775 35989 21787 36023
rect 21729 35983 21787 35989
rect 24394 35980 24400 36032
rect 24452 35980 24458 36032
rect 24762 35980 24768 36032
rect 24820 35980 24826 36032
rect 29178 35980 29184 36032
rect 29236 35980 29242 36032
rect 29288 36020 29316 36060
rect 30668 36020 30696 36060
rect 32858 36048 32864 36100
rect 32916 36048 32922 36100
rect 35710 36048 35716 36100
rect 35768 36088 35774 36100
rect 36556 36088 36584 36332
rect 39206 36320 39212 36332
rect 39264 36320 39270 36372
rect 40208 36363 40266 36369
rect 40208 36329 40220 36363
rect 40254 36360 40266 36363
rect 40310 36360 40316 36372
rect 40254 36332 40316 36360
rect 40254 36329 40266 36332
rect 40208 36323 40266 36329
rect 40310 36320 40316 36332
rect 40368 36320 40374 36372
rect 41690 36320 41696 36372
rect 41748 36320 41754 36372
rect 42702 36320 42708 36372
rect 42760 36360 42766 36372
rect 42797 36363 42855 36369
rect 42797 36360 42809 36363
rect 42760 36332 42809 36360
rect 42760 36320 42766 36332
rect 42797 36329 42809 36332
rect 42843 36329 42855 36363
rect 42797 36323 42855 36329
rect 43714 36320 43720 36372
rect 43772 36320 43778 36372
rect 38746 36184 38752 36236
rect 38804 36224 38810 36236
rect 39209 36227 39267 36233
rect 39209 36224 39221 36227
rect 38804 36196 39221 36224
rect 38804 36184 38810 36196
rect 39209 36193 39221 36196
rect 39255 36193 39267 36227
rect 39209 36187 39267 36193
rect 39485 36227 39543 36233
rect 39485 36193 39497 36227
rect 39531 36224 39543 36227
rect 39850 36224 39856 36236
rect 39531 36196 39856 36224
rect 39531 36193 39543 36196
rect 39485 36187 39543 36193
rect 39850 36184 39856 36196
rect 39908 36224 39914 36236
rect 39945 36227 40003 36233
rect 39945 36224 39957 36227
rect 39908 36196 39957 36224
rect 39908 36184 39914 36196
rect 39945 36193 39957 36196
rect 39991 36224 40003 36227
rect 40218 36224 40224 36236
rect 39991 36196 40224 36224
rect 39991 36193 40003 36196
rect 39945 36187 40003 36193
rect 40218 36184 40224 36196
rect 40276 36184 40282 36236
rect 41708 36224 41736 36320
rect 42153 36227 42211 36233
rect 42153 36224 42165 36227
rect 41708 36196 42165 36224
rect 42153 36193 42165 36196
rect 42199 36193 42211 36227
rect 42153 36187 42211 36193
rect 43732 36156 43760 36320
rect 41354 36142 43760 36156
rect 41340 36128 43760 36142
rect 35768 36060 36584 36088
rect 35768 36048 35774 36060
rect 37182 36048 37188 36100
rect 37240 36088 37246 36100
rect 39206 36088 39212 36100
rect 37240 36060 37872 36088
rect 38778 36060 39212 36088
rect 37240 36048 37246 36060
rect 29288 35992 30696 36020
rect 34698 35980 34704 36032
rect 34756 35980 34762 36032
rect 37734 35980 37740 36032
rect 37792 35980 37798 36032
rect 37844 36020 37872 36060
rect 39206 36048 39212 36060
rect 39264 36048 39270 36100
rect 41340 36020 41368 36128
rect 37844 35992 41368 36020
rect 41598 35980 41604 36032
rect 41656 36020 41662 36032
rect 41693 36023 41751 36029
rect 41693 36020 41705 36023
rect 41656 35992 41705 36020
rect 41656 35980 41662 35992
rect 41693 35989 41705 35992
rect 41739 36020 41751 36023
rect 42058 36020 42064 36032
rect 41739 35992 42064 36020
rect 41739 35989 41751 35992
rect 41693 35983 41751 35989
rect 42058 35980 42064 35992
rect 42116 35980 42122 36032
rect 1104 35930 45172 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 45172 35930
rect 1104 35856 45172 35878
rect 4433 35819 4491 35825
rect 4433 35785 4445 35819
rect 4479 35816 4491 35819
rect 4706 35816 4712 35828
rect 4479 35788 4712 35816
rect 4479 35785 4491 35788
rect 4433 35779 4491 35785
rect 4706 35776 4712 35788
rect 4764 35816 4770 35828
rect 4764 35788 5120 35816
rect 4764 35776 4770 35788
rect 3326 35689 3332 35692
rect 3320 35643 3332 35689
rect 3326 35640 3332 35643
rect 3384 35640 3390 35692
rect 5092 35689 5120 35788
rect 5350 35776 5356 35828
rect 5408 35816 5414 35828
rect 5445 35819 5503 35825
rect 5445 35816 5457 35819
rect 5408 35788 5457 35816
rect 5408 35776 5414 35788
rect 5445 35785 5457 35788
rect 5491 35785 5503 35819
rect 5445 35779 5503 35785
rect 5902 35776 5908 35828
rect 5960 35776 5966 35828
rect 5994 35776 6000 35828
rect 6052 35816 6058 35828
rect 6270 35816 6276 35828
rect 6052 35788 6276 35816
rect 6052 35776 6058 35788
rect 6270 35776 6276 35788
rect 6328 35816 6334 35828
rect 9398 35816 9404 35828
rect 6328 35788 9404 35816
rect 6328 35776 6334 35788
rect 9398 35776 9404 35788
rect 9456 35776 9462 35828
rect 11241 35819 11299 35825
rect 9508 35788 11192 35816
rect 9508 35760 9536 35788
rect 6457 35751 6515 35757
rect 6457 35748 6469 35751
rect 5736 35720 6469 35748
rect 5077 35683 5135 35689
rect 5077 35649 5089 35683
rect 5123 35649 5135 35683
rect 5077 35643 5135 35649
rect 3053 35615 3111 35621
rect 3053 35612 3065 35615
rect 2976 35584 3065 35612
rect 2976 35488 3004 35584
rect 3053 35581 3065 35584
rect 3099 35581 3111 35615
rect 3053 35575 3111 35581
rect 2958 35436 2964 35488
rect 3016 35436 3022 35488
rect 4525 35479 4583 35485
rect 4525 35445 4537 35479
rect 4571 35476 4583 35479
rect 4614 35476 4620 35488
rect 4571 35448 4620 35476
rect 4571 35445 4583 35448
rect 4525 35439 4583 35445
rect 4614 35436 4620 35448
rect 4672 35436 4678 35488
rect 5736 35476 5764 35720
rect 6457 35717 6469 35720
rect 6503 35717 6515 35751
rect 6457 35711 6515 35717
rect 6673 35751 6731 35757
rect 6673 35717 6685 35751
rect 6719 35748 6731 35751
rect 7929 35751 7987 35757
rect 7929 35748 7941 35751
rect 6719 35720 7941 35748
rect 6719 35717 6731 35720
rect 6673 35711 6731 35717
rect 7929 35717 7941 35720
rect 7975 35717 7987 35751
rect 7929 35711 7987 35717
rect 9490 35708 9496 35760
rect 9548 35708 9554 35760
rect 9766 35708 9772 35760
rect 9824 35708 9830 35760
rect 5813 35683 5871 35689
rect 5813 35649 5825 35683
rect 5859 35680 5871 35683
rect 7006 35680 7012 35692
rect 5859 35652 7012 35680
rect 5859 35649 5871 35652
rect 5813 35643 5871 35649
rect 7006 35640 7012 35652
rect 7064 35640 7070 35692
rect 7098 35640 7104 35692
rect 7156 35680 7162 35692
rect 7377 35683 7435 35689
rect 7377 35680 7389 35683
rect 7156 35652 7389 35680
rect 7156 35640 7162 35652
rect 7377 35649 7389 35652
rect 7423 35649 7435 35683
rect 7377 35643 7435 35649
rect 7561 35683 7619 35689
rect 7561 35649 7573 35683
rect 7607 35680 7619 35683
rect 7834 35680 7840 35692
rect 7607 35652 7840 35680
rect 7607 35649 7619 35652
rect 7561 35643 7619 35649
rect 7834 35640 7840 35652
rect 7892 35640 7898 35692
rect 8021 35683 8079 35689
rect 8021 35649 8033 35683
rect 8067 35649 8079 35683
rect 8021 35643 8079 35649
rect 5994 35572 6000 35624
rect 6052 35572 6058 35624
rect 6914 35572 6920 35624
rect 6972 35572 6978 35624
rect 7285 35615 7343 35621
rect 7285 35581 7297 35615
rect 7331 35612 7343 35615
rect 8036 35612 8064 35643
rect 8294 35640 8300 35692
rect 8352 35680 8358 35692
rect 8938 35680 8944 35692
rect 8352 35652 8944 35680
rect 8352 35640 8358 35652
rect 8938 35640 8944 35652
rect 8996 35640 9002 35692
rect 11164 35689 11192 35788
rect 11241 35785 11253 35819
rect 11287 35816 11299 35819
rect 12894 35816 12900 35828
rect 11287 35788 12900 35816
rect 11287 35785 11299 35788
rect 11241 35779 11299 35785
rect 12894 35776 12900 35788
rect 12952 35776 12958 35828
rect 13814 35776 13820 35828
rect 13872 35776 13878 35828
rect 13906 35776 13912 35828
rect 13964 35816 13970 35828
rect 14185 35819 14243 35825
rect 14185 35816 14197 35819
rect 13964 35788 14197 35816
rect 13964 35776 13970 35788
rect 14185 35785 14197 35788
rect 14231 35785 14243 35819
rect 14185 35779 14243 35785
rect 16666 35776 16672 35828
rect 16724 35776 16730 35828
rect 17862 35816 17868 35828
rect 17696 35788 17868 35816
rect 13832 35689 13860 35776
rect 13998 35708 14004 35760
rect 14056 35748 14062 35760
rect 14093 35751 14151 35757
rect 14093 35748 14105 35751
rect 14056 35720 14105 35748
rect 14056 35708 14062 35720
rect 14093 35717 14105 35720
rect 14139 35717 14151 35751
rect 14093 35711 14151 35717
rect 11149 35683 11207 35689
rect 11149 35649 11161 35683
rect 11195 35649 11207 35683
rect 11149 35643 11207 35649
rect 11333 35683 11391 35689
rect 11333 35649 11345 35683
rect 11379 35680 11391 35683
rect 11609 35683 11667 35689
rect 11609 35680 11621 35683
rect 11379 35652 11621 35680
rect 11379 35649 11391 35652
rect 11333 35643 11391 35649
rect 11609 35649 11621 35652
rect 11655 35649 11667 35683
rect 11609 35643 11667 35649
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35649 11759 35683
rect 11701 35643 11759 35649
rect 13817 35683 13875 35689
rect 13817 35649 13829 35683
rect 13863 35649 13875 35683
rect 13817 35643 13875 35649
rect 8386 35612 8392 35624
rect 7331 35584 8392 35612
rect 7331 35581 7343 35584
rect 7285 35575 7343 35581
rect 8386 35572 8392 35584
rect 8444 35572 8450 35624
rect 9217 35615 9275 35621
rect 9217 35581 9229 35615
rect 9263 35612 9275 35615
rect 9674 35612 9680 35624
rect 9263 35584 9680 35612
rect 9263 35581 9275 35584
rect 9217 35575 9275 35581
rect 9674 35572 9680 35584
rect 9732 35572 9738 35624
rect 11054 35572 11060 35624
rect 11112 35612 11118 35624
rect 11348 35612 11376 35643
rect 11112 35584 11376 35612
rect 11716 35612 11744 35643
rect 14550 35640 14556 35692
rect 14608 35680 14614 35692
rect 14734 35680 14740 35692
rect 14608 35652 14740 35680
rect 14608 35640 14614 35652
rect 14734 35640 14740 35652
rect 14792 35640 14798 35692
rect 16301 35683 16359 35689
rect 16301 35649 16313 35683
rect 16347 35680 16359 35683
rect 16684 35680 16712 35776
rect 17696 35757 17724 35788
rect 17862 35776 17868 35788
rect 17920 35776 17926 35828
rect 19426 35776 19432 35828
rect 19484 35816 19490 35828
rect 20073 35819 20131 35825
rect 20073 35816 20085 35819
rect 19484 35788 20085 35816
rect 19484 35776 19490 35788
rect 20073 35785 20085 35788
rect 20119 35785 20131 35819
rect 20073 35779 20131 35785
rect 20346 35776 20352 35828
rect 20404 35776 20410 35828
rect 20438 35776 20444 35828
rect 20496 35816 20502 35828
rect 20901 35819 20959 35825
rect 20901 35816 20913 35819
rect 20496 35788 20913 35816
rect 20496 35776 20502 35788
rect 20901 35785 20913 35788
rect 20947 35785 20959 35819
rect 20901 35779 20959 35785
rect 23845 35819 23903 35825
rect 23845 35785 23857 35819
rect 23891 35785 23903 35819
rect 23845 35779 23903 35785
rect 17681 35751 17739 35757
rect 17681 35717 17693 35751
rect 17727 35717 17739 35751
rect 17681 35711 17739 35717
rect 17954 35708 17960 35760
rect 18012 35748 18018 35760
rect 20364 35748 20392 35776
rect 20533 35751 20591 35757
rect 20533 35748 20545 35751
rect 18012 35720 18170 35748
rect 20364 35720 20545 35748
rect 18012 35708 18018 35720
rect 20533 35717 20545 35720
rect 20579 35717 20591 35751
rect 23860 35748 23888 35779
rect 24394 35776 24400 35828
rect 24452 35776 24458 35828
rect 25317 35819 25375 35825
rect 25317 35785 25329 35819
rect 25363 35816 25375 35819
rect 25774 35816 25780 35828
rect 25363 35788 25780 35816
rect 25363 35785 25375 35788
rect 25317 35779 25375 35785
rect 25774 35776 25780 35788
rect 25832 35776 25838 35828
rect 29917 35819 29975 35825
rect 29917 35785 29929 35819
rect 29963 35816 29975 35819
rect 30926 35816 30932 35828
rect 29963 35788 30932 35816
rect 29963 35785 29975 35788
rect 29917 35779 29975 35785
rect 30926 35776 30932 35788
rect 30984 35776 30990 35828
rect 31205 35819 31263 35825
rect 31205 35785 31217 35819
rect 31251 35816 31263 35819
rect 32398 35816 32404 35828
rect 31251 35788 32404 35816
rect 31251 35785 31263 35788
rect 31205 35779 31263 35785
rect 32398 35776 32404 35788
rect 32456 35776 32462 35828
rect 32677 35819 32735 35825
rect 32677 35785 32689 35819
rect 32723 35816 32735 35819
rect 32766 35816 32772 35828
rect 32723 35788 32772 35816
rect 32723 35785 32735 35788
rect 32677 35779 32735 35785
rect 32766 35776 32772 35788
rect 32824 35776 32830 35828
rect 32858 35776 32864 35828
rect 32916 35776 32922 35828
rect 33873 35819 33931 35825
rect 33873 35785 33885 35819
rect 33919 35816 33931 35819
rect 33962 35816 33968 35828
rect 33919 35788 33968 35816
rect 33919 35785 33931 35788
rect 33873 35779 33931 35785
rect 33962 35776 33968 35788
rect 34020 35776 34026 35828
rect 34054 35776 34060 35828
rect 34112 35816 34118 35828
rect 34333 35819 34391 35825
rect 34333 35816 34345 35819
rect 34112 35788 34345 35816
rect 34112 35776 34118 35788
rect 34333 35785 34345 35788
rect 34379 35785 34391 35819
rect 34333 35779 34391 35785
rect 34517 35819 34575 35825
rect 34517 35785 34529 35819
rect 34563 35816 34575 35819
rect 34606 35816 34612 35828
rect 34563 35788 34612 35816
rect 34563 35785 34575 35788
rect 34517 35779 34575 35785
rect 34606 35776 34612 35788
rect 34664 35776 34670 35828
rect 35710 35776 35716 35828
rect 35768 35776 35774 35828
rect 37918 35776 37924 35828
rect 37976 35816 37982 35828
rect 38378 35816 38384 35828
rect 37976 35788 38384 35816
rect 37976 35776 37982 35788
rect 38378 35776 38384 35788
rect 38436 35776 38442 35828
rect 24182 35751 24240 35757
rect 24182 35748 24194 35751
rect 23860 35720 24194 35748
rect 20533 35711 20591 35717
rect 24182 35717 24194 35720
rect 24228 35717 24240 35751
rect 24182 35711 24240 35717
rect 16347 35652 16712 35680
rect 17405 35683 17463 35689
rect 16347 35649 16359 35652
rect 16301 35643 16359 35649
rect 17405 35649 17417 35683
rect 17451 35649 17463 35683
rect 17405 35643 17463 35649
rect 11974 35612 11980 35624
rect 11716 35584 11980 35612
rect 11112 35572 11118 35584
rect 11974 35572 11980 35584
rect 12032 35612 12038 35624
rect 12526 35612 12532 35624
rect 12032 35584 12532 35612
rect 12032 35572 12038 35584
rect 12526 35572 12532 35584
rect 12584 35572 12590 35624
rect 15654 35572 15660 35624
rect 15712 35572 15718 35624
rect 16942 35572 16948 35624
rect 17000 35572 17006 35624
rect 17420 35612 17448 35643
rect 20898 35640 20904 35692
rect 20956 35680 20962 35692
rect 21453 35683 21511 35689
rect 21453 35680 21465 35683
rect 20956 35652 21465 35680
rect 20956 35640 20962 35652
rect 21453 35649 21465 35652
rect 21499 35649 21511 35683
rect 21453 35643 21511 35649
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35680 23719 35683
rect 24412 35680 24440 35776
rect 32493 35751 32551 35757
rect 32493 35717 32505 35751
rect 32539 35748 32551 35751
rect 32876 35748 32904 35776
rect 35437 35751 35495 35757
rect 32539 35720 32904 35748
rect 32968 35720 34192 35748
rect 32539 35717 32551 35720
rect 32493 35711 32551 35717
rect 23707 35652 24440 35680
rect 23707 35649 23719 35652
rect 23661 35643 23719 35649
rect 27614 35640 27620 35692
rect 27672 35680 27678 35692
rect 27985 35683 28043 35689
rect 27985 35680 27997 35683
rect 27672 35652 27997 35680
rect 27672 35640 27678 35652
rect 27985 35649 27997 35652
rect 28031 35649 28043 35683
rect 27985 35643 28043 35649
rect 29457 35683 29515 35689
rect 29457 35649 29469 35683
rect 29503 35680 29515 35683
rect 29546 35680 29552 35692
rect 29503 35652 29552 35680
rect 29503 35649 29515 35652
rect 29457 35643 29515 35649
rect 29546 35640 29552 35652
rect 29604 35680 29610 35692
rect 30006 35680 30012 35692
rect 29604 35652 30012 35680
rect 29604 35640 29610 35652
rect 30006 35640 30012 35652
rect 30064 35680 30070 35692
rect 30377 35683 30435 35689
rect 30377 35680 30389 35683
rect 30064 35652 30389 35680
rect 30064 35640 30070 35652
rect 30377 35649 30389 35652
rect 30423 35649 30435 35683
rect 30377 35643 30435 35649
rect 32401 35683 32459 35689
rect 32401 35649 32413 35683
rect 32447 35649 32459 35683
rect 32401 35643 32459 35649
rect 32585 35683 32643 35689
rect 32585 35649 32597 35683
rect 32631 35680 32643 35683
rect 32861 35683 32919 35689
rect 32861 35680 32873 35683
rect 32631 35652 32873 35680
rect 32631 35649 32643 35652
rect 32585 35643 32643 35649
rect 32861 35649 32873 35652
rect 32907 35680 32919 35683
rect 32968 35680 32996 35720
rect 34164 35692 34192 35720
rect 35437 35717 35449 35751
rect 35483 35748 35495 35751
rect 37182 35748 37188 35760
rect 35483 35720 37188 35748
rect 35483 35717 35495 35720
rect 35437 35711 35495 35717
rect 37182 35708 37188 35720
rect 37240 35708 37246 35760
rect 32907 35652 32996 35680
rect 33045 35683 33103 35689
rect 32907 35649 32919 35652
rect 32861 35643 32919 35649
rect 33045 35649 33057 35683
rect 33091 35649 33103 35683
rect 33045 35643 33103 35649
rect 17770 35612 17776 35624
rect 17420 35584 17776 35612
rect 17770 35572 17776 35584
rect 17828 35572 17834 35624
rect 20625 35615 20683 35621
rect 20625 35581 20637 35615
rect 20671 35612 20683 35615
rect 20671 35584 22094 35612
rect 20671 35581 20683 35584
rect 20625 35575 20683 35581
rect 7745 35547 7803 35553
rect 7745 35544 7757 35547
rect 6656 35516 7757 35544
rect 5810 35476 5816 35488
rect 5736 35448 5816 35476
rect 5810 35436 5816 35448
rect 5868 35436 5874 35488
rect 6656 35485 6684 35516
rect 7745 35513 7757 35516
rect 7791 35513 7803 35547
rect 7745 35507 7803 35513
rect 14093 35547 14151 35553
rect 14093 35513 14105 35547
rect 14139 35544 14151 35547
rect 15672 35544 15700 35572
rect 14139 35516 15700 35544
rect 16485 35547 16543 35553
rect 14139 35513 14151 35516
rect 14093 35507 14151 35513
rect 16485 35513 16497 35547
rect 16531 35544 16543 35547
rect 16960 35544 16988 35572
rect 16531 35516 16988 35544
rect 22066 35544 22094 35584
rect 22370 35572 22376 35624
rect 22428 35572 22434 35624
rect 23290 35572 23296 35624
rect 23348 35572 23354 35624
rect 23937 35615 23995 35621
rect 23937 35581 23949 35615
rect 23983 35581 23995 35615
rect 23937 35575 23995 35581
rect 27709 35615 27767 35621
rect 27709 35581 27721 35615
rect 27755 35581 27767 35615
rect 27709 35575 27767 35581
rect 29733 35615 29791 35621
rect 29733 35581 29745 35615
rect 29779 35612 29791 35615
rect 29914 35612 29920 35624
rect 29779 35584 29920 35612
rect 29779 35581 29791 35584
rect 29733 35575 29791 35581
rect 23308 35544 23336 35572
rect 22066 35516 23336 35544
rect 16531 35513 16543 35516
rect 16485 35507 16543 35513
rect 6641 35479 6699 35485
rect 6641 35445 6653 35479
rect 6687 35445 6699 35479
rect 6641 35439 6699 35445
rect 6825 35479 6883 35485
rect 6825 35445 6837 35479
rect 6871 35476 6883 35479
rect 6914 35476 6920 35488
rect 6871 35448 6920 35476
rect 6871 35445 6883 35448
rect 6825 35439 6883 35445
rect 6914 35436 6920 35448
rect 6972 35436 6978 35488
rect 9582 35436 9588 35488
rect 9640 35476 9646 35488
rect 10686 35476 10692 35488
rect 9640 35448 10692 35476
rect 9640 35436 9646 35448
rect 10686 35436 10692 35448
rect 10744 35436 10750 35488
rect 19150 35436 19156 35488
rect 19208 35436 19214 35488
rect 21542 35436 21548 35488
rect 21600 35476 21606 35488
rect 21821 35479 21879 35485
rect 21821 35476 21833 35479
rect 21600 35448 21833 35476
rect 21600 35436 21606 35448
rect 21821 35445 21833 35448
rect 21867 35445 21879 35479
rect 23952 35476 23980 35575
rect 27614 35504 27620 35556
rect 27672 35544 27678 35556
rect 27724 35544 27752 35575
rect 29914 35572 29920 35584
rect 29972 35572 29978 35624
rect 30282 35572 30288 35624
rect 30340 35572 30346 35624
rect 32416 35612 32444 35643
rect 33060 35612 33088 35643
rect 33410 35640 33416 35692
rect 33468 35680 33474 35692
rect 33505 35683 33563 35689
rect 33505 35680 33517 35683
rect 33468 35652 33517 35680
rect 33468 35640 33474 35652
rect 33505 35649 33517 35652
rect 33551 35680 33563 35683
rect 33965 35683 34023 35689
rect 33965 35680 33977 35683
rect 33551 35652 33977 35680
rect 33551 35649 33563 35652
rect 33505 35643 33563 35649
rect 33965 35649 33977 35652
rect 34011 35649 34023 35683
rect 33965 35643 34023 35649
rect 34146 35640 34152 35692
rect 34204 35640 34210 35692
rect 34698 35640 34704 35692
rect 34756 35680 34762 35692
rect 35069 35683 35127 35689
rect 35069 35680 35081 35683
rect 34756 35652 35081 35680
rect 34756 35640 34762 35652
rect 35069 35649 35081 35652
rect 35115 35649 35127 35683
rect 35069 35643 35127 35649
rect 32416 35584 33548 35612
rect 33520 35556 33548 35584
rect 33594 35572 33600 35624
rect 33652 35572 33658 35624
rect 37369 35615 37427 35621
rect 37369 35581 37381 35615
rect 37415 35612 37427 35615
rect 37734 35612 37740 35624
rect 37415 35584 37740 35612
rect 37415 35581 37427 35584
rect 37369 35575 37427 35581
rect 37734 35572 37740 35584
rect 37792 35612 37798 35624
rect 38470 35612 38476 35624
rect 37792 35584 38476 35612
rect 37792 35572 37798 35584
rect 38470 35572 38476 35584
rect 38528 35572 38534 35624
rect 41506 35572 41512 35624
rect 41564 35572 41570 35624
rect 27672 35516 27752 35544
rect 29549 35547 29607 35553
rect 27672 35504 27678 35516
rect 29549 35513 29561 35547
rect 29595 35544 29607 35547
rect 29822 35544 29828 35556
rect 29595 35516 29828 35544
rect 29595 35513 29607 35516
rect 29549 35507 29607 35513
rect 29822 35504 29828 35516
rect 29880 35544 29886 35556
rect 30098 35544 30104 35556
rect 29880 35516 30104 35544
rect 29880 35504 29886 35516
rect 30098 35504 30104 35516
rect 30156 35504 30162 35556
rect 33502 35504 33508 35556
rect 33560 35504 33566 35556
rect 25222 35476 25228 35488
rect 23952 35448 25228 35476
rect 21821 35439 21879 35445
rect 25222 35436 25228 35448
rect 25280 35476 25286 35488
rect 25866 35476 25872 35488
rect 25280 35448 25872 35476
rect 25280 35436 25286 35448
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 40954 35436 40960 35488
rect 41012 35436 41018 35488
rect 1104 35386 45172 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 45172 35386
rect 1104 35312 45172 35334
rect 3326 35232 3332 35284
rect 3384 35272 3390 35284
rect 3421 35275 3479 35281
rect 3421 35272 3433 35275
rect 3384 35244 3433 35272
rect 3384 35232 3390 35244
rect 3421 35241 3433 35244
rect 3467 35241 3479 35275
rect 4614 35272 4620 35284
rect 3421 35235 3479 35241
rect 4264 35244 4620 35272
rect 3881 35207 3939 35213
rect 3881 35173 3893 35207
rect 3927 35173 3939 35207
rect 3881 35167 3939 35173
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 2958 35068 2964 35080
rect 1719 35040 2964 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 2958 35028 2964 35040
rect 3016 35028 3022 35080
rect 3605 35071 3663 35077
rect 3605 35037 3617 35071
rect 3651 35068 3663 35071
rect 3896 35068 3924 35167
rect 4264 35080 4292 35244
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 4798 35232 4804 35284
rect 4856 35232 4862 35284
rect 6546 35232 6552 35284
rect 6604 35272 6610 35284
rect 6825 35275 6883 35281
rect 6825 35272 6837 35275
rect 6604 35244 6837 35272
rect 6604 35232 6610 35244
rect 6825 35241 6837 35244
rect 6871 35241 6883 35275
rect 6825 35235 6883 35241
rect 6914 35232 6920 35284
rect 6972 35232 6978 35284
rect 9217 35275 9275 35281
rect 9217 35241 9229 35275
rect 9263 35272 9275 35275
rect 9306 35272 9312 35284
rect 9263 35244 9312 35272
rect 9263 35241 9275 35244
rect 9217 35235 9275 35241
rect 9306 35232 9312 35244
rect 9364 35232 9370 35284
rect 9401 35275 9459 35281
rect 9401 35241 9413 35275
rect 9447 35272 9459 35275
rect 9858 35272 9864 35284
rect 9447 35244 9864 35272
rect 9447 35241 9459 35244
rect 9401 35235 9459 35241
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 10686 35232 10692 35284
rect 10744 35232 10750 35284
rect 17865 35275 17923 35281
rect 17865 35241 17877 35275
rect 17911 35272 17923 35275
rect 18046 35272 18052 35284
rect 17911 35244 18052 35272
rect 17911 35241 17923 35244
rect 17865 35235 17923 35241
rect 18046 35232 18052 35244
rect 18104 35232 18110 35284
rect 19150 35232 19156 35284
rect 19208 35232 19214 35284
rect 22005 35275 22063 35281
rect 22005 35241 22017 35275
rect 22051 35272 22063 35275
rect 22370 35272 22376 35284
rect 22051 35244 22376 35272
rect 22051 35241 22063 35244
rect 22005 35235 22063 35241
rect 22370 35232 22376 35244
rect 22428 35232 22434 35284
rect 24213 35275 24271 35281
rect 24213 35241 24225 35275
rect 24259 35272 24271 35275
rect 25881 35275 25939 35281
rect 25881 35272 25893 35275
rect 24259 35244 25893 35272
rect 24259 35241 24271 35244
rect 24213 35235 24271 35241
rect 25881 35241 25893 35244
rect 25927 35241 25939 35275
rect 25881 35235 25939 35241
rect 26142 35232 26148 35284
rect 26200 35272 26206 35284
rect 26200 35244 30236 35272
rect 26200 35232 26206 35244
rect 4816 35204 4844 35232
rect 4540 35176 4844 35204
rect 4540 35145 4568 35176
rect 4525 35139 4583 35145
rect 4525 35105 4537 35139
rect 4571 35136 4583 35139
rect 4614 35136 4620 35148
rect 4571 35108 4620 35136
rect 4571 35105 4583 35108
rect 4525 35099 4583 35105
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 6178 35136 6184 35148
rect 4724 35108 6184 35136
rect 3651 35040 3924 35068
rect 3651 35037 3663 35040
rect 3605 35031 3663 35037
rect 4246 35028 4252 35080
rect 4304 35028 4310 35080
rect 4724 35077 4752 35108
rect 6178 35096 6184 35108
rect 6236 35096 6242 35148
rect 4709 35071 4767 35077
rect 4709 35037 4721 35071
rect 4755 35037 4767 35071
rect 6932 35068 6960 35232
rect 7009 35071 7067 35077
rect 7009 35068 7021 35071
rect 6932 35040 7021 35068
rect 4709 35031 4767 35037
rect 7009 35037 7021 35040
rect 7055 35037 7067 35071
rect 10704 35068 10732 35232
rect 12434 35204 12440 35216
rect 12406 35164 12440 35204
rect 12492 35204 12498 35216
rect 13170 35204 13176 35216
rect 12492 35176 13176 35204
rect 12492 35164 12498 35176
rect 13170 35164 13176 35176
rect 13228 35164 13234 35216
rect 11701 35071 11759 35077
rect 11701 35068 11713 35071
rect 10704 35040 11713 35068
rect 7009 35031 7067 35037
rect 11701 35037 11713 35040
rect 11747 35037 11759 35071
rect 11701 35031 11759 35037
rect 1940 35003 1998 35009
rect 1940 34969 1952 35003
rect 1986 35000 1998 35003
rect 2130 35000 2136 35012
rect 1986 34972 2136 35000
rect 1986 34969 1998 34972
rect 1940 34963 1998 34969
rect 2130 34960 2136 34972
rect 2188 34960 2194 35012
rect 2976 35000 3004 35028
rect 4724 35000 4752 35031
rect 2976 34972 4752 35000
rect 4985 35003 5043 35009
rect 4985 34969 4997 35003
rect 5031 35000 5043 35003
rect 5074 35000 5080 35012
rect 5031 34972 5080 35000
rect 5031 34969 5043 34972
rect 4985 34963 5043 34969
rect 5074 34960 5080 34972
rect 5132 34960 5138 35012
rect 5534 34960 5540 35012
rect 5592 34960 5598 35012
rect 9033 35003 9091 35009
rect 9033 35000 9045 35003
rect 6380 34972 9045 35000
rect 3050 34892 3056 34944
rect 3108 34892 3114 34944
rect 4341 34935 4399 34941
rect 4341 34901 4353 34935
rect 4387 34932 4399 34935
rect 5350 34932 5356 34944
rect 4387 34904 5356 34932
rect 4387 34901 4399 34904
rect 4341 34895 4399 34901
rect 5350 34892 5356 34904
rect 5408 34892 5414 34944
rect 5810 34892 5816 34944
rect 5868 34932 5874 34944
rect 6380 34932 6408 34972
rect 9033 34969 9045 34972
rect 9079 34969 9091 35003
rect 9033 34963 9091 34969
rect 9249 35003 9307 35009
rect 9249 34969 9261 35003
rect 9295 35000 9307 35003
rect 9490 35000 9496 35012
rect 9295 34972 9496 35000
rect 9295 34969 9307 34972
rect 9249 34963 9307 34969
rect 5868 34904 6408 34932
rect 6457 34935 6515 34941
rect 5868 34892 5874 34904
rect 6457 34901 6469 34935
rect 6503 34932 6515 34935
rect 6914 34932 6920 34944
rect 6503 34904 6920 34932
rect 6503 34901 6515 34904
rect 6457 34895 6515 34901
rect 6914 34892 6920 34904
rect 6972 34892 6978 34944
rect 9048 34932 9076 34963
rect 9490 34960 9496 34972
rect 9548 34960 9554 35012
rect 12406 35000 12434 35164
rect 18138 35096 18144 35148
rect 18196 35136 18202 35148
rect 18325 35139 18383 35145
rect 18325 35136 18337 35139
rect 18196 35108 18337 35136
rect 18196 35096 18202 35108
rect 18325 35105 18337 35108
rect 18371 35105 18383 35139
rect 18325 35099 18383 35105
rect 18414 35096 18420 35148
rect 18472 35096 18478 35148
rect 18230 35028 18236 35080
rect 18288 35068 18294 35080
rect 19168 35068 19196 35232
rect 30208 35204 30236 35244
rect 30282 35232 30288 35284
rect 30340 35232 30346 35284
rect 33594 35232 33600 35284
rect 33652 35272 33658 35284
rect 33781 35275 33839 35281
rect 33781 35272 33793 35275
rect 33652 35244 33793 35272
rect 33652 35232 33658 35244
rect 33781 35241 33793 35244
rect 33827 35241 33839 35275
rect 33781 35235 33839 35241
rect 34146 35232 34152 35284
rect 34204 35232 34210 35284
rect 35710 35232 35716 35284
rect 35768 35232 35774 35284
rect 33229 35207 33287 35213
rect 30208 35176 31754 35204
rect 22462 35096 22468 35148
rect 22520 35096 22526 35148
rect 22649 35139 22707 35145
rect 22649 35105 22661 35139
rect 22695 35136 22707 35139
rect 23290 35136 23296 35148
rect 22695 35108 23296 35136
rect 22695 35105 22707 35108
rect 22649 35099 22707 35105
rect 23290 35096 23296 35108
rect 23348 35096 23354 35148
rect 25866 35096 25872 35148
rect 25924 35136 25930 35148
rect 26145 35139 26203 35145
rect 26145 35136 26157 35139
rect 25924 35108 26157 35136
rect 25924 35096 25930 35108
rect 26145 35105 26157 35108
rect 26191 35105 26203 35139
rect 26145 35099 26203 35105
rect 27798 35096 27804 35148
rect 27856 35136 27862 35148
rect 28169 35139 28227 35145
rect 28169 35136 28181 35139
rect 27856 35108 28181 35136
rect 27856 35096 27862 35108
rect 28169 35105 28181 35108
rect 28215 35105 28227 35139
rect 28169 35099 28227 35105
rect 18288 35040 19196 35068
rect 18288 35028 18294 35040
rect 19426 35028 19432 35080
rect 19484 35068 19490 35080
rect 20441 35071 20499 35077
rect 20441 35068 20453 35071
rect 19484 35040 20453 35068
rect 19484 35028 19490 35040
rect 20441 35037 20453 35040
rect 20487 35037 20499 35071
rect 20441 35031 20499 35037
rect 23382 35028 23388 35080
rect 23440 35028 23446 35080
rect 24026 35028 24032 35080
rect 24084 35028 24090 35080
rect 29914 35028 29920 35080
rect 29972 35028 29978 35080
rect 30098 35028 30104 35080
rect 30156 35068 30162 35080
rect 30156 35040 30328 35068
rect 30156 35028 30162 35040
rect 11717 34972 12434 35000
rect 11717 34932 11745 34972
rect 22094 34960 22100 35012
rect 22152 35000 22158 35012
rect 22373 35003 22431 35009
rect 22373 35000 22385 35003
rect 22152 34972 22385 35000
rect 22152 34960 22158 34972
rect 22373 34969 22385 34972
rect 22419 35000 22431 35003
rect 22833 35003 22891 35009
rect 22833 35000 22845 35003
rect 22419 34972 22845 35000
rect 22419 34969 22431 34972
rect 22373 34963 22431 34969
rect 22833 34969 22845 34972
rect 22879 34969 22891 35003
rect 25438 34972 26726 35000
rect 22833 34963 22891 34969
rect 26068 34944 26096 34972
rect 27890 34960 27896 35012
rect 27948 34960 27954 35012
rect 30300 34944 30328 35040
rect 9048 34904 11745 34932
rect 11793 34935 11851 34941
rect 11793 34901 11805 34935
rect 11839 34932 11851 34935
rect 12250 34932 12256 34944
rect 11839 34904 12256 34932
rect 11839 34901 11851 34904
rect 11793 34895 11851 34901
rect 12250 34892 12256 34904
rect 12308 34892 12314 34944
rect 19889 34935 19947 34941
rect 19889 34901 19901 34935
rect 19935 34932 19947 34935
rect 19978 34932 19984 34944
rect 19935 34904 19984 34932
rect 19935 34901 19947 34904
rect 19889 34895 19947 34901
rect 19978 34892 19984 34904
rect 20036 34892 20042 34944
rect 24397 34935 24455 34941
rect 24397 34901 24409 34935
rect 24443 34932 24455 34935
rect 24578 34932 24584 34944
rect 24443 34904 24584 34932
rect 24443 34901 24455 34904
rect 24397 34895 24455 34901
rect 24578 34892 24584 34904
rect 24636 34892 24642 34944
rect 26050 34892 26056 34944
rect 26108 34892 26114 34944
rect 26421 34935 26479 34941
rect 26421 34901 26433 34935
rect 26467 34932 26479 34935
rect 26510 34932 26516 34944
rect 26467 34904 26516 34932
rect 26467 34901 26479 34904
rect 26421 34895 26479 34901
rect 26510 34892 26516 34904
rect 26568 34892 26574 34944
rect 26602 34892 26608 34944
rect 26660 34932 26666 34944
rect 28074 34932 28080 34944
rect 26660 34904 28080 34932
rect 26660 34892 26666 34904
rect 28074 34892 28080 34904
rect 28132 34892 28138 34944
rect 30282 34892 30288 34944
rect 30340 34892 30346 34944
rect 31726 34932 31754 35176
rect 33229 35173 33241 35207
rect 33275 35204 33287 35207
rect 34164 35204 34192 35232
rect 33275 35176 34192 35204
rect 33275 35173 33287 35176
rect 33229 35167 33287 35173
rect 33689 35139 33747 35145
rect 33689 35136 33701 35139
rect 33152 35108 33701 35136
rect 33152 35080 33180 35108
rect 33689 35105 33701 35108
rect 33735 35105 33747 35139
rect 33689 35099 33747 35105
rect 33134 35028 33140 35080
rect 33192 35028 33198 35080
rect 33318 35028 33324 35080
rect 33376 35028 33382 35080
rect 33502 35028 33508 35080
rect 33560 35068 33566 35080
rect 33873 35071 33931 35077
rect 33873 35068 33885 35071
rect 33560 35040 33885 35068
rect 33560 35028 33566 35040
rect 33873 35037 33885 35040
rect 33919 35037 33931 35071
rect 33873 35031 33931 35037
rect 33965 35071 34023 35077
rect 33965 35037 33977 35071
rect 34011 35068 34023 35071
rect 34164 35068 34192 35176
rect 34011 35040 34192 35068
rect 35728 35068 35756 35232
rect 40218 35096 40224 35148
rect 40276 35136 40282 35148
rect 40681 35139 40739 35145
rect 40681 35136 40693 35139
rect 40276 35108 40693 35136
rect 40276 35096 40282 35108
rect 40681 35105 40693 35108
rect 40727 35105 40739 35139
rect 40681 35099 40739 35105
rect 40954 35096 40960 35148
rect 41012 35096 41018 35148
rect 42429 35139 42487 35145
rect 42429 35105 42441 35139
rect 42475 35136 42487 35139
rect 43073 35139 43131 35145
rect 43073 35136 43085 35139
rect 42475 35108 43085 35136
rect 42475 35105 42487 35108
rect 42429 35099 42487 35105
rect 43073 35105 43085 35108
rect 43119 35105 43131 35139
rect 43073 35099 43131 35105
rect 35728 35040 35834 35068
rect 34011 35037 34023 35040
rect 33965 35031 34023 35037
rect 37182 35028 37188 35080
rect 37240 35028 37246 35080
rect 38654 35028 38660 35080
rect 38712 35028 38718 35080
rect 40034 35028 40040 35080
rect 40092 35068 40098 35080
rect 40405 35071 40463 35077
rect 40405 35068 40417 35071
rect 40092 35040 40417 35068
rect 40092 35028 40098 35040
rect 40405 35037 40417 35040
rect 40451 35037 40463 35071
rect 40405 35031 40463 35037
rect 44821 35071 44879 35077
rect 44821 35037 44833 35071
rect 44867 35068 44879 35071
rect 44867 35040 45324 35068
rect 44867 35037 44879 35040
rect 44821 35031 44879 35037
rect 36909 35003 36967 35009
rect 36909 34969 36921 35003
rect 36955 34969 36967 35003
rect 36909 34963 36967 34969
rect 35437 34935 35495 34941
rect 35437 34932 35449 34935
rect 31726 34904 35449 34932
rect 35437 34901 35449 34904
rect 35483 34932 35495 34935
rect 36170 34932 36176 34944
rect 35483 34904 36176 34932
rect 35483 34901 35495 34904
rect 35437 34895 35495 34901
rect 36170 34892 36176 34904
rect 36228 34892 36234 34944
rect 36262 34892 36268 34944
rect 36320 34932 36326 34944
rect 36924 34932 36952 34963
rect 39298 34960 39304 35012
rect 39356 35000 39362 35012
rect 39356 34972 41446 35000
rect 39356 34960 39362 34972
rect 45296 34944 45324 35040
rect 36320 34904 36952 34932
rect 36320 34892 36326 34904
rect 38010 34892 38016 34944
rect 38068 34932 38074 34944
rect 38105 34935 38163 34941
rect 38105 34932 38117 34935
rect 38068 34904 38117 34932
rect 38068 34892 38074 34904
rect 38105 34901 38117 34904
rect 38151 34901 38163 34935
rect 38105 34895 38163 34901
rect 38746 34892 38752 34944
rect 38804 34932 38810 34944
rect 39853 34935 39911 34941
rect 39853 34932 39865 34935
rect 38804 34904 39865 34932
rect 38804 34892 38810 34904
rect 39853 34901 39865 34904
rect 39899 34901 39911 34935
rect 39853 34895 39911 34901
rect 41966 34892 41972 34944
rect 42024 34932 42030 34944
rect 42521 34935 42579 34941
rect 42521 34932 42533 34935
rect 42024 34904 42533 34932
rect 42024 34892 42030 34904
rect 42521 34901 42533 34904
rect 42567 34901 42579 34935
rect 42521 34895 42579 34901
rect 44082 34892 44088 34944
rect 44140 34932 44146 34944
rect 44637 34935 44695 34941
rect 44637 34932 44649 34935
rect 44140 34904 44649 34932
rect 44140 34892 44146 34904
rect 44637 34901 44649 34904
rect 44683 34901 44695 34935
rect 44637 34895 44695 34901
rect 45278 34892 45284 34944
rect 45336 34892 45342 34944
rect 1104 34842 45172 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 45172 34842
rect 1104 34768 45172 34790
rect 2130 34688 2136 34740
rect 2188 34688 2194 34740
rect 2685 34731 2743 34737
rect 2685 34697 2697 34731
rect 2731 34697 2743 34731
rect 2685 34691 2743 34697
rect 3145 34731 3203 34737
rect 3145 34697 3157 34731
rect 3191 34728 3203 34731
rect 4246 34728 4252 34740
rect 3191 34700 4252 34728
rect 3191 34697 3203 34700
rect 3145 34691 3203 34697
rect 2317 34595 2375 34601
rect 2317 34561 2329 34595
rect 2363 34592 2375 34595
rect 2700 34592 2728 34691
rect 4246 34688 4252 34700
rect 4304 34688 4310 34740
rect 13262 34688 13268 34740
rect 13320 34728 13326 34740
rect 13320 34700 14136 34728
rect 13320 34688 13326 34700
rect 13722 34660 13728 34672
rect 13096 34632 13728 34660
rect 2363 34564 2728 34592
rect 3053 34595 3111 34601
rect 2363 34561 2375 34564
rect 2317 34555 2375 34561
rect 3053 34561 3065 34595
rect 3099 34592 3111 34595
rect 3786 34592 3792 34604
rect 3099 34564 3792 34592
rect 3099 34561 3111 34564
rect 3053 34555 3111 34561
rect 3786 34552 3792 34564
rect 3844 34552 3850 34604
rect 5166 34552 5172 34604
rect 5224 34592 5230 34604
rect 5353 34595 5411 34601
rect 5353 34592 5365 34595
rect 5224 34564 5365 34592
rect 5224 34552 5230 34564
rect 5353 34561 5365 34564
rect 5399 34561 5411 34595
rect 5353 34555 5411 34561
rect 7558 34552 7564 34604
rect 7616 34552 7622 34604
rect 8570 34552 8576 34604
rect 8628 34552 8634 34604
rect 10137 34595 10195 34601
rect 10137 34561 10149 34595
rect 10183 34592 10195 34595
rect 10226 34592 10232 34604
rect 10183 34564 10232 34592
rect 10183 34561 10195 34564
rect 10137 34555 10195 34561
rect 10226 34552 10232 34564
rect 10284 34552 10290 34604
rect 13096 34601 13124 34632
rect 13722 34620 13728 34632
rect 13780 34660 13786 34672
rect 13780 34632 13952 34660
rect 13780 34620 13786 34632
rect 13081 34595 13139 34601
rect 13081 34561 13093 34595
rect 13127 34561 13139 34595
rect 13081 34555 13139 34561
rect 13173 34595 13231 34601
rect 13173 34561 13185 34595
rect 13219 34592 13231 34595
rect 13262 34592 13268 34604
rect 13219 34564 13268 34592
rect 13219 34561 13231 34564
rect 13173 34555 13231 34561
rect 13262 34552 13268 34564
rect 13320 34552 13326 34604
rect 13354 34552 13360 34604
rect 13412 34592 13418 34604
rect 13924 34601 13952 34632
rect 14108 34601 14136 34700
rect 14550 34688 14556 34740
rect 14608 34728 14614 34740
rect 16850 34728 16856 34740
rect 14608 34700 16856 34728
rect 14608 34688 14614 34700
rect 16850 34688 16856 34700
rect 16908 34728 16914 34740
rect 18046 34728 18052 34740
rect 16908 34700 18052 34728
rect 16908 34688 16914 34700
rect 18046 34688 18052 34700
rect 18104 34688 18110 34740
rect 18230 34688 18236 34740
rect 18288 34688 18294 34740
rect 19426 34688 19432 34740
rect 19484 34728 19490 34740
rect 19889 34731 19947 34737
rect 19889 34728 19901 34731
rect 19484 34700 19901 34728
rect 19484 34688 19490 34700
rect 19889 34697 19901 34700
rect 19935 34697 19947 34731
rect 19889 34691 19947 34697
rect 19978 34688 19984 34740
rect 20036 34688 20042 34740
rect 20349 34731 20407 34737
rect 20349 34697 20361 34731
rect 20395 34728 20407 34731
rect 20438 34728 20444 34740
rect 20395 34700 20444 34728
rect 20395 34697 20407 34700
rect 20349 34691 20407 34697
rect 20438 34688 20444 34700
rect 20496 34688 20502 34740
rect 21542 34688 21548 34740
rect 21600 34688 21606 34740
rect 21637 34731 21695 34737
rect 21637 34697 21649 34731
rect 21683 34728 21695 34731
rect 23201 34731 23259 34737
rect 21683 34700 22094 34728
rect 21683 34697 21695 34700
rect 21637 34691 21695 34697
rect 13541 34595 13599 34601
rect 13541 34592 13553 34595
rect 13412 34564 13553 34592
rect 13412 34552 13418 34564
rect 13541 34561 13553 34564
rect 13587 34592 13599 34595
rect 13633 34595 13691 34601
rect 13633 34592 13645 34595
rect 13587 34564 13645 34592
rect 13587 34561 13599 34564
rect 13541 34555 13599 34561
rect 13633 34561 13645 34564
rect 13679 34561 13691 34595
rect 13633 34555 13691 34561
rect 13817 34595 13875 34601
rect 13817 34561 13829 34595
rect 13863 34561 13875 34595
rect 13817 34555 13875 34561
rect 13909 34595 13967 34601
rect 13909 34561 13921 34595
rect 13955 34561 13967 34595
rect 13909 34555 13967 34561
rect 14093 34595 14151 34601
rect 14093 34561 14105 34595
rect 14139 34561 14151 34595
rect 14093 34555 14151 34561
rect 3329 34527 3387 34533
rect 3329 34493 3341 34527
rect 3375 34493 3387 34527
rect 3329 34487 3387 34493
rect 2866 34416 2872 34468
rect 2924 34456 2930 34468
rect 3344 34456 3372 34487
rect 8846 34484 8852 34536
rect 8904 34484 8910 34536
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13832 34524 13860 34555
rect 14182 34552 14188 34604
rect 14240 34552 14246 34604
rect 17957 34595 18015 34601
rect 17957 34561 17969 34595
rect 18003 34592 18015 34595
rect 18248 34592 18276 34688
rect 18003 34564 18276 34592
rect 19797 34595 19855 34601
rect 18003 34561 18015 34564
rect 17957 34555 18015 34561
rect 19797 34561 19809 34595
rect 19843 34592 19855 34595
rect 19996 34592 20024 34688
rect 19843 34564 20024 34592
rect 19843 34561 19855 34564
rect 19797 34555 19855 34561
rect 20254 34552 20260 34604
rect 20312 34552 20318 34604
rect 21453 34595 21511 34601
rect 21453 34561 21465 34595
rect 21499 34592 21511 34595
rect 21560 34592 21588 34688
rect 22066 34669 22094 34700
rect 23201 34697 23213 34731
rect 23247 34728 23259 34731
rect 23382 34728 23388 34740
rect 23247 34700 23388 34728
rect 23247 34697 23259 34700
rect 23201 34691 23259 34697
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 24026 34688 24032 34740
rect 24084 34728 24090 34740
rect 24305 34731 24363 34737
rect 24305 34728 24317 34731
rect 24084 34700 24317 34728
rect 24084 34688 24090 34700
rect 24305 34697 24317 34700
rect 24351 34697 24363 34731
rect 24305 34691 24363 34697
rect 24762 34688 24768 34740
rect 24820 34688 24826 34740
rect 27801 34731 27859 34737
rect 27801 34697 27813 34731
rect 27847 34728 27859 34731
rect 27890 34728 27896 34740
rect 27847 34700 27896 34728
rect 27847 34697 27859 34700
rect 27801 34691 27859 34697
rect 27890 34688 27896 34700
rect 27948 34688 27954 34740
rect 33134 34688 33140 34740
rect 33192 34688 33198 34740
rect 33318 34688 33324 34740
rect 33376 34728 33382 34740
rect 33689 34731 33747 34737
rect 33689 34728 33701 34731
rect 33376 34700 33701 34728
rect 33376 34688 33382 34700
rect 33689 34697 33701 34700
rect 33735 34697 33747 34731
rect 33689 34691 33747 34697
rect 36262 34688 36268 34740
rect 36320 34688 36326 34740
rect 36449 34731 36507 34737
rect 36449 34697 36461 34731
rect 36495 34697 36507 34731
rect 36449 34691 36507 34697
rect 38197 34731 38255 34737
rect 38197 34697 38209 34731
rect 38243 34728 38255 34731
rect 38654 34728 38660 34740
rect 38243 34700 38660 34728
rect 38243 34697 38255 34700
rect 38197 34691 38255 34697
rect 22066 34663 22124 34669
rect 22066 34629 22078 34663
rect 22112 34629 22124 34663
rect 22066 34623 22124 34629
rect 26418 34620 26424 34672
rect 26476 34620 26482 34672
rect 28534 34660 28540 34672
rect 26620 34632 28540 34660
rect 21499 34564 21588 34592
rect 21499 34561 21511 34564
rect 21453 34555 21511 34561
rect 22646 34552 22652 34604
rect 22704 34592 22710 34604
rect 23385 34595 23443 34601
rect 23385 34592 23397 34595
rect 22704 34564 23397 34592
rect 22704 34552 22710 34564
rect 23385 34561 23397 34564
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 24670 34552 24676 34604
rect 24728 34552 24734 34604
rect 26234 34552 26240 34604
rect 26292 34552 26298 34604
rect 26510 34552 26516 34604
rect 26568 34552 26574 34604
rect 26620 34601 26648 34632
rect 27632 34604 27660 34632
rect 28534 34620 28540 34632
rect 28592 34660 28598 34672
rect 31662 34660 31668 34672
rect 28592 34632 31668 34660
rect 28592 34620 28598 34632
rect 31662 34620 31668 34632
rect 31720 34620 31726 34672
rect 32582 34660 32588 34672
rect 32140 34632 32588 34660
rect 26605 34595 26663 34601
rect 26605 34561 26617 34595
rect 26651 34561 26663 34595
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 26605 34555 26663 34561
rect 26804 34564 27169 34592
rect 14200 34524 14228 34552
rect 13495 34496 14228 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 17862 34484 17868 34536
rect 17920 34484 17926 34536
rect 18414 34484 18420 34536
rect 18472 34484 18478 34536
rect 20441 34527 20499 34533
rect 20441 34493 20453 34527
rect 20487 34493 20499 34527
rect 20441 34487 20499 34493
rect 5718 34456 5724 34468
rect 2924 34428 5724 34456
rect 2924 34416 2930 34428
rect 5718 34416 5724 34428
rect 5776 34416 5782 34468
rect 12434 34416 12440 34468
rect 12492 34456 12498 34468
rect 13633 34459 13691 34465
rect 13633 34456 13645 34459
rect 12492 34428 13645 34456
rect 12492 34416 12498 34428
rect 13633 34425 13645 34428
rect 13679 34425 13691 34459
rect 18432 34456 18460 34484
rect 20456 34456 20484 34487
rect 20990 34484 20996 34536
rect 21048 34524 21054 34536
rect 21821 34527 21879 34533
rect 21821 34524 21833 34527
rect 21048 34496 21833 34524
rect 21048 34484 21054 34496
rect 21821 34493 21833 34496
rect 21867 34493 21879 34527
rect 24486 34524 24492 34536
rect 21821 34487 21879 34493
rect 23492 34496 24492 34524
rect 18432 34428 20484 34456
rect 13633 34419 13691 34425
rect 4798 34348 4804 34400
rect 4856 34348 4862 34400
rect 7374 34348 7380 34400
rect 7432 34348 7438 34400
rect 8754 34348 8760 34400
rect 8812 34348 8818 34400
rect 9490 34348 9496 34400
rect 9548 34348 9554 34400
rect 9861 34391 9919 34397
rect 9861 34357 9873 34391
rect 9907 34388 9919 34391
rect 9950 34388 9956 34400
rect 9907 34360 9956 34388
rect 9907 34357 9919 34360
rect 9861 34351 9919 34357
rect 9950 34348 9956 34360
rect 10008 34348 10014 34400
rect 12894 34348 12900 34400
rect 12952 34348 12958 34400
rect 13814 34348 13820 34400
rect 13872 34388 13878 34400
rect 14001 34391 14059 34397
rect 14001 34388 14013 34391
rect 13872 34360 14013 34388
rect 13872 34348 13878 34360
rect 14001 34357 14013 34360
rect 14047 34357 14059 34391
rect 14001 34351 14059 34357
rect 14274 34348 14280 34400
rect 14332 34388 14338 34400
rect 15746 34388 15752 34400
rect 14332 34360 15752 34388
rect 14332 34348 14338 34360
rect 15746 34348 15752 34360
rect 15804 34348 15810 34400
rect 16114 34348 16120 34400
rect 16172 34388 16178 34400
rect 17034 34388 17040 34400
rect 16172 34360 17040 34388
rect 16172 34348 16178 34360
rect 17034 34348 17040 34360
rect 17092 34348 17098 34400
rect 19610 34348 19616 34400
rect 19668 34348 19674 34400
rect 20456 34388 20484 34428
rect 21082 34388 21088 34400
rect 20456 34360 21088 34388
rect 21082 34348 21088 34360
rect 21140 34388 21146 34400
rect 22002 34388 22008 34400
rect 21140 34360 22008 34388
rect 21140 34348 21146 34360
rect 22002 34348 22008 34360
rect 22060 34388 22066 34400
rect 23492 34397 23520 34496
rect 24486 34484 24492 34496
rect 24544 34524 24550 34536
rect 24857 34527 24915 34533
rect 24857 34524 24869 34527
rect 24544 34496 24869 34524
rect 24544 34484 24550 34496
rect 24857 34493 24869 34496
rect 24903 34493 24915 34527
rect 26528 34524 26556 34552
rect 26528 34496 26740 34524
rect 24857 34487 24915 34493
rect 23477 34391 23535 34397
rect 23477 34388 23489 34391
rect 22060 34360 23489 34388
rect 22060 34348 22066 34360
rect 23477 34357 23489 34360
rect 23523 34357 23535 34391
rect 26712 34388 26740 34496
rect 26804 34465 26832 34564
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 27157 34555 27215 34561
rect 27614 34552 27620 34604
rect 27672 34552 27678 34604
rect 28166 34552 28172 34604
rect 28224 34552 28230 34604
rect 32140 34601 32168 34632
rect 32582 34620 32588 34632
rect 32640 34620 32646 34672
rect 36280 34660 36308 34688
rect 36357 34663 36415 34669
rect 36357 34660 36369 34663
rect 36280 34632 36369 34660
rect 36357 34629 36369 34632
rect 36403 34629 36415 34663
rect 36357 34623 36415 34629
rect 32125 34595 32183 34601
rect 32125 34561 32137 34595
rect 32171 34561 32183 34595
rect 32125 34555 32183 34561
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34592 32367 34595
rect 33226 34592 33232 34604
rect 32355 34564 33232 34592
rect 32355 34561 32367 34564
rect 32309 34555 32367 34561
rect 33226 34552 33232 34564
rect 33284 34552 33290 34604
rect 33321 34595 33379 34601
rect 33321 34561 33333 34595
rect 33367 34561 33379 34595
rect 33321 34555 33379 34561
rect 33505 34595 33563 34601
rect 33505 34561 33517 34595
rect 33551 34592 33563 34595
rect 33594 34592 33600 34604
rect 33551 34564 33600 34592
rect 33551 34561 33563 34564
rect 33505 34555 33563 34561
rect 28184 34524 28212 34552
rect 26896 34496 28212 34524
rect 26789 34459 26847 34465
rect 26789 34425 26801 34459
rect 26835 34425 26847 34459
rect 26789 34419 26847 34425
rect 26896 34388 26924 34496
rect 31478 34484 31484 34536
rect 31536 34524 31542 34536
rect 32217 34527 32275 34533
rect 32217 34524 32229 34527
rect 31536 34496 32229 34524
rect 31536 34484 31542 34496
rect 32217 34493 32229 34496
rect 32263 34493 32275 34527
rect 33336 34524 33364 34555
rect 33594 34552 33600 34564
rect 33652 34552 33658 34604
rect 33781 34595 33839 34601
rect 33781 34561 33793 34595
rect 33827 34592 33839 34595
rect 34054 34592 34060 34604
rect 33827 34564 34060 34592
rect 33827 34561 33839 34564
rect 33781 34555 33839 34561
rect 33796 34524 33824 34555
rect 34054 34552 34060 34564
rect 34112 34552 34118 34604
rect 35805 34595 35863 34601
rect 35805 34561 35817 34595
rect 35851 34592 35863 34595
rect 36464 34592 36492 34691
rect 38654 34688 38660 34700
rect 38712 34688 38718 34740
rect 39758 34688 39764 34740
rect 39816 34728 39822 34740
rect 41417 34731 41475 34737
rect 39816 34700 40724 34728
rect 39816 34688 39822 34700
rect 36725 34663 36783 34669
rect 36725 34660 36737 34663
rect 36556 34632 36737 34660
rect 36556 34604 36584 34632
rect 36725 34629 36737 34632
rect 36771 34660 36783 34663
rect 37366 34660 37372 34672
rect 36771 34632 37372 34660
rect 36771 34629 36783 34632
rect 36725 34623 36783 34629
rect 37366 34620 37372 34632
rect 37424 34620 37430 34672
rect 38838 34660 38844 34672
rect 38672 34632 38844 34660
rect 35851 34564 36492 34592
rect 35851 34561 35863 34564
rect 35805 34555 35863 34561
rect 36538 34552 36544 34604
rect 36596 34552 36602 34604
rect 36633 34595 36691 34601
rect 36633 34561 36645 34595
rect 36679 34561 36691 34595
rect 36633 34555 36691 34561
rect 33336 34496 33824 34524
rect 32217 34487 32275 34493
rect 34514 34484 34520 34536
rect 34572 34524 34578 34536
rect 36648 34524 36676 34555
rect 36814 34552 36820 34604
rect 36872 34552 36878 34604
rect 37001 34595 37059 34601
rect 37001 34561 37013 34595
rect 37047 34592 37059 34595
rect 37918 34592 37924 34604
rect 37047 34564 37924 34592
rect 37047 34561 37059 34564
rect 37001 34555 37059 34561
rect 37918 34552 37924 34564
rect 37976 34552 37982 34604
rect 38286 34552 38292 34604
rect 38344 34592 38350 34604
rect 38381 34595 38439 34601
rect 38381 34592 38393 34595
rect 38344 34564 38393 34592
rect 38344 34552 38350 34564
rect 38381 34561 38393 34564
rect 38427 34561 38439 34595
rect 38381 34555 38439 34561
rect 38470 34552 38476 34604
rect 38528 34552 38534 34604
rect 34572 34496 36676 34524
rect 34572 34484 34578 34496
rect 37090 34484 37096 34536
rect 37148 34524 37154 34536
rect 38672 34533 38700 34632
rect 38838 34620 38844 34632
rect 38896 34620 38902 34672
rect 40586 34660 40592 34672
rect 40342 34632 40592 34660
rect 40586 34620 40592 34632
rect 40644 34620 40650 34672
rect 40696 34660 40724 34700
rect 41417 34697 41429 34731
rect 41463 34728 41475 34731
rect 41506 34728 41512 34740
rect 41463 34700 41512 34728
rect 41463 34697 41475 34700
rect 41417 34691 41475 34697
rect 41506 34688 41512 34700
rect 41564 34688 41570 34740
rect 41690 34688 41696 34740
rect 41748 34728 41754 34740
rect 42705 34731 42763 34737
rect 41748 34700 41920 34728
rect 41748 34688 41754 34700
rect 40696 34632 41736 34660
rect 38746 34552 38752 34604
rect 38804 34552 38810 34604
rect 40512 34564 41414 34592
rect 37461 34527 37519 34533
rect 37461 34524 37473 34527
rect 37148 34496 37473 34524
rect 37148 34484 37154 34496
rect 37461 34493 37473 34496
rect 37507 34493 37519 34527
rect 38657 34527 38715 34533
rect 38657 34524 38669 34527
rect 37461 34487 37519 34493
rect 38212 34496 38669 34524
rect 36998 34416 37004 34468
rect 37056 34456 37062 34468
rect 38212 34456 38240 34496
rect 38657 34493 38669 34496
rect 38703 34493 38715 34527
rect 38657 34487 38715 34493
rect 38841 34527 38899 34533
rect 38841 34493 38853 34527
rect 38887 34493 38899 34527
rect 38841 34487 38899 34493
rect 37056 34428 38240 34456
rect 37056 34416 37062 34428
rect 38378 34416 38384 34468
rect 38436 34456 38442 34468
rect 38856 34456 38884 34487
rect 39114 34484 39120 34536
rect 39172 34484 39178 34536
rect 39574 34484 39580 34536
rect 39632 34524 39638 34536
rect 40512 34524 40540 34564
rect 39632 34496 40540 34524
rect 40589 34527 40647 34533
rect 39632 34484 39638 34496
rect 40589 34493 40601 34527
rect 40635 34524 40647 34527
rect 41233 34527 41291 34533
rect 41233 34524 41245 34527
rect 40635 34496 41245 34524
rect 40635 34493 40647 34496
rect 40589 34487 40647 34493
rect 41233 34493 41245 34496
rect 41279 34493 41291 34527
rect 41386 34524 41414 34564
rect 41598 34552 41604 34604
rect 41656 34552 41662 34604
rect 41708 34601 41736 34632
rect 41693 34595 41751 34601
rect 41693 34561 41705 34595
rect 41739 34561 41751 34595
rect 41693 34555 41751 34561
rect 41892 34533 41920 34700
rect 42705 34697 42717 34731
rect 42751 34728 42763 34731
rect 42751 34700 43116 34728
rect 42751 34697 42763 34700
rect 42705 34691 42763 34697
rect 43088 34669 43116 34700
rect 43073 34663 43131 34669
rect 43073 34629 43085 34663
rect 43119 34629 43131 34663
rect 43073 34623 43131 34629
rect 43530 34620 43536 34672
rect 43588 34620 43594 34672
rect 41966 34552 41972 34604
rect 42024 34552 42030 34604
rect 42518 34552 42524 34604
rect 42576 34552 42582 34604
rect 41877 34527 41935 34533
rect 41877 34524 41889 34527
rect 41386 34496 41889 34524
rect 41233 34487 41291 34493
rect 41877 34493 41889 34496
rect 41923 34493 41935 34527
rect 41877 34487 41935 34493
rect 42794 34484 42800 34536
rect 42852 34484 42858 34536
rect 43070 34484 43076 34536
rect 43128 34524 43134 34536
rect 44821 34527 44879 34533
rect 44821 34524 44833 34527
rect 43128 34496 44833 34524
rect 43128 34484 43134 34496
rect 44821 34493 44833 34496
rect 44867 34493 44879 34527
rect 44821 34487 44879 34493
rect 38436 34428 38884 34456
rect 38436 34416 38442 34428
rect 26712 34360 26924 34388
rect 23477 34351 23535 34357
rect 32582 34348 32588 34400
rect 32640 34388 32646 34400
rect 33318 34388 33324 34400
rect 32640 34360 33324 34388
rect 32640 34348 32646 34360
rect 33318 34348 33324 34360
rect 33376 34348 33382 34400
rect 38102 34348 38108 34400
rect 38160 34348 38166 34400
rect 38856 34388 38884 34428
rect 40402 34388 40408 34400
rect 38856 34360 40408 34388
rect 40402 34348 40408 34360
rect 40460 34348 40466 34400
rect 40678 34348 40684 34400
rect 40736 34348 40742 34400
rect 40770 34348 40776 34400
rect 40828 34388 40834 34400
rect 43530 34388 43536 34400
rect 40828 34360 43536 34388
rect 40828 34348 40834 34360
rect 43530 34348 43536 34360
rect 43588 34348 43594 34400
rect 1104 34298 45172 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 45172 34298
rect 1104 34224 45172 34246
rect 5166 34144 5172 34196
rect 5224 34144 5230 34196
rect 8481 34187 8539 34193
rect 8481 34153 8493 34187
rect 8527 34184 8539 34187
rect 8846 34184 8852 34196
rect 8527 34156 8852 34184
rect 8527 34153 8539 34156
rect 8481 34147 8539 34153
rect 8846 34144 8852 34156
rect 8904 34144 8910 34196
rect 12621 34187 12679 34193
rect 12621 34153 12633 34187
rect 12667 34184 12679 34187
rect 13633 34187 13691 34193
rect 12667 34156 12940 34184
rect 12667 34153 12679 34156
rect 12621 34147 12679 34153
rect 8938 34008 8944 34060
rect 8996 34008 9002 34060
rect 12434 34008 12440 34060
rect 12492 34008 12498 34060
rect 12912 33992 12940 34156
rect 13633 34153 13645 34187
rect 13679 34184 13691 34187
rect 13722 34184 13728 34196
rect 13679 34156 13728 34184
rect 13679 34153 13691 34156
rect 13633 34147 13691 34153
rect 13722 34144 13728 34156
rect 13780 34144 13786 34196
rect 14550 34144 14556 34196
rect 14608 34144 14614 34196
rect 14642 34144 14648 34196
rect 14700 34144 14706 34196
rect 14737 34187 14795 34193
rect 14737 34153 14749 34187
rect 14783 34184 14795 34187
rect 15654 34184 15660 34196
rect 14783 34156 15660 34184
rect 14783 34153 14795 34156
rect 14737 34147 14795 34153
rect 15654 34144 15660 34156
rect 15712 34144 15718 34196
rect 15746 34144 15752 34196
rect 15804 34144 15810 34196
rect 16022 34144 16028 34196
rect 16080 34144 16086 34196
rect 16666 34144 16672 34196
rect 16724 34184 16730 34196
rect 17957 34187 18015 34193
rect 17957 34184 17969 34187
rect 16724 34156 17969 34184
rect 16724 34144 16730 34156
rect 17957 34153 17969 34156
rect 18003 34153 18015 34187
rect 17957 34147 18015 34153
rect 20254 34144 20260 34196
rect 20312 34184 20318 34196
rect 20993 34187 21051 34193
rect 20993 34184 21005 34187
rect 20312 34156 21005 34184
rect 20312 34144 20318 34156
rect 20993 34153 21005 34156
rect 21039 34153 21051 34187
rect 20993 34147 21051 34153
rect 22002 34144 22008 34196
rect 22060 34184 22066 34196
rect 22060 34156 22416 34184
rect 22060 34144 22066 34156
rect 13357 34119 13415 34125
rect 13357 34085 13369 34119
rect 13403 34116 13415 34119
rect 14568 34116 14596 34144
rect 13403 34088 14596 34116
rect 14921 34119 14979 34125
rect 13403 34085 13415 34088
rect 13357 34079 13415 34085
rect 14921 34085 14933 34119
rect 14967 34116 14979 34119
rect 16040 34116 16068 34144
rect 14967 34088 16068 34116
rect 16301 34119 16359 34125
rect 14967 34085 14979 34088
rect 14921 34079 14979 34085
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 14384 34020 14749 34048
rect 14384 33992 14412 34020
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 3234 33940 3240 33992
rect 3292 33940 3298 33992
rect 3789 33983 3847 33989
rect 3789 33949 3801 33983
rect 3835 33980 3847 33983
rect 5166 33980 5172 33992
rect 3835 33952 5172 33980
rect 3835 33949 3847 33952
rect 3789 33943 3847 33949
rect 4172 33924 4200 33952
rect 5166 33940 5172 33952
rect 5224 33940 5230 33992
rect 5718 33940 5724 33992
rect 5776 33940 5782 33992
rect 7098 33940 7104 33992
rect 7156 33940 7162 33992
rect 7374 33989 7380 33992
rect 7368 33980 7380 33989
rect 7335 33952 7380 33980
rect 7368 33943 7380 33952
rect 7374 33940 7380 33943
rect 7432 33940 7438 33992
rect 8754 33940 8760 33992
rect 8812 33940 8818 33992
rect 10781 33983 10839 33989
rect 10781 33980 10793 33983
rect 10704 33952 10793 33980
rect 3878 33872 3884 33924
rect 3936 33912 3942 33924
rect 4034 33915 4092 33921
rect 4034 33912 4046 33915
rect 3936 33884 4046 33912
rect 3936 33872 3942 33884
rect 4034 33881 4046 33884
rect 4080 33881 4092 33915
rect 4034 33875 4092 33881
rect 4154 33872 4160 33924
rect 4212 33872 4218 33924
rect 8772 33912 8800 33940
rect 9217 33915 9275 33921
rect 9217 33912 9229 33915
rect 8772 33884 9229 33912
rect 9217 33881 9229 33884
rect 9263 33881 9275 33915
rect 9217 33875 9275 33881
rect 9950 33872 9956 33924
rect 10008 33872 10014 33924
rect 2406 33804 2412 33856
rect 2464 33844 2470 33856
rect 2685 33847 2743 33853
rect 2685 33844 2697 33847
rect 2464 33816 2697 33844
rect 2464 33804 2470 33816
rect 2685 33813 2697 33816
rect 2731 33813 2743 33847
rect 2685 33807 2743 33813
rect 6086 33804 6092 33856
rect 6144 33844 6150 33856
rect 6365 33847 6423 33853
rect 6365 33844 6377 33847
rect 6144 33816 6377 33844
rect 6144 33804 6150 33816
rect 6365 33813 6377 33816
rect 6411 33813 6423 33847
rect 6365 33807 6423 33813
rect 9122 33804 9128 33856
rect 9180 33844 9186 33856
rect 10704 33853 10732 33952
rect 10781 33949 10793 33952
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 12713 33983 12771 33989
rect 12713 33949 12725 33983
rect 12759 33949 12771 33983
rect 12713 33943 12771 33949
rect 10870 33872 10876 33924
rect 10928 33912 10934 33924
rect 11241 33915 11299 33921
rect 11241 33912 11253 33915
rect 10928 33884 11253 33912
rect 10928 33872 10934 33884
rect 11241 33881 11253 33884
rect 11287 33881 11299 33915
rect 11241 33875 11299 33881
rect 11425 33915 11483 33921
rect 11425 33881 11437 33915
rect 11471 33881 11483 33915
rect 12728 33912 12756 33943
rect 12894 33940 12900 33992
rect 12952 33989 12958 33992
rect 12952 33983 12988 33989
rect 12976 33949 12988 33983
rect 12952 33943 12988 33949
rect 12952 33940 12958 33943
rect 13354 33940 13360 33992
rect 13412 33980 13418 33992
rect 13449 33983 13507 33989
rect 13449 33980 13461 33983
rect 13412 33952 13461 33980
rect 13412 33940 13418 33952
rect 13449 33949 13461 33952
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 13538 33940 13544 33992
rect 13596 33980 13602 33992
rect 13722 33980 13728 33992
rect 13596 33952 13728 33980
rect 13596 33940 13602 33952
rect 13722 33940 13728 33952
rect 13780 33940 13786 33992
rect 14366 33940 14372 33992
rect 14424 33940 14430 33992
rect 14458 33940 14464 33992
rect 14516 33980 14522 33992
rect 14553 33983 14611 33989
rect 14553 33980 14565 33983
rect 14516 33952 14565 33980
rect 14516 33940 14522 33952
rect 14553 33949 14565 33952
rect 14599 33949 14611 33983
rect 14752 33980 14780 34011
rect 15212 33989 15240 34088
rect 16301 34085 16313 34119
rect 16347 34116 16359 34119
rect 18325 34119 18383 34125
rect 18325 34116 18337 34119
rect 16347 34088 17448 34116
rect 16347 34085 16359 34088
rect 16301 34079 16359 34085
rect 17420 34057 17448 34088
rect 17687 34088 18337 34116
rect 16945 34051 17003 34057
rect 16945 34048 16957 34051
rect 15672 34020 16957 34048
rect 15672 33989 15700 34020
rect 16945 34017 16957 34020
rect 16991 34017 17003 34051
rect 16945 34011 17003 34017
rect 17405 34051 17463 34057
rect 17405 34017 17417 34051
rect 17451 34017 17463 34051
rect 17405 34011 17463 34017
rect 15013 33983 15071 33989
rect 15013 33980 15025 33983
rect 14752 33952 15025 33980
rect 14553 33943 14611 33949
rect 15013 33949 15025 33952
rect 15059 33949 15071 33983
rect 15013 33943 15071 33949
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33949 15255 33983
rect 15197 33943 15255 33949
rect 15657 33983 15715 33989
rect 15657 33949 15669 33983
rect 15703 33949 15715 33983
rect 15657 33943 15715 33949
rect 16022 33940 16028 33992
rect 16080 33940 16086 33992
rect 16114 33940 16120 33992
rect 16172 33940 16178 33992
rect 16206 33940 16212 33992
rect 16264 33980 16270 33992
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 16264 33952 17049 33980
rect 16264 33940 16270 33952
rect 17037 33949 17049 33952
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 17126 33940 17132 33992
rect 17184 33940 17190 33992
rect 17310 33940 17316 33992
rect 17368 33980 17374 33992
rect 17687 33980 17715 34088
rect 18325 34085 18337 34088
rect 18371 34085 18383 34119
rect 21361 34119 21419 34125
rect 21361 34116 21373 34119
rect 18325 34079 18383 34085
rect 20640 34088 21373 34116
rect 17368 33952 17715 33980
rect 17368 33940 17374 33952
rect 18046 33940 18052 33992
rect 18104 33940 18110 33992
rect 18322 33940 18328 33992
rect 18380 33940 18386 33992
rect 19242 33940 19248 33992
rect 19300 33940 19306 33992
rect 20640 33966 20668 34088
rect 21361 34085 21373 34088
rect 21407 34116 21419 34119
rect 22278 34116 22284 34128
rect 21407 34088 22284 34116
rect 21407 34085 21419 34088
rect 21361 34079 21419 34085
rect 22278 34076 22284 34088
rect 22336 34076 22342 34128
rect 22094 34008 22100 34060
rect 22152 34008 22158 34060
rect 22189 34051 22247 34057
rect 22189 34017 22201 34051
rect 22235 34048 22247 34051
rect 22388 34048 22416 34156
rect 29362 34144 29368 34196
rect 29420 34184 29426 34196
rect 33042 34184 33048 34196
rect 29420 34156 33048 34184
rect 29420 34144 29426 34156
rect 33042 34144 33048 34156
rect 33100 34144 33106 34196
rect 33229 34187 33287 34193
rect 33229 34153 33241 34187
rect 33275 34184 33287 34187
rect 33318 34184 33324 34196
rect 33275 34156 33324 34184
rect 33275 34153 33287 34156
rect 33229 34147 33287 34153
rect 33318 34144 33324 34156
rect 33376 34184 33382 34196
rect 33686 34184 33692 34196
rect 33376 34156 33692 34184
rect 33376 34144 33382 34156
rect 33686 34144 33692 34156
rect 33744 34144 33750 34196
rect 33870 34144 33876 34196
rect 33928 34144 33934 34196
rect 34054 34144 34060 34196
rect 34112 34144 34118 34196
rect 36998 34144 37004 34196
rect 37056 34184 37062 34196
rect 37093 34187 37151 34193
rect 37093 34184 37105 34187
rect 37056 34156 37105 34184
rect 37056 34144 37062 34156
rect 37093 34153 37105 34156
rect 37139 34153 37151 34187
rect 37093 34147 37151 34153
rect 39393 34187 39451 34193
rect 39393 34153 39405 34187
rect 39439 34184 39451 34187
rect 40034 34184 40040 34196
rect 39439 34156 40040 34184
rect 39439 34153 39451 34156
rect 39393 34147 39451 34153
rect 40034 34144 40040 34156
rect 40092 34144 40098 34196
rect 42518 34144 42524 34196
rect 42576 34184 42582 34196
rect 42613 34187 42671 34193
rect 42613 34184 42625 34187
rect 42576 34156 42625 34184
rect 42576 34144 42582 34156
rect 42613 34153 42625 34156
rect 42659 34153 42671 34187
rect 42613 34147 42671 34153
rect 42794 34144 42800 34196
rect 42852 34144 42858 34196
rect 33888 34116 33916 34144
rect 32968 34088 33916 34116
rect 32968 34048 32996 34088
rect 22235 34020 22416 34048
rect 31726 34020 32996 34048
rect 22235 34017 22247 34020
rect 22189 34011 22247 34017
rect 23474 33980 23480 33992
rect 21100 33952 23480 33980
rect 13814 33912 13820 33924
rect 12728 33884 13820 33912
rect 11425 33875 11483 33881
rect 10689 33847 10747 33853
rect 10689 33844 10701 33847
rect 9180 33816 10701 33844
rect 9180 33804 9186 33816
rect 10689 33813 10701 33816
rect 10735 33813 10747 33847
rect 10689 33807 10747 33813
rect 10962 33804 10968 33856
rect 11020 33844 11026 33856
rect 11440 33844 11468 33875
rect 11020 33816 11468 33844
rect 11020 33804 11026 33816
rect 11606 33804 11612 33856
rect 11664 33804 11670 33856
rect 11882 33804 11888 33856
rect 11940 33844 11946 33856
rect 12161 33847 12219 33853
rect 12161 33844 12173 33847
rect 11940 33816 12173 33844
rect 11940 33804 11946 33816
rect 12161 33813 12173 33816
rect 12207 33813 12219 33847
rect 12161 33807 12219 33813
rect 12802 33804 12808 33856
rect 12860 33804 12866 33856
rect 13004 33853 13032 33884
rect 13814 33872 13820 33884
rect 13872 33872 13878 33924
rect 15105 33915 15163 33921
rect 15105 33881 15117 33915
rect 15151 33912 15163 33915
rect 15746 33912 15752 33924
rect 15151 33884 15752 33912
rect 15151 33881 15163 33884
rect 15105 33875 15163 33881
rect 15746 33872 15752 33884
rect 15804 33912 15810 33924
rect 16393 33915 16451 33921
rect 16393 33912 16405 33915
rect 15804 33884 16405 33912
rect 15804 33872 15810 33884
rect 16393 33881 16405 33884
rect 16439 33881 16451 33915
rect 16393 33875 16451 33881
rect 16669 33915 16727 33921
rect 16669 33881 16681 33915
rect 16715 33912 16727 33915
rect 17218 33912 17224 33924
rect 16715 33884 17224 33912
rect 16715 33881 16727 33884
rect 16669 33875 16727 33881
rect 17218 33872 17224 33884
rect 17276 33872 17282 33924
rect 17497 33915 17555 33921
rect 17497 33881 17509 33915
rect 17543 33881 17555 33915
rect 17497 33875 17555 33881
rect 12989 33847 13047 33853
rect 12989 33813 13001 33847
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 15010 33804 15016 33856
rect 15068 33844 15074 33856
rect 16577 33847 16635 33853
rect 16577 33844 16589 33847
rect 15068 33816 16589 33844
rect 15068 33804 15074 33816
rect 16577 33813 16589 33816
rect 16623 33813 16635 33847
rect 16577 33807 16635 33813
rect 16761 33847 16819 33853
rect 16761 33813 16773 33847
rect 16807 33844 16819 33847
rect 16850 33844 16856 33856
rect 16807 33816 16856 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 16850 33804 16856 33816
rect 16908 33804 16914 33856
rect 17512 33844 17540 33875
rect 17586 33872 17592 33924
rect 17644 33872 17650 33924
rect 17678 33872 17684 33924
rect 17736 33912 17742 33924
rect 17773 33915 17831 33921
rect 17773 33912 17785 33915
rect 17736 33884 17785 33912
rect 17736 33872 17742 33884
rect 17773 33881 17785 33884
rect 17819 33881 17831 33915
rect 19521 33915 19579 33921
rect 17773 33875 17831 33881
rect 17880 33884 19472 33912
rect 17880 33844 17908 33884
rect 17512 33816 17908 33844
rect 18138 33804 18144 33856
rect 18196 33804 18202 33856
rect 19444 33844 19472 33884
rect 19521 33881 19533 33915
rect 19567 33912 19579 33915
rect 19610 33912 19616 33924
rect 19567 33884 19616 33912
rect 19567 33881 19579 33884
rect 19521 33875 19579 33881
rect 19610 33872 19616 33884
rect 19668 33872 19674 33924
rect 21100 33844 21128 33952
rect 23474 33940 23480 33952
rect 23532 33940 23538 33992
rect 24578 33940 24584 33992
rect 24636 33940 24642 33992
rect 27982 33940 27988 33992
rect 28040 33980 28046 33992
rect 28718 33980 28724 33992
rect 28040 33952 28724 33980
rect 28040 33940 28046 33952
rect 28718 33940 28724 33952
rect 28776 33980 28782 33992
rect 29273 33983 29331 33989
rect 29273 33980 29285 33983
rect 28776 33952 29285 33980
rect 28776 33940 28782 33952
rect 29273 33949 29285 33952
rect 29319 33980 29331 33983
rect 31205 33983 31263 33989
rect 31205 33980 31217 33983
rect 29319 33952 31217 33980
rect 29319 33949 29331 33952
rect 29273 33943 29331 33949
rect 31205 33949 31217 33952
rect 31251 33980 31263 33983
rect 31726 33980 31754 34020
rect 33042 34008 33048 34060
rect 33100 34008 33106 34060
rect 33226 34008 33232 34060
rect 33284 34048 33290 34060
rect 37274 34048 37280 34060
rect 33284 34020 33364 34048
rect 33284 34008 33290 34020
rect 32953 33983 33011 33989
rect 32953 33980 32965 33983
rect 31251 33952 31754 33980
rect 32876 33952 32965 33980
rect 31251 33949 31263 33952
rect 31205 33943 31263 33949
rect 32876 33924 32904 33952
rect 32953 33949 32965 33952
rect 32999 33949 33011 33983
rect 32953 33943 33011 33949
rect 33134 33940 33140 33992
rect 33192 33940 33198 33992
rect 33336 33989 33364 34020
rect 36924 34020 37280 34048
rect 33321 33983 33379 33989
rect 33321 33949 33333 33983
rect 33367 33949 33379 33983
rect 33321 33943 33379 33949
rect 33410 33940 33416 33992
rect 33468 33940 33474 33992
rect 33594 33940 33600 33992
rect 33652 33940 33658 33992
rect 33962 33940 33968 33992
rect 34020 33940 34026 33992
rect 36924 33989 36952 34020
rect 37274 34008 37280 34020
rect 37332 34008 37338 34060
rect 37642 34008 37648 34060
rect 37700 34048 37706 34060
rect 38378 34048 38384 34060
rect 37700 34020 38384 34048
rect 37700 34008 37706 34020
rect 38378 34008 38384 34020
rect 38436 34008 38442 34060
rect 40770 34048 40776 34060
rect 39040 34020 40776 34048
rect 39040 33992 39068 34020
rect 40770 34008 40776 34020
rect 40828 34008 40834 34060
rect 41322 34008 41328 34060
rect 41380 34048 41386 34060
rect 41969 34051 42027 34057
rect 41969 34048 41981 34051
rect 41380 34020 41981 34048
rect 41380 34008 41386 34020
rect 41969 34017 41981 34020
rect 42015 34017 42027 34051
rect 41969 34011 42027 34017
rect 42705 34051 42763 34057
rect 42705 34017 42717 34051
rect 42751 34048 42763 34051
rect 42812 34048 42840 34144
rect 42751 34020 42840 34048
rect 42751 34017 42763 34020
rect 42705 34011 42763 34017
rect 35989 33983 36047 33989
rect 35989 33949 36001 33983
rect 36035 33980 36047 33983
rect 36633 33983 36691 33989
rect 36633 33980 36645 33983
rect 36035 33952 36645 33980
rect 36035 33949 36047 33952
rect 35989 33943 36047 33949
rect 36633 33949 36645 33952
rect 36679 33949 36691 33983
rect 36633 33943 36691 33949
rect 36817 33983 36875 33989
rect 36817 33949 36829 33983
rect 36863 33949 36875 33983
rect 36817 33943 36875 33949
rect 36909 33983 36967 33989
rect 36909 33949 36921 33983
rect 36955 33949 36967 33983
rect 36909 33943 36967 33949
rect 21174 33872 21180 33924
rect 21232 33872 21238 33924
rect 32858 33872 32864 33924
rect 32916 33872 32922 33924
rect 33152 33912 33180 33940
rect 35161 33915 35219 33921
rect 35161 33912 35173 33915
rect 33152 33884 35173 33912
rect 35161 33881 35173 33884
rect 35207 33881 35219 33915
rect 35161 33875 35219 33881
rect 19444 33816 21128 33844
rect 21634 33804 21640 33856
rect 21692 33804 21698 33856
rect 22002 33804 22008 33856
rect 22060 33804 22066 33856
rect 24765 33847 24823 33853
rect 24765 33813 24777 33847
rect 24811 33844 24823 33847
rect 25222 33844 25228 33856
rect 24811 33816 25228 33844
rect 24811 33813 24823 33816
rect 24765 33807 24823 33813
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 27522 33804 27528 33856
rect 27580 33844 27586 33856
rect 27801 33847 27859 33853
rect 27801 33844 27813 33847
rect 27580 33816 27813 33844
rect 27580 33804 27586 33816
rect 27801 33813 27813 33816
rect 27847 33813 27859 33847
rect 27801 33807 27859 33813
rect 33045 33847 33103 33853
rect 33045 33813 33057 33847
rect 33091 33844 33103 33847
rect 33134 33844 33140 33856
rect 33091 33816 33140 33844
rect 33091 33813 33103 33816
rect 33045 33807 33103 33813
rect 33134 33804 33140 33816
rect 33192 33804 33198 33856
rect 33410 33804 33416 33856
rect 33468 33804 33474 33856
rect 35437 33847 35495 33853
rect 35437 33813 35449 33847
rect 35483 33844 35495 33847
rect 35894 33844 35900 33856
rect 35483 33816 35900 33844
rect 35483 33813 35495 33816
rect 35437 33807 35495 33813
rect 35894 33804 35900 33816
rect 35952 33804 35958 33856
rect 36541 33847 36599 33853
rect 36541 33813 36553 33847
rect 36587 33844 36599 33847
rect 36630 33844 36636 33856
rect 36587 33816 36636 33844
rect 36587 33813 36599 33816
rect 36541 33807 36599 33813
rect 36630 33804 36636 33816
rect 36688 33804 36694 33856
rect 36832 33844 36860 33943
rect 36998 33940 37004 33992
rect 37056 33980 37062 33992
rect 37185 33983 37243 33989
rect 37185 33980 37197 33983
rect 37056 33952 37197 33980
rect 37056 33940 37062 33952
rect 37185 33949 37197 33952
rect 37231 33949 37243 33983
rect 37185 33943 37243 33949
rect 39022 33940 39028 33992
rect 39080 33940 39086 33992
rect 40402 33940 40408 33992
rect 40460 33980 40466 33992
rect 41601 33983 41659 33989
rect 41601 33980 41613 33983
rect 40460 33952 41613 33980
rect 40460 33940 40466 33952
rect 41601 33949 41613 33952
rect 41647 33980 41659 33983
rect 42720 33980 42748 34011
rect 41647 33952 42748 33980
rect 41647 33949 41659 33952
rect 41601 33943 41659 33949
rect 37921 33915 37979 33921
rect 37921 33881 37933 33915
rect 37967 33912 37979 33915
rect 38010 33912 38016 33924
rect 37967 33884 38016 33912
rect 37967 33881 37979 33884
rect 37921 33875 37979 33881
rect 38010 33872 38016 33884
rect 38068 33872 38074 33924
rect 39853 33915 39911 33921
rect 39853 33881 39865 33915
rect 39899 33912 39911 33915
rect 39942 33912 39948 33924
rect 39899 33884 39948 33912
rect 39899 33881 39911 33884
rect 39853 33875 39911 33881
rect 39942 33872 39948 33884
rect 40000 33872 40006 33924
rect 41966 33872 41972 33924
rect 42024 33912 42030 33924
rect 42153 33915 42211 33921
rect 42153 33912 42165 33915
rect 42024 33884 42165 33912
rect 42024 33872 42030 33884
rect 42153 33881 42165 33884
rect 42199 33881 42211 33915
rect 42153 33875 42211 33881
rect 42978 33872 42984 33924
rect 43036 33872 43042 33924
rect 43070 33872 43076 33924
rect 43128 33872 43134 33924
rect 43438 33872 43444 33924
rect 43496 33872 43502 33924
rect 37274 33844 37280 33856
rect 36832 33816 37280 33844
rect 37274 33804 37280 33816
rect 37332 33844 37338 33856
rect 38286 33844 38292 33856
rect 37332 33816 38292 33844
rect 37332 33804 37338 33816
rect 38286 33804 38292 33816
rect 38344 33804 38350 33856
rect 38838 33804 38844 33856
rect 38896 33844 38902 33856
rect 39574 33844 39580 33856
rect 38896 33816 39580 33844
rect 38896 33804 38902 33816
rect 39574 33804 39580 33816
rect 39632 33804 39638 33856
rect 42245 33847 42303 33853
rect 42245 33813 42257 33847
rect 42291 33844 42303 33847
rect 43088 33844 43116 33872
rect 42291 33816 43116 33844
rect 42291 33813 42303 33816
rect 42245 33807 42303 33813
rect 43622 33804 43628 33856
rect 43680 33844 43686 33856
rect 44453 33847 44511 33853
rect 44453 33844 44465 33847
rect 43680 33816 44465 33844
rect 43680 33804 43686 33816
rect 44453 33813 44465 33816
rect 44499 33813 44511 33847
rect 44453 33807 44511 33813
rect 1104 33754 45172 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 45172 33754
rect 1104 33680 45172 33702
rect 3329 33643 3387 33649
rect 3329 33609 3341 33643
rect 3375 33609 3387 33643
rect 3329 33603 3387 33609
rect 2992 33575 3050 33581
rect 2992 33541 3004 33575
rect 3038 33572 3050 33575
rect 3344 33572 3372 33603
rect 3878 33600 3884 33652
rect 3936 33600 3942 33652
rect 3973 33643 4031 33649
rect 3973 33609 3985 33643
rect 4019 33609 4031 33643
rect 3973 33603 4031 33609
rect 4341 33643 4399 33649
rect 4341 33609 4353 33643
rect 4387 33640 4399 33643
rect 4798 33640 4804 33652
rect 4387 33612 4804 33640
rect 4387 33609 4399 33612
rect 4341 33603 4399 33609
rect 3038 33544 3372 33572
rect 3038 33541 3050 33544
rect 2992 33535 3050 33541
rect 3510 33464 3516 33516
rect 3568 33464 3574 33516
rect 3697 33507 3755 33513
rect 3697 33473 3709 33507
rect 3743 33504 3755 33507
rect 3988 33504 4016 33603
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 5074 33600 5080 33652
rect 5132 33600 5138 33652
rect 5537 33643 5595 33649
rect 5537 33609 5549 33643
rect 5583 33640 5595 33643
rect 5718 33640 5724 33652
rect 5583 33612 5724 33640
rect 5583 33609 5595 33612
rect 5537 33603 5595 33609
rect 5718 33600 5724 33612
rect 5776 33600 5782 33652
rect 7558 33600 7564 33652
rect 7616 33600 7622 33652
rect 8570 33600 8576 33652
rect 8628 33640 8634 33652
rect 8757 33643 8815 33649
rect 8757 33640 8769 33643
rect 8628 33612 8769 33640
rect 8628 33600 8634 33612
rect 8757 33609 8769 33612
rect 8803 33609 8815 33643
rect 8757 33603 8815 33609
rect 9122 33600 9128 33652
rect 9180 33600 9186 33652
rect 9217 33643 9275 33649
rect 9217 33609 9229 33643
rect 9263 33640 9275 33643
rect 9490 33640 9496 33652
rect 9263 33612 9496 33640
rect 9263 33609 9275 33612
rect 9217 33603 9275 33609
rect 5626 33572 5632 33584
rect 5000 33544 5632 33572
rect 3743 33476 4016 33504
rect 3743 33473 3755 33476
rect 3697 33467 3755 33473
rect 4154 33464 4160 33516
rect 4212 33464 4218 33516
rect 3237 33439 3295 33445
rect 3237 33405 3249 33439
rect 3283 33436 3295 33439
rect 4172 33436 4200 33464
rect 3283 33408 4200 33436
rect 4433 33439 4491 33445
rect 3283 33405 3295 33408
rect 3237 33399 3295 33405
rect 4433 33405 4445 33439
rect 4479 33405 4491 33439
rect 4433 33399 4491 33405
rect 1857 33303 1915 33309
rect 1857 33269 1869 33303
rect 1903 33300 1915 33303
rect 2498 33300 2504 33312
rect 1903 33272 2504 33300
rect 1903 33269 1915 33272
rect 1857 33263 1915 33269
rect 2498 33260 2504 33272
rect 2556 33260 2562 33312
rect 2590 33260 2596 33312
rect 2648 33300 2654 33312
rect 3252 33300 3280 33399
rect 4448 33368 4476 33399
rect 4614 33396 4620 33448
rect 4672 33396 4678 33448
rect 5000 33445 5028 33544
rect 5626 33532 5632 33544
rect 5684 33572 5690 33584
rect 7929 33575 7987 33581
rect 5684 33544 7880 33572
rect 5684 33532 5690 33544
rect 5169 33507 5227 33513
rect 5169 33473 5181 33507
rect 5215 33473 5227 33507
rect 5169 33467 5227 33473
rect 5813 33507 5871 33513
rect 5813 33473 5825 33507
rect 5859 33504 5871 33507
rect 6086 33504 6092 33516
rect 5859 33476 6092 33504
rect 5859 33473 5871 33476
rect 5813 33467 5871 33473
rect 4985 33439 5043 33445
rect 4985 33405 4997 33439
rect 5031 33405 5043 33439
rect 5184 33436 5212 33467
rect 6086 33464 6092 33476
rect 6144 33464 6150 33516
rect 6914 33464 6920 33516
rect 6972 33504 6978 33516
rect 7101 33507 7159 33513
rect 7101 33504 7113 33507
rect 6972 33476 7113 33504
rect 6972 33464 6978 33476
rect 7101 33473 7113 33476
rect 7147 33473 7159 33507
rect 7852 33504 7880 33544
rect 7929 33541 7941 33575
rect 7975 33572 7987 33575
rect 9232 33572 9260 33603
rect 9490 33600 9496 33612
rect 9548 33600 9554 33652
rect 10870 33600 10876 33652
rect 10928 33600 10934 33652
rect 11238 33600 11244 33652
rect 11296 33600 11302 33652
rect 12158 33600 12164 33652
rect 12216 33600 12222 33652
rect 12802 33600 12808 33652
rect 12860 33600 12866 33652
rect 14550 33640 14556 33652
rect 13832 33612 14556 33640
rect 7975 33544 9260 33572
rect 10781 33575 10839 33581
rect 7975 33541 7987 33544
rect 7929 33535 7987 33541
rect 10781 33541 10793 33575
rect 10827 33572 10839 33575
rect 10888 33572 10916 33600
rect 10827 33544 10916 33572
rect 10827 33541 10839 33544
rect 10781 33535 10839 33541
rect 7852 33476 8156 33504
rect 7101 33467 7159 33473
rect 5184 33408 6316 33436
rect 4985 33399 5043 33405
rect 5534 33368 5540 33380
rect 4448 33340 5540 33368
rect 5534 33328 5540 33340
rect 5592 33328 5598 33380
rect 6288 33368 6316 33408
rect 6362 33396 6368 33448
rect 6420 33396 6426 33448
rect 8018 33396 8024 33448
rect 8076 33396 8082 33448
rect 8128 33445 8156 33476
rect 11054 33464 11060 33516
rect 11112 33504 11118 33516
rect 11256 33504 11284 33600
rect 11112 33476 11284 33504
rect 11112 33464 11118 33476
rect 11606 33464 11612 33516
rect 11664 33464 11670 33516
rect 11698 33464 11704 33516
rect 11756 33464 11762 33516
rect 11882 33513 11888 33516
rect 11839 33507 11888 33513
rect 11839 33473 11851 33507
rect 11885 33473 11888 33507
rect 11839 33467 11888 33473
rect 11882 33464 11888 33467
rect 11940 33464 11946 33516
rect 12161 33507 12219 33513
rect 12161 33473 12173 33507
rect 12207 33504 12219 33507
rect 12820 33504 12848 33600
rect 12207 33476 12848 33504
rect 13832 33502 13860 33612
rect 14550 33600 14556 33612
rect 14608 33600 14614 33652
rect 14921 33643 14979 33649
rect 14921 33609 14933 33643
rect 14967 33609 14979 33643
rect 14921 33603 14979 33609
rect 14093 33575 14151 33581
rect 14093 33541 14105 33575
rect 14139 33572 14151 33575
rect 14139 33544 14596 33572
rect 14139 33541 14151 33544
rect 14093 33535 14151 33541
rect 14001 33507 14059 33513
rect 14001 33502 14013 33507
rect 12207 33473 12219 33476
rect 13832 33474 14013 33502
rect 12161 33467 12219 33473
rect 14001 33473 14013 33474
rect 14047 33473 14059 33507
rect 14001 33467 14059 33473
rect 14185 33507 14243 33513
rect 14185 33473 14197 33507
rect 14231 33504 14243 33507
rect 14458 33504 14464 33516
rect 14231 33476 14464 33504
rect 14231 33473 14243 33476
rect 14185 33467 14243 33473
rect 14458 33464 14464 33476
rect 14516 33464 14522 33516
rect 14568 33504 14596 33544
rect 14642 33532 14648 33584
rect 14700 33532 14706 33584
rect 14936 33572 14964 33603
rect 16022 33600 16028 33652
rect 16080 33640 16086 33652
rect 16669 33643 16727 33649
rect 16669 33640 16681 33643
rect 16080 33612 16681 33640
rect 16080 33600 16086 33612
rect 16669 33609 16681 33612
rect 16715 33609 16727 33643
rect 16669 33603 16727 33609
rect 16850 33600 16856 33652
rect 16908 33600 16914 33652
rect 17218 33600 17224 33652
rect 17276 33640 17282 33652
rect 17497 33643 17555 33649
rect 17497 33640 17509 33643
rect 17276 33612 17509 33640
rect 17276 33600 17282 33612
rect 17497 33609 17509 33612
rect 17543 33609 17555 33643
rect 18046 33640 18052 33652
rect 17497 33603 17555 33609
rect 17972 33612 18052 33640
rect 16868 33572 16896 33600
rect 14936 33544 16896 33572
rect 17310 33532 17316 33584
rect 17368 33532 17374 33584
rect 14918 33504 14924 33516
rect 14568 33476 14924 33504
rect 14918 33464 14924 33476
rect 14976 33464 14982 33516
rect 16206 33504 16212 33516
rect 15488 33476 16212 33504
rect 8113 33439 8171 33445
rect 8113 33405 8125 33439
rect 8159 33405 8171 33439
rect 8113 33399 8171 33405
rect 9398 33396 9404 33448
rect 9456 33396 9462 33448
rect 10594 33396 10600 33448
rect 10652 33436 10658 33448
rect 10689 33439 10747 33445
rect 10689 33436 10701 33439
rect 10652 33408 10701 33436
rect 10652 33396 10658 33408
rect 10689 33405 10701 33408
rect 10735 33436 10747 33439
rect 10962 33436 10968 33448
rect 10735 33408 10968 33436
rect 10735 33405 10747 33408
rect 10689 33399 10747 33405
rect 10962 33396 10968 33408
rect 11020 33396 11026 33448
rect 11149 33439 11207 33445
rect 11149 33405 11161 33439
rect 11195 33436 11207 33439
rect 11238 33436 11244 33448
rect 11195 33408 11244 33436
rect 11195 33405 11207 33408
rect 11149 33399 11207 33405
rect 11238 33396 11244 33408
rect 11296 33396 11302 33448
rect 11624 33436 11652 33464
rect 15080 33439 15138 33445
rect 15080 33436 15092 33439
rect 11624 33408 15092 33436
rect 6822 33368 6828 33380
rect 6288 33340 6828 33368
rect 6822 33328 6828 33340
rect 6880 33368 6886 33380
rect 7009 33371 7067 33377
rect 7009 33368 7021 33371
rect 6880 33340 7021 33368
rect 6880 33328 6886 33340
rect 7009 33337 7021 33340
rect 7055 33337 7067 33371
rect 7009 33331 7067 33337
rect 11333 33371 11391 33377
rect 11333 33337 11345 33371
rect 11379 33368 11391 33371
rect 11379 33340 12572 33368
rect 11379 33337 11391 33340
rect 11333 33331 11391 33337
rect 2648 33272 3280 33300
rect 2648 33260 2654 33272
rect 5626 33260 5632 33312
rect 5684 33260 5690 33312
rect 7193 33303 7251 33309
rect 7193 33269 7205 33303
rect 7239 33300 7251 33303
rect 9582 33300 9588 33312
rect 7239 33272 9588 33300
rect 7239 33269 7251 33272
rect 7193 33263 7251 33269
rect 9582 33260 9588 33272
rect 9640 33260 9646 33312
rect 11974 33260 11980 33312
rect 12032 33260 12038 33312
rect 12544 33300 12572 33340
rect 14274 33328 14280 33380
rect 14332 33328 14338 33380
rect 14090 33300 14096 33312
rect 12544 33272 14096 33300
rect 14090 33260 14096 33272
rect 14148 33260 14154 33312
rect 14651 33309 14679 33408
rect 15080 33405 15092 33408
rect 15126 33405 15138 33439
rect 15080 33399 15138 33405
rect 15194 33396 15200 33448
rect 15252 33396 15258 33448
rect 15286 33396 15292 33448
rect 15344 33396 15350 33448
rect 14829 33371 14887 33377
rect 14829 33337 14841 33371
rect 14875 33368 14887 33371
rect 15488 33368 15516 33476
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 16390 33464 16396 33516
rect 16448 33464 16454 33516
rect 16482 33464 16488 33516
rect 16540 33504 16546 33516
rect 16853 33507 16911 33513
rect 16853 33504 16865 33507
rect 16540 33476 16865 33504
rect 16540 33464 16546 33476
rect 16853 33473 16865 33476
rect 16899 33473 16911 33507
rect 16853 33467 16911 33473
rect 17681 33507 17739 33513
rect 17681 33473 17693 33507
rect 17727 33473 17739 33507
rect 17681 33467 17739 33473
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33436 15623 33439
rect 16298 33436 16304 33448
rect 15611 33408 16304 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 17037 33439 17095 33445
rect 17037 33405 17049 33439
rect 17083 33405 17095 33439
rect 17696 33436 17724 33467
rect 17770 33464 17776 33516
rect 17828 33464 17834 33516
rect 17696 33408 17908 33436
rect 17037 33399 17095 33405
rect 14875 33340 15516 33368
rect 17052 33368 17080 33399
rect 17678 33368 17684 33380
rect 17052 33340 17684 33368
rect 14875 33337 14887 33340
rect 14829 33331 14887 33337
rect 17678 33328 17684 33340
rect 17736 33328 17742 33380
rect 14645 33303 14703 33309
rect 14645 33269 14657 33303
rect 14691 33269 14703 33303
rect 14645 33263 14703 33269
rect 15838 33260 15844 33312
rect 15896 33260 15902 33312
rect 15930 33260 15936 33312
rect 15988 33300 15994 33312
rect 16853 33303 16911 33309
rect 16853 33300 16865 33303
rect 15988 33272 16865 33300
rect 15988 33260 15994 33272
rect 16853 33269 16865 33272
rect 16899 33269 16911 33303
rect 17880 33300 17908 33408
rect 17972 33377 18000 33612
rect 18046 33600 18052 33612
rect 18104 33600 18110 33652
rect 19889 33643 19947 33649
rect 19889 33609 19901 33643
rect 19935 33640 19947 33643
rect 20070 33640 20076 33652
rect 19935 33612 20076 33640
rect 19935 33609 19947 33612
rect 19889 33603 19947 33609
rect 20070 33600 20076 33612
rect 20128 33600 20134 33652
rect 21634 33600 21640 33652
rect 21692 33600 21698 33652
rect 24394 33600 24400 33652
rect 24452 33640 24458 33652
rect 25038 33640 25044 33652
rect 24452 33612 25044 33640
rect 24452 33600 24458 33612
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 25222 33600 25228 33652
rect 25280 33640 25286 33652
rect 25280 33612 25912 33640
rect 25280 33600 25286 33612
rect 21542 33572 21548 33584
rect 18156 33544 21548 33572
rect 18156 33516 18184 33544
rect 21542 33532 21548 33544
rect 21600 33532 21606 33584
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33504 18107 33507
rect 18138 33504 18144 33516
rect 18095 33476 18144 33504
rect 18095 33473 18107 33476
rect 18049 33467 18107 33473
rect 18138 33464 18144 33476
rect 18196 33464 18202 33516
rect 18877 33507 18935 33513
rect 18877 33473 18889 33507
rect 18923 33504 18935 33507
rect 20165 33507 20223 33513
rect 18923 33476 19564 33504
rect 18923 33473 18935 33476
rect 18877 33467 18935 33473
rect 18892 33436 18920 33467
rect 18064 33408 18920 33436
rect 17957 33371 18015 33377
rect 17957 33337 17969 33371
rect 18003 33337 18015 33371
rect 17957 33331 18015 33337
rect 18064 33300 18092 33408
rect 19150 33396 19156 33448
rect 19208 33436 19214 33448
rect 19245 33439 19303 33445
rect 19245 33436 19257 33439
rect 19208 33408 19257 33436
rect 19208 33396 19214 33408
rect 19245 33405 19257 33408
rect 19291 33405 19303 33439
rect 19536 33436 19564 33476
rect 20165 33473 20177 33507
rect 20211 33504 20223 33507
rect 20254 33504 20260 33516
rect 20211 33476 20260 33504
rect 20211 33473 20223 33476
rect 20165 33467 20223 33473
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 21453 33507 21511 33513
rect 21453 33473 21465 33507
rect 21499 33504 21511 33507
rect 21652 33504 21680 33600
rect 23934 33532 23940 33584
rect 23992 33572 23998 33584
rect 25884 33581 25912 33612
rect 27522 33600 27528 33652
rect 27580 33640 27586 33652
rect 33781 33643 33839 33649
rect 27580 33612 29546 33640
rect 27580 33600 27586 33612
rect 24029 33575 24087 33581
rect 24029 33572 24041 33575
rect 23992 33544 24041 33572
rect 23992 33532 23998 33544
rect 24029 33541 24041 33544
rect 24075 33541 24087 33575
rect 24029 33535 24087 33541
rect 25869 33575 25927 33581
rect 25869 33541 25881 33575
rect 25915 33541 25927 33575
rect 25869 33535 25927 33541
rect 21499 33476 21680 33504
rect 24213 33507 24271 33513
rect 21499 33473 21511 33476
rect 21453 33467 21511 33473
rect 24213 33473 24225 33507
rect 24259 33504 24271 33507
rect 24762 33504 24768 33516
rect 24259 33476 24768 33504
rect 24259 33473 24271 33476
rect 24213 33467 24271 33473
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 26145 33507 26203 33513
rect 26145 33473 26157 33507
rect 26191 33504 26203 33507
rect 26326 33504 26332 33516
rect 26191 33476 26332 33504
rect 26191 33473 26203 33476
rect 26145 33467 26203 33473
rect 26326 33464 26332 33476
rect 26384 33504 26390 33516
rect 27540 33504 27568 33600
rect 26384 33476 27568 33504
rect 27617 33507 27675 33513
rect 26384 33464 26390 33476
rect 27617 33473 27629 33507
rect 27663 33504 27675 33507
rect 27706 33504 27712 33516
rect 27663 33476 27712 33504
rect 27663 33473 27675 33476
rect 27617 33467 27675 33473
rect 27706 33464 27712 33476
rect 27764 33464 27770 33516
rect 27908 33513 27936 33612
rect 27893 33507 27951 33513
rect 27893 33473 27905 33507
rect 27939 33473 27951 33507
rect 29518 33504 29546 33612
rect 33781 33609 33793 33643
rect 33827 33640 33839 33643
rect 33962 33640 33968 33652
rect 33827 33612 33968 33640
rect 33827 33609 33839 33612
rect 33781 33603 33839 33609
rect 30009 33507 30067 33513
rect 30009 33504 30021 33507
rect 27893 33467 27951 33473
rect 24670 33436 24676 33448
rect 19536 33408 24676 33436
rect 19245 33399 19303 33405
rect 24670 33396 24676 33408
rect 24728 33396 24734 33448
rect 28169 33439 28227 33445
rect 28169 33436 28181 33439
rect 27816 33408 28181 33436
rect 23934 33328 23940 33380
rect 23992 33328 23998 33380
rect 27816 33377 27844 33408
rect 28169 33405 28181 33408
rect 28215 33405 28227 33439
rect 29288 33436 29316 33490
rect 29518 33476 30021 33504
rect 30009 33473 30021 33476
rect 30055 33473 30067 33507
rect 33137 33507 33195 33513
rect 30009 33467 30067 33473
rect 29454 33436 29460 33448
rect 29288 33408 29460 33436
rect 28169 33399 28227 33405
rect 29454 33396 29460 33408
rect 29512 33436 29518 33448
rect 30285 33439 30343 33445
rect 29512 33408 29776 33436
rect 29512 33396 29518 33408
rect 27801 33371 27859 33377
rect 27801 33337 27813 33371
rect 27847 33337 27859 33371
rect 27801 33331 27859 33337
rect 17880 33272 18092 33300
rect 16853 33263 16911 33269
rect 18782 33260 18788 33312
rect 18840 33260 18846 33312
rect 18874 33260 18880 33312
rect 18932 33300 18938 33312
rect 20073 33303 20131 33309
rect 20073 33300 20085 33303
rect 18932 33272 20085 33300
rect 18932 33260 18938 33272
rect 20073 33269 20085 33272
rect 20119 33269 20131 33303
rect 20073 33263 20131 33269
rect 21266 33260 21272 33312
rect 21324 33260 21330 33312
rect 23952 33300 23980 33328
rect 29362 33300 29368 33312
rect 23952 33272 29368 33300
rect 29362 33260 29368 33272
rect 29420 33260 29426 33312
rect 29546 33260 29552 33312
rect 29604 33300 29610 33312
rect 29641 33303 29699 33309
rect 29641 33300 29653 33303
rect 29604 33272 29653 33300
rect 29604 33260 29610 33272
rect 29641 33269 29653 33272
rect 29687 33269 29699 33303
rect 29748 33300 29776 33408
rect 30285 33405 30297 33439
rect 30331 33436 30343 33439
rect 30742 33436 30748 33448
rect 30331 33408 30748 33436
rect 30331 33405 30343 33408
rect 30285 33399 30343 33405
rect 30742 33396 30748 33408
rect 30800 33396 30806 33448
rect 31404 33300 31432 33490
rect 33137 33473 33149 33507
rect 33183 33504 33195 33507
rect 33796 33504 33824 33603
rect 33962 33600 33968 33612
rect 34020 33600 34026 33652
rect 35526 33640 35532 33652
rect 35452 33612 35532 33640
rect 35452 33572 35480 33612
rect 35526 33600 35532 33612
rect 35584 33640 35590 33652
rect 35989 33643 36047 33649
rect 35989 33640 36001 33643
rect 35584 33612 36001 33640
rect 35584 33600 35590 33612
rect 35989 33609 36001 33612
rect 36035 33640 36047 33643
rect 40313 33643 40371 33649
rect 40313 33640 40325 33643
rect 36035 33612 38884 33640
rect 36035 33609 36047 33612
rect 35989 33603 36047 33609
rect 37182 33572 37188 33584
rect 34822 33544 35480 33572
rect 35544 33544 37188 33572
rect 35544 33513 35572 33544
rect 37182 33532 37188 33544
rect 37240 33572 37246 33584
rect 37642 33572 37648 33584
rect 37240 33544 37648 33572
rect 37240 33532 37246 33544
rect 33183 33476 33824 33504
rect 35529 33507 35587 33513
rect 33183 33473 33195 33476
rect 33137 33467 33195 33473
rect 35529 33473 35541 33507
rect 35575 33473 35587 33507
rect 35529 33467 35587 33473
rect 35713 33507 35771 33513
rect 35713 33473 35725 33507
rect 35759 33504 35771 33507
rect 35894 33504 35900 33516
rect 35759 33476 35900 33504
rect 35759 33473 35771 33476
rect 35713 33467 35771 33473
rect 35894 33464 35900 33476
rect 35952 33504 35958 33516
rect 36814 33504 36820 33516
rect 35952 33476 36820 33504
rect 35952 33464 35958 33476
rect 36814 33464 36820 33476
rect 36872 33464 36878 33516
rect 37292 33513 37320 33544
rect 37642 33532 37648 33544
rect 37700 33532 37706 33584
rect 38856 33572 38884 33612
rect 39224 33612 40325 33640
rect 39022 33572 39028 33584
rect 38778 33544 39028 33572
rect 39022 33532 39028 33544
rect 39080 33532 39086 33584
rect 37277 33507 37335 33513
rect 37277 33473 37289 33507
rect 37323 33473 37335 33507
rect 37277 33467 37335 33473
rect 38838 33464 38844 33516
rect 38896 33504 38902 33516
rect 39224 33513 39252 33612
rect 40313 33609 40325 33612
rect 40359 33640 40371 33643
rect 40678 33640 40684 33652
rect 40359 33612 40684 33640
rect 40359 33609 40371 33612
rect 40313 33603 40371 33609
rect 40678 33600 40684 33612
rect 40736 33600 40742 33652
rect 42886 33600 42892 33652
rect 42944 33600 42950 33652
rect 42978 33600 42984 33652
rect 43036 33640 43042 33652
rect 43441 33643 43499 33649
rect 43441 33640 43453 33643
rect 43036 33612 43453 33640
rect 43036 33600 43042 33612
rect 43441 33609 43453 33612
rect 43487 33609 43499 33643
rect 43441 33603 43499 33609
rect 43622 33600 43628 33652
rect 43680 33600 43686 33652
rect 43162 33572 43168 33584
rect 42996 33544 43168 33572
rect 39209 33507 39267 33513
rect 38896 33476 39160 33504
rect 38896 33464 38902 33476
rect 31754 33396 31760 33448
rect 31812 33436 31818 33448
rect 32677 33439 32735 33445
rect 32677 33436 32689 33439
rect 31812 33408 32689 33436
rect 31812 33396 31818 33408
rect 32677 33405 32689 33408
rect 32723 33405 32735 33439
rect 32677 33399 32735 33405
rect 34790 33396 34796 33448
rect 34848 33436 34854 33448
rect 35253 33439 35311 33445
rect 35253 33436 35265 33439
rect 34848 33408 35265 33436
rect 34848 33396 34854 33408
rect 35253 33405 35265 33408
rect 35299 33405 35311 33439
rect 35253 33399 35311 33405
rect 35986 33396 35992 33448
rect 36044 33436 36050 33448
rect 36449 33439 36507 33445
rect 36449 33436 36461 33439
rect 36044 33408 36461 33436
rect 36044 33396 36050 33408
rect 36449 33405 36461 33408
rect 36495 33405 36507 33439
rect 36449 33399 36507 33405
rect 37553 33439 37611 33445
rect 37553 33405 37565 33439
rect 37599 33436 37611 33439
rect 38102 33436 38108 33448
rect 37599 33408 38108 33436
rect 37599 33405 37611 33408
rect 37553 33399 37611 33405
rect 38102 33396 38108 33408
rect 38160 33396 38166 33448
rect 38286 33396 38292 33448
rect 38344 33436 38350 33448
rect 39132 33436 39160 33476
rect 39209 33473 39221 33507
rect 39255 33473 39267 33507
rect 39209 33467 39267 33473
rect 39482 33464 39488 33516
rect 39540 33464 39546 33516
rect 39577 33507 39635 33513
rect 39577 33473 39589 33507
rect 39623 33473 39635 33507
rect 39577 33467 39635 33473
rect 39301 33439 39359 33445
rect 39301 33436 39313 33439
rect 38344 33408 39068 33436
rect 39132 33408 39313 33436
rect 38344 33396 38350 33408
rect 33689 33371 33747 33377
rect 33689 33337 33701 33371
rect 33735 33368 33747 33371
rect 34054 33368 34060 33380
rect 33735 33340 34060 33368
rect 33735 33337 33747 33340
rect 33689 33331 33747 33337
rect 34054 33328 34060 33340
rect 34112 33328 34118 33380
rect 39040 33368 39068 33408
rect 39301 33405 39313 33408
rect 39347 33405 39359 33439
rect 39301 33399 39359 33405
rect 39592 33368 39620 33467
rect 40218 33464 40224 33516
rect 40276 33464 40282 33516
rect 40681 33507 40739 33513
rect 40681 33504 40693 33507
rect 40328 33476 40693 33504
rect 40328 33436 40356 33476
rect 40681 33473 40693 33476
rect 40727 33473 40739 33507
rect 41322 33504 41328 33516
rect 40681 33467 40739 33473
rect 41156 33476 41328 33504
rect 39040 33340 39620 33368
rect 39684 33408 40356 33436
rect 29748 33272 31432 33300
rect 29641 33263 29699 33269
rect 32122 33260 32128 33312
rect 32180 33260 32186 33312
rect 36538 33260 36544 33312
rect 36596 33300 36602 33312
rect 36998 33300 37004 33312
rect 36596 33272 37004 33300
rect 36596 33260 36602 33272
rect 36998 33260 37004 33272
rect 37056 33300 37062 33312
rect 37093 33303 37151 33309
rect 37093 33300 37105 33303
rect 37056 33272 37105 33300
rect 37056 33260 37062 33272
rect 37093 33269 37105 33272
rect 37139 33269 37151 33303
rect 37093 33263 37151 33269
rect 39022 33260 39028 33312
rect 39080 33260 39086 33312
rect 39206 33260 39212 33312
rect 39264 33300 39270 33312
rect 39684 33300 39712 33408
rect 40494 33396 40500 33448
rect 40552 33436 40558 33448
rect 41156 33436 41184 33476
rect 41322 33464 41328 33476
rect 41380 33504 41386 33516
rect 41380 33464 41414 33504
rect 42058 33464 42064 33516
rect 42116 33464 42122 33516
rect 42996 33513 43024 33544
rect 43162 33532 43168 33544
rect 43220 33572 43226 33584
rect 43640 33572 43668 33600
rect 43220 33544 43668 33572
rect 43220 33532 43226 33544
rect 42981 33507 43039 33513
rect 42981 33473 42993 33507
rect 43027 33473 43039 33507
rect 43625 33507 43683 33513
rect 43625 33504 43637 33507
rect 42981 33467 43039 33473
rect 43364 33476 43637 33504
rect 40552 33408 41184 33436
rect 41233 33439 41291 33445
rect 40552 33396 40558 33408
rect 41233 33405 41245 33439
rect 41279 33405 41291 33439
rect 41386 33436 41414 33464
rect 42705 33439 42763 33445
rect 42705 33436 42717 33439
rect 41386 33408 42717 33436
rect 41233 33399 41291 33405
rect 42705 33405 42717 33408
rect 42751 33436 42763 33439
rect 42886 33436 42892 33448
rect 42751 33408 42892 33436
rect 42751 33405 42763 33408
rect 42705 33399 42763 33405
rect 39761 33371 39819 33377
rect 39761 33337 39773 33371
rect 39807 33368 39819 33371
rect 41248 33368 41276 33399
rect 42886 33396 42892 33408
rect 42944 33396 42950 33448
rect 43364 33377 43392 33476
rect 43625 33473 43637 33476
rect 43671 33473 43683 33507
rect 43625 33467 43683 33473
rect 44266 33396 44272 33448
rect 44324 33436 44330 33448
rect 44361 33439 44419 33445
rect 44361 33436 44373 33439
rect 44324 33408 44373 33436
rect 44324 33396 44330 33408
rect 44361 33405 44373 33408
rect 44407 33405 44419 33439
rect 44361 33399 44419 33405
rect 39807 33340 41276 33368
rect 43349 33371 43407 33377
rect 39807 33337 39819 33340
rect 39761 33331 39819 33337
rect 43349 33337 43361 33371
rect 43395 33337 43407 33371
rect 43349 33331 43407 33337
rect 44082 33328 44088 33380
rect 44140 33328 44146 33380
rect 39264 33272 39712 33300
rect 39264 33260 39270 33272
rect 39850 33260 39856 33312
rect 39908 33260 39914 33312
rect 41506 33260 41512 33312
rect 41564 33260 41570 33312
rect 43898 33260 43904 33312
rect 43956 33260 43962 33312
rect 1104 33210 45172 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 45172 33210
rect 1104 33136 45172 33158
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 3605 33099 3663 33105
rect 3605 33096 3617 33099
rect 3568 33068 3617 33096
rect 3568 33056 3574 33068
rect 3605 33065 3617 33068
rect 3651 33065 3663 33099
rect 4614 33096 4620 33108
rect 3605 33059 3663 33065
rect 4448 33068 4620 33096
rect 2041 33031 2099 33037
rect 2041 32997 2053 33031
rect 2087 32997 2099 33031
rect 2041 32991 2099 32997
rect 1949 32895 2007 32901
rect 1949 32861 1961 32895
rect 1995 32892 2007 32895
rect 2056 32892 2084 32991
rect 2498 32920 2504 32972
rect 2556 32920 2562 32972
rect 2685 32963 2743 32969
rect 2685 32929 2697 32963
rect 2731 32960 2743 32963
rect 2866 32960 2872 32972
rect 2731 32932 2872 32960
rect 2731 32929 2743 32932
rect 2685 32923 2743 32929
rect 2866 32920 2872 32932
rect 2924 32920 2930 32972
rect 3053 32963 3111 32969
rect 3053 32929 3065 32963
rect 3099 32960 3111 32963
rect 4448 32960 4476 33068
rect 4614 33056 4620 33068
rect 4672 33096 4678 33108
rect 5813 33099 5871 33105
rect 4672 33068 5764 33096
rect 4672 33056 4678 33068
rect 3099 32932 4476 32960
rect 5736 32960 5764 33068
rect 5813 33065 5825 33099
rect 5859 33096 5871 33099
rect 6362 33096 6368 33108
rect 5859 33068 6368 33096
rect 5859 33065 5871 33068
rect 5813 33059 5871 33065
rect 6362 33056 6368 33068
rect 6420 33056 6426 33108
rect 7098 33096 7104 33108
rect 6748 33068 7104 33096
rect 6748 32969 6776 33068
rect 7098 33056 7104 33068
rect 7156 33056 7162 33108
rect 8110 33056 8116 33108
rect 8168 33056 8174 33108
rect 11793 33099 11851 33105
rect 9232 33068 11192 33096
rect 6733 32963 6791 32969
rect 5736 32932 6684 32960
rect 3099 32929 3111 32932
rect 3053 32923 3111 32929
rect 1995 32864 2084 32892
rect 1995 32861 2007 32864
rect 1949 32855 2007 32861
rect 2406 32852 2412 32904
rect 2464 32852 2470 32904
rect 2516 32824 2544 32920
rect 3237 32895 3295 32901
rect 3237 32892 3249 32895
rect 2746 32864 3249 32892
rect 2746 32824 2774 32864
rect 3237 32861 3249 32864
rect 3283 32892 3295 32895
rect 3694 32892 3700 32904
rect 3283 32864 3700 32892
rect 3283 32861 3295 32864
rect 3237 32855 3295 32861
rect 3694 32852 3700 32864
rect 3752 32852 3758 32904
rect 4433 32895 4491 32901
rect 4433 32861 4445 32895
rect 4479 32892 4491 32895
rect 5166 32892 5172 32904
rect 4479 32864 5172 32892
rect 4479 32861 4491 32864
rect 4433 32855 4491 32861
rect 5166 32852 5172 32864
rect 5224 32852 5230 32904
rect 5626 32852 5632 32904
rect 5684 32852 5690 32904
rect 6086 32852 6092 32904
rect 6144 32852 6150 32904
rect 6656 32892 6684 32932
rect 6733 32929 6745 32963
rect 6779 32929 6791 32963
rect 8128 32960 8156 33056
rect 9232 33040 9260 33068
rect 9214 32988 9220 33040
rect 9272 32988 9278 33040
rect 11054 32988 11060 33040
rect 11112 32988 11118 33040
rect 11164 33028 11192 33068
rect 11793 33065 11805 33099
rect 11839 33096 11851 33099
rect 11882 33096 11888 33108
rect 11839 33068 11888 33096
rect 11839 33065 11851 33068
rect 11793 33059 11851 33065
rect 11882 33056 11888 33068
rect 11940 33056 11946 33108
rect 11977 33099 12035 33105
rect 11977 33065 11989 33099
rect 12023 33096 12035 33099
rect 14274 33096 14280 33108
rect 12023 33068 14280 33096
rect 12023 33065 12035 33068
rect 11977 33059 12035 33065
rect 14274 33056 14280 33068
rect 14332 33056 14338 33108
rect 14642 33056 14648 33108
rect 14700 33096 14706 33108
rect 14829 33099 14887 33105
rect 14829 33096 14841 33099
rect 14700 33068 14841 33096
rect 14700 33056 14706 33068
rect 14829 33065 14841 33068
rect 14875 33065 14887 33099
rect 16482 33096 16488 33108
rect 14829 33059 14887 33065
rect 14937 33068 16488 33096
rect 12894 33028 12900 33040
rect 11164 33000 12900 33028
rect 12894 32988 12900 33000
rect 12952 33028 12958 33040
rect 13173 33031 13231 33037
rect 13173 33028 13185 33031
rect 12952 33000 13185 33028
rect 12952 32988 12958 33000
rect 13173 32997 13185 33000
rect 13219 32997 13231 33031
rect 14937 33028 14965 33068
rect 15194 33028 15200 33040
rect 13173 32991 13231 32997
rect 14108 33000 14965 33028
rect 15028 33000 15200 33028
rect 9493 32963 9551 32969
rect 9493 32960 9505 32963
rect 8128 32932 9505 32960
rect 6733 32923 6791 32929
rect 9493 32929 9505 32932
rect 9539 32929 9551 32963
rect 9493 32923 9551 32929
rect 10060 32932 11008 32960
rect 10060 32904 10088 32932
rect 7282 32892 7288 32904
rect 6656 32864 7288 32892
rect 7282 32852 7288 32864
rect 7340 32852 7346 32904
rect 8018 32852 8024 32904
rect 8076 32892 8082 32904
rect 8941 32895 8999 32901
rect 8941 32892 8953 32895
rect 8076 32864 8953 32892
rect 8076 32852 8082 32864
rect 8941 32861 8953 32864
rect 8987 32861 8999 32895
rect 8941 32855 8999 32861
rect 10042 32852 10048 32904
rect 10100 32852 10106 32904
rect 10980 32901 11008 32932
rect 10781 32895 10839 32901
rect 10781 32892 10793 32895
rect 10244 32864 10793 32892
rect 4700 32827 4758 32833
rect 2516 32796 2774 32824
rect 3160 32796 4660 32824
rect 1762 32716 1768 32768
rect 1820 32716 1826 32768
rect 3160 32765 3188 32796
rect 3145 32759 3203 32765
rect 3145 32725 3157 32759
rect 3191 32725 3203 32759
rect 4632 32756 4660 32796
rect 4700 32793 4712 32827
rect 4746 32824 4758 32827
rect 5644 32824 5672 32852
rect 4746 32796 5672 32824
rect 7000 32827 7058 32833
rect 4746 32793 4758 32796
rect 4700 32787 4758 32793
rect 7000 32793 7012 32827
rect 7046 32824 7058 32827
rect 7190 32824 7196 32836
rect 7046 32796 7196 32824
rect 7046 32793 7058 32796
rect 7000 32787 7058 32793
rect 7190 32784 7196 32796
rect 7248 32784 7254 32836
rect 10244 32768 10272 32864
rect 10781 32861 10793 32864
rect 10827 32861 10839 32895
rect 10781 32855 10839 32861
rect 10965 32895 11023 32901
rect 10965 32861 10977 32895
rect 11011 32861 11023 32895
rect 11072 32892 11100 32988
rect 14108 32972 14136 33000
rect 11149 32963 11207 32969
rect 11149 32929 11161 32963
rect 11195 32960 11207 32963
rect 11698 32960 11704 32972
rect 11195 32932 11704 32960
rect 11195 32929 11207 32932
rect 11149 32923 11207 32929
rect 11698 32920 11704 32932
rect 11756 32920 11762 32972
rect 13538 32960 13544 32972
rect 12912 32932 13544 32960
rect 11241 32895 11299 32901
rect 11241 32892 11253 32895
rect 11072 32864 11253 32892
rect 10965 32855 11023 32861
rect 11241 32861 11253 32864
rect 11287 32861 11299 32895
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 11241 32855 11299 32861
rect 11348 32864 11437 32892
rect 11348 32824 11376 32864
rect 11425 32861 11437 32864
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11606 32852 11612 32904
rect 11664 32852 11670 32904
rect 12912 32901 12940 32932
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 14090 32920 14096 32972
rect 14148 32920 14154 32972
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 12986 32852 12992 32904
rect 13044 32852 13050 32904
rect 13265 32895 13323 32901
rect 13265 32861 13277 32895
rect 13311 32892 13323 32895
rect 13722 32892 13728 32904
rect 13311 32864 13728 32892
rect 13311 32861 13323 32864
rect 13265 32855 13323 32861
rect 13722 32852 13728 32864
rect 13780 32892 13786 32904
rect 14458 32892 14464 32904
rect 13780 32864 14464 32892
rect 13780 32852 13786 32864
rect 14458 32852 14464 32864
rect 14516 32852 14522 32904
rect 15028 32901 15056 33000
rect 15194 32988 15200 33000
rect 15252 32988 15258 33040
rect 15102 32920 15108 32972
rect 15160 32920 15166 32972
rect 15304 32969 15332 33068
rect 16482 33056 16488 33068
rect 16540 33056 16546 33108
rect 16758 33056 16764 33108
rect 16816 33056 16822 33108
rect 17678 33056 17684 33108
rect 17736 33096 17742 33108
rect 17865 33099 17923 33105
rect 17865 33096 17877 33099
rect 17736 33068 17877 33096
rect 17736 33056 17742 33068
rect 17865 33065 17877 33068
rect 17911 33065 17923 33099
rect 17865 33059 17923 33065
rect 18414 33056 18420 33108
rect 18472 33056 18478 33108
rect 24578 33056 24584 33108
rect 24636 33096 24642 33108
rect 24673 33099 24731 33105
rect 24673 33096 24685 33099
rect 24636 33068 24685 33096
rect 24636 33056 24642 33068
rect 24673 33065 24685 33068
rect 24719 33065 24731 33099
rect 24673 33059 24731 33065
rect 24762 33056 24768 33108
rect 24820 33096 24826 33108
rect 24820 33068 27660 33096
rect 24820 33056 24826 33068
rect 27632 33028 27660 33068
rect 27706 33056 27712 33108
rect 27764 33096 27770 33108
rect 28169 33099 28227 33105
rect 28169 33096 28181 33099
rect 27764 33068 28181 33096
rect 27764 33056 27770 33068
rect 28169 33065 28181 33068
rect 28215 33065 28227 33099
rect 28169 33059 28227 33065
rect 28902 33056 28908 33108
rect 28960 33096 28966 33108
rect 30193 33099 30251 33105
rect 30193 33096 30205 33099
rect 28960 33068 30205 33096
rect 28960 33056 28966 33068
rect 30193 33065 30205 33068
rect 30239 33065 30251 33099
rect 30193 33059 30251 33065
rect 30282 33056 30288 33108
rect 30340 33096 30346 33108
rect 30561 33099 30619 33105
rect 30561 33096 30573 33099
rect 30340 33068 30573 33096
rect 30340 33056 30346 33068
rect 30561 33065 30573 33068
rect 30607 33065 30619 33099
rect 30561 33059 30619 33065
rect 30742 33056 30748 33108
rect 30800 33096 30806 33108
rect 31205 33099 31263 33105
rect 31205 33096 31217 33099
rect 30800 33068 31217 33096
rect 30800 33056 30806 33068
rect 31205 33065 31217 33068
rect 31251 33065 31263 33099
rect 31205 33059 31263 33065
rect 31938 33056 31944 33108
rect 31996 33096 32002 33108
rect 32674 33096 32680 33108
rect 31996 33068 32680 33096
rect 31996 33056 32002 33068
rect 32674 33056 32680 33068
rect 32732 33056 32738 33108
rect 34333 33099 34391 33105
rect 34333 33065 34345 33099
rect 34379 33096 34391 33099
rect 34790 33096 34796 33108
rect 34379 33068 34796 33096
rect 34379 33065 34391 33068
rect 34333 33059 34391 33065
rect 34790 33056 34796 33068
rect 34848 33056 34854 33108
rect 35253 33099 35311 33105
rect 35253 33065 35265 33099
rect 35299 33096 35311 33099
rect 35986 33096 35992 33108
rect 35299 33068 35992 33096
rect 35299 33065 35311 33068
rect 35253 33059 35311 33065
rect 35986 33056 35992 33068
rect 36044 33056 36050 33108
rect 36906 33056 36912 33108
rect 36964 33056 36970 33108
rect 37090 33056 37096 33108
rect 37148 33056 37154 33108
rect 39850 33096 39856 33108
rect 39500 33068 39856 33096
rect 29454 33028 29460 33040
rect 15580 33000 19104 33028
rect 15289 32963 15347 32969
rect 15289 32929 15301 32963
rect 15335 32929 15347 32963
rect 15289 32923 15347 32929
rect 15013 32895 15071 32901
rect 15013 32861 15025 32895
rect 15059 32861 15071 32895
rect 15013 32855 15071 32861
rect 15028 32824 15056 32855
rect 15194 32852 15200 32904
rect 15252 32852 15258 32904
rect 15470 32852 15476 32904
rect 15528 32852 15534 32904
rect 11256 32796 11376 32824
rect 11440 32796 15056 32824
rect 11256 32768 11284 32796
rect 5718 32756 5724 32768
rect 4632 32728 5724 32756
rect 3145 32719 3203 32725
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 5902 32716 5908 32768
rect 5960 32716 5966 32768
rect 10226 32716 10232 32768
rect 10284 32716 10290 32768
rect 11238 32716 11244 32768
rect 11296 32716 11302 32768
rect 11440 32765 11468 32796
rect 15102 32784 15108 32836
rect 15160 32824 15166 32836
rect 15580 32824 15608 33000
rect 18708 32932 19012 32960
rect 16206 32852 16212 32904
rect 16264 32892 16270 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 16264 32864 17325 32892
rect 16264 32852 16270 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17589 32895 17647 32901
rect 17589 32892 17601 32895
rect 17313 32855 17371 32861
rect 17420 32864 17601 32892
rect 15160 32796 15608 32824
rect 15160 32784 15166 32796
rect 17126 32784 17132 32836
rect 17184 32824 17190 32836
rect 17420 32824 17448 32864
rect 17589 32861 17601 32864
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 17681 32895 17739 32901
rect 17681 32861 17693 32895
rect 17727 32892 17739 32895
rect 17862 32892 17868 32904
rect 17727 32864 17868 32892
rect 17727 32861 17739 32864
rect 17681 32855 17739 32861
rect 17862 32852 17868 32864
rect 17920 32852 17926 32904
rect 18708 32901 18736 32932
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32861 18751 32895
rect 18693 32855 18751 32861
rect 18874 32852 18880 32904
rect 18932 32852 18938 32904
rect 17184 32796 17448 32824
rect 17497 32827 17555 32833
rect 17184 32784 17190 32796
rect 17497 32793 17509 32827
rect 17543 32824 17555 32827
rect 18892 32824 18920 32852
rect 17543 32796 18920 32824
rect 17543 32793 17555 32796
rect 17497 32787 17555 32793
rect 11425 32759 11483 32765
rect 11425 32725 11437 32759
rect 11471 32725 11483 32759
rect 11425 32719 11483 32725
rect 12710 32716 12716 32768
rect 12768 32716 12774 32768
rect 13262 32716 13268 32768
rect 13320 32756 13326 32768
rect 13630 32756 13636 32768
rect 13320 32728 13636 32756
rect 13320 32716 13326 32728
rect 13630 32716 13636 32728
rect 13688 32716 13694 32768
rect 17402 32716 17408 32768
rect 17460 32756 17466 32768
rect 17512 32756 17540 32787
rect 18984 32768 19012 32932
rect 19076 32836 19104 33000
rect 25976 33000 26464 33028
rect 27632 33000 29460 33028
rect 19242 32920 19248 32972
rect 19300 32960 19306 32972
rect 20717 32963 20775 32969
rect 20717 32960 20729 32963
rect 19300 32932 20729 32960
rect 19300 32920 19306 32932
rect 20717 32929 20729 32932
rect 20763 32960 20775 32963
rect 20990 32960 20996 32972
rect 20763 32932 20996 32960
rect 20763 32929 20775 32932
rect 20717 32923 20775 32929
rect 20990 32920 20996 32932
rect 21048 32920 21054 32972
rect 24486 32920 24492 32972
rect 24544 32960 24550 32972
rect 25225 32963 25283 32969
rect 25225 32960 25237 32963
rect 24544 32932 25237 32960
rect 24544 32920 24550 32932
rect 25225 32929 25237 32932
rect 25271 32929 25283 32963
rect 25225 32923 25283 32929
rect 23474 32852 23480 32904
rect 23532 32892 23538 32904
rect 23845 32895 23903 32901
rect 23845 32892 23857 32895
rect 23532 32864 23857 32892
rect 23532 32852 23538 32864
rect 23845 32861 23857 32864
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 25038 32852 25044 32904
rect 25096 32852 25102 32904
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32892 25191 32895
rect 25976 32892 26004 33000
rect 26326 32920 26332 32972
rect 26384 32920 26390 32972
rect 26436 32960 26464 33000
rect 26602 32960 26608 32972
rect 26436 32932 26608 32960
rect 26602 32920 26608 32932
rect 26660 32920 26666 32972
rect 25179 32864 26004 32892
rect 25179 32861 25191 32864
rect 25133 32855 25191 32861
rect 26050 32852 26056 32904
rect 26108 32852 26114 32904
rect 27724 32878 27752 33000
rect 29454 32988 29460 33000
rect 29512 32988 29518 33040
rect 30098 32988 30104 33040
rect 30156 32988 30162 33040
rect 31021 33031 31079 33037
rect 31021 32997 31033 33031
rect 31067 33028 31079 33031
rect 31067 33000 32260 33028
rect 31067 32997 31079 33000
rect 31021 32991 31079 32997
rect 28810 32920 28816 32972
rect 28868 32920 28874 32972
rect 29638 32920 29644 32972
rect 29696 32920 29702 32972
rect 30285 32963 30343 32969
rect 30285 32960 30297 32963
rect 29748 32932 30297 32960
rect 29748 32901 29776 32932
rect 30285 32929 30297 32932
rect 30331 32929 30343 32963
rect 31754 32960 31760 32972
rect 30285 32923 30343 32929
rect 31128 32932 31760 32960
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 28092 32864 29745 32892
rect 19058 32784 19064 32836
rect 19116 32784 19122 32836
rect 20993 32827 21051 32833
rect 20993 32793 21005 32827
rect 21039 32824 21051 32827
rect 21266 32824 21272 32836
rect 21039 32796 21272 32824
rect 21039 32793 21051 32796
rect 20993 32787 21051 32793
rect 21266 32784 21272 32796
rect 21324 32784 21330 32836
rect 22278 32824 22284 32836
rect 22218 32796 22284 32824
rect 22278 32784 22284 32796
rect 22336 32784 22342 32836
rect 24213 32827 24271 32833
rect 24213 32793 24225 32827
rect 24259 32824 24271 32827
rect 24578 32824 24584 32836
rect 24259 32796 24584 32824
rect 24259 32793 24271 32796
rect 24213 32787 24271 32793
rect 24578 32784 24584 32796
rect 24636 32784 24642 32836
rect 26605 32827 26663 32833
rect 26605 32824 26617 32827
rect 26252 32796 26617 32824
rect 17460 32728 17540 32756
rect 17460 32716 17466 32728
rect 18230 32716 18236 32768
rect 18288 32716 18294 32768
rect 18966 32716 18972 32768
rect 19024 32756 19030 32768
rect 22002 32756 22008 32768
rect 19024 32728 22008 32756
rect 19024 32716 19030 32728
rect 22002 32716 22008 32728
rect 22060 32756 22066 32768
rect 26252 32765 26280 32796
rect 26605 32793 26617 32796
rect 26651 32793 26663 32827
rect 26605 32787 26663 32793
rect 22465 32759 22523 32765
rect 22465 32756 22477 32759
rect 22060 32728 22477 32756
rect 22060 32716 22066 32728
rect 22465 32725 22477 32728
rect 22511 32725 22523 32759
rect 22465 32719 22523 32725
rect 26237 32759 26295 32765
rect 26237 32725 26249 32759
rect 26283 32725 26295 32759
rect 26237 32719 26295 32725
rect 27338 32716 27344 32768
rect 27396 32756 27402 32768
rect 28092 32765 28120 32864
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 30926 32852 30932 32904
rect 30984 32852 30990 32904
rect 31128 32901 31156 32932
rect 31754 32920 31760 32932
rect 31812 32920 31818 32972
rect 31849 32963 31907 32969
rect 31849 32929 31861 32963
rect 31895 32960 31907 32963
rect 32122 32960 32128 32972
rect 31895 32932 32128 32960
rect 31895 32929 31907 32932
rect 31849 32923 31907 32929
rect 32122 32920 32128 32932
rect 32180 32920 32186 32972
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32861 31171 32895
rect 31113 32855 31171 32861
rect 31386 32852 31392 32904
rect 31444 32852 31450 32904
rect 31478 32852 31484 32904
rect 31536 32852 31542 32904
rect 31573 32895 31631 32901
rect 31573 32861 31585 32895
rect 31619 32892 31631 32895
rect 31938 32892 31944 32904
rect 31619 32864 31944 32892
rect 31619 32861 31631 32864
rect 31573 32855 31631 32861
rect 31938 32852 31944 32864
rect 31996 32852 32002 32904
rect 32232 32892 32260 33000
rect 32950 32988 32956 33040
rect 33008 32988 33014 33040
rect 33042 32988 33048 33040
rect 33100 32988 33106 33040
rect 33686 33028 33692 33040
rect 33236 33000 33692 33028
rect 32490 32920 32496 32972
rect 32548 32960 32554 32972
rect 32968 32960 32996 32988
rect 32548 32932 32996 32960
rect 33133 32963 33191 32969
rect 32548 32920 32554 32932
rect 33133 32929 33145 32963
rect 33179 32960 33191 32963
rect 33236 32960 33264 33000
rect 33686 32988 33692 33000
rect 33744 32988 33750 33040
rect 35526 32988 35532 33040
rect 35584 32988 35590 33040
rect 36924 33028 36952 33056
rect 37553 33031 37611 33037
rect 37553 33028 37565 33031
rect 36924 33000 37565 33028
rect 37553 32997 37565 33000
rect 37599 32997 37611 33031
rect 37553 32991 37611 32997
rect 33179 32932 33264 32960
rect 33179 32929 33191 32932
rect 33133 32923 33191 32929
rect 33318 32920 33324 32972
rect 33376 32920 33382 32972
rect 32585 32895 32643 32901
rect 32585 32892 32597 32895
rect 32232 32864 32597 32892
rect 32585 32861 32597 32864
rect 32631 32861 32643 32895
rect 32585 32855 32643 32861
rect 32769 32895 32827 32901
rect 32769 32861 32781 32895
rect 32815 32892 32827 32895
rect 32953 32895 33011 32901
rect 32953 32894 32965 32895
rect 32876 32892 32965 32894
rect 32815 32866 32965 32892
rect 32815 32864 32904 32866
rect 32815 32861 32827 32864
rect 32769 32855 32827 32861
rect 32953 32861 32965 32866
rect 32999 32861 33011 32895
rect 32953 32855 33011 32861
rect 28537 32827 28595 32833
rect 28537 32793 28549 32827
rect 28583 32824 28595 32827
rect 29546 32824 29552 32836
rect 28583 32796 29552 32824
rect 28583 32793 28595 32796
rect 28537 32787 28595 32793
rect 29546 32784 29552 32796
rect 29604 32784 29610 32836
rect 31662 32784 31668 32836
rect 31720 32833 31726 32836
rect 31720 32827 31769 32833
rect 31720 32793 31723 32827
rect 31757 32824 31769 32827
rect 32600 32824 32628 32855
rect 33226 32852 33232 32904
rect 33284 32852 33290 32904
rect 33336 32824 33364 32920
rect 33502 32852 33508 32904
rect 33560 32852 33566 32904
rect 33778 32852 33784 32904
rect 33836 32852 33842 32904
rect 34149 32895 34207 32901
rect 34149 32861 34161 32895
rect 34195 32892 34207 32895
rect 34330 32892 34336 32904
rect 34195 32864 34336 32892
rect 34195 32861 34207 32864
rect 34149 32855 34207 32861
rect 34330 32852 34336 32864
rect 34388 32852 34394 32904
rect 35544 32892 35572 32988
rect 35710 32920 35716 32972
rect 35768 32960 35774 32972
rect 38657 32963 38715 32969
rect 35768 32932 37044 32960
rect 35768 32920 35774 32932
rect 37016 32901 37044 32932
rect 38657 32929 38669 32963
rect 38703 32960 38715 32963
rect 39022 32960 39028 32972
rect 38703 32932 39028 32960
rect 38703 32929 38715 32932
rect 38657 32923 38715 32929
rect 39022 32920 39028 32932
rect 39080 32920 39086 32972
rect 37001 32895 37059 32901
rect 35544 32864 35650 32892
rect 37001 32861 37013 32895
rect 37047 32861 37059 32895
rect 37001 32855 37059 32861
rect 37274 32852 37280 32904
rect 37332 32852 37338 32904
rect 37366 32852 37372 32904
rect 37424 32852 37430 32904
rect 39500 32901 39528 33068
rect 39850 33056 39856 33068
rect 39908 33056 39914 33108
rect 40218 33056 40224 33108
rect 40276 33096 40282 33108
rect 41601 33099 41659 33105
rect 41601 33096 41613 33099
rect 40276 33068 41613 33096
rect 40276 33056 40282 33068
rect 41601 33065 41613 33068
rect 41647 33065 41659 33099
rect 41601 33059 41659 33065
rect 39669 33031 39727 33037
rect 39669 32997 39681 33031
rect 39715 32997 39727 33031
rect 39669 32991 39727 32997
rect 39684 32960 39712 32991
rect 40129 32963 40187 32969
rect 40129 32960 40141 32963
rect 39684 32932 40141 32960
rect 40129 32929 40141 32932
rect 40175 32929 40187 32963
rect 40129 32923 40187 32929
rect 40678 32920 40684 32972
rect 40736 32960 40742 32972
rect 40736 32932 41828 32960
rect 40736 32920 40742 32932
rect 41800 32901 41828 32932
rect 37645 32895 37703 32901
rect 37645 32861 37657 32895
rect 37691 32892 37703 32895
rect 39485 32895 39543 32901
rect 37691 32864 38056 32892
rect 37691 32861 37703 32864
rect 37645 32855 37703 32861
rect 31757 32796 32536 32824
rect 32600 32796 33364 32824
rect 31757 32793 31769 32796
rect 31720 32787 31769 32793
rect 31720 32784 31726 32787
rect 28077 32759 28135 32765
rect 28077 32756 28089 32759
rect 27396 32728 28089 32756
rect 27396 32716 27402 32728
rect 28077 32725 28089 32728
rect 28123 32725 28135 32759
rect 28077 32719 28135 32725
rect 28626 32716 28632 32768
rect 28684 32716 28690 32768
rect 32125 32759 32183 32765
rect 32125 32725 32137 32759
rect 32171 32756 32183 32759
rect 32214 32756 32220 32768
rect 32171 32728 32220 32756
rect 32171 32725 32183 32728
rect 32125 32719 32183 32725
rect 32214 32716 32220 32728
rect 32272 32716 32278 32768
rect 32508 32756 32536 32796
rect 33870 32784 33876 32836
rect 33928 32824 33934 32836
rect 33965 32827 34023 32833
rect 33965 32824 33977 32827
rect 33928 32796 33977 32824
rect 33928 32784 33934 32796
rect 33965 32793 33977 32796
rect 34011 32793 34023 32827
rect 33965 32787 34023 32793
rect 34054 32784 34060 32836
rect 34112 32784 34118 32836
rect 34514 32784 34520 32836
rect 34572 32784 34578 32836
rect 36630 32784 36636 32836
rect 36688 32824 36694 32836
rect 36725 32827 36783 32833
rect 36725 32824 36737 32827
rect 36688 32796 36737 32824
rect 36688 32784 36694 32796
rect 36725 32793 36737 32796
rect 36771 32793 36783 32827
rect 36725 32787 36783 32793
rect 33318 32756 33324 32768
rect 32508 32728 33324 32756
rect 33318 32716 33324 32728
rect 33376 32756 33382 32768
rect 34532 32756 34560 32784
rect 38028 32768 38056 32864
rect 39485 32861 39497 32895
rect 39531 32861 39543 32895
rect 39485 32855 39543 32861
rect 39853 32895 39911 32901
rect 39853 32861 39865 32895
rect 39899 32861 39911 32895
rect 39853 32855 39911 32861
rect 41785 32895 41843 32901
rect 41785 32861 41797 32895
rect 41831 32861 41843 32895
rect 41785 32855 41843 32861
rect 33376 32728 34560 32756
rect 33376 32716 33382 32728
rect 38010 32716 38016 32768
rect 38068 32716 38074 32768
rect 39868 32756 39896 32855
rect 40402 32784 40408 32836
rect 40460 32784 40466 32836
rect 40586 32824 40592 32836
rect 40512 32796 40592 32824
rect 40420 32756 40448 32784
rect 39868 32728 40448 32756
rect 40512 32756 40540 32796
rect 40586 32784 40592 32796
rect 40644 32784 40650 32836
rect 41138 32756 41144 32768
rect 40512 32728 41144 32756
rect 41138 32716 41144 32728
rect 41196 32756 41202 32768
rect 41877 32759 41935 32765
rect 41877 32756 41889 32759
rect 41196 32728 41889 32756
rect 41196 32716 41202 32728
rect 41877 32725 41889 32728
rect 41923 32756 41935 32759
rect 43438 32756 43444 32768
rect 41923 32728 43444 32756
rect 41923 32725 41935 32728
rect 41877 32719 41935 32725
rect 43438 32716 43444 32728
rect 43496 32716 43502 32768
rect 1104 32666 45172 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 45172 32666
rect 1104 32592 45172 32614
rect 2869 32555 2927 32561
rect 2869 32521 2881 32555
rect 2915 32552 2927 32555
rect 3234 32552 3240 32564
rect 2915 32524 3240 32552
rect 2915 32521 2927 32524
rect 2869 32515 2927 32521
rect 3234 32512 3240 32524
rect 3292 32512 3298 32564
rect 3786 32512 3792 32564
rect 3844 32512 3850 32564
rect 6454 32552 6460 32564
rect 3896 32524 6460 32552
rect 1762 32493 1768 32496
rect 1756 32484 1768 32493
rect 1723 32456 1768 32484
rect 1756 32447 1768 32456
rect 1762 32444 1768 32447
rect 1820 32444 1826 32496
rect 3896 32493 3924 32524
rect 6454 32512 6460 32524
rect 6512 32512 6518 32564
rect 6730 32512 6736 32564
rect 6788 32512 6794 32564
rect 6822 32512 6828 32564
rect 6880 32512 6886 32564
rect 7098 32512 7104 32564
rect 7156 32512 7162 32564
rect 7190 32512 7196 32564
rect 7248 32512 7254 32564
rect 7282 32512 7288 32564
rect 7340 32512 7346 32564
rect 7837 32555 7895 32561
rect 7837 32521 7849 32555
rect 7883 32552 7895 32555
rect 8018 32552 8024 32564
rect 7883 32524 8024 32552
rect 7883 32521 7895 32524
rect 7837 32515 7895 32521
rect 8018 32512 8024 32524
rect 8076 32512 8082 32564
rect 8386 32512 8392 32564
rect 8444 32552 8450 32564
rect 10134 32552 10140 32564
rect 8444 32524 10140 32552
rect 8444 32512 8450 32524
rect 10134 32512 10140 32524
rect 10192 32512 10198 32564
rect 10226 32512 10232 32564
rect 10284 32552 10290 32564
rect 10284 32524 12434 32552
rect 10284 32512 10290 32524
rect 3881 32487 3939 32493
rect 3881 32453 3893 32487
rect 3927 32453 3939 32487
rect 3881 32447 3939 32453
rect 5166 32444 5172 32496
rect 5224 32484 5230 32496
rect 5629 32487 5687 32493
rect 5629 32484 5641 32487
rect 5224 32456 5641 32484
rect 5224 32444 5230 32456
rect 5629 32453 5641 32456
rect 5675 32484 5687 32487
rect 7116 32484 7144 32512
rect 5675 32456 7144 32484
rect 7300 32484 7328 32512
rect 7300 32456 8064 32484
rect 5675 32453 5687 32456
rect 5629 32447 5687 32453
rect 3050 32376 3056 32428
rect 3108 32416 3114 32428
rect 3145 32419 3203 32425
rect 3145 32416 3157 32419
rect 3108 32388 3157 32416
rect 3108 32376 3114 32388
rect 3145 32385 3157 32388
rect 3191 32385 3203 32419
rect 3145 32379 3203 32385
rect 6086 32376 6092 32428
rect 6144 32376 6150 32428
rect 6181 32419 6239 32425
rect 6181 32385 6193 32419
rect 6227 32385 6239 32419
rect 6181 32379 6239 32385
rect 1486 32308 1492 32360
rect 1544 32308 1550 32360
rect 6104 32280 6132 32376
rect 6196 32348 6224 32379
rect 6270 32376 6276 32428
rect 6328 32416 6334 32428
rect 7377 32419 7435 32425
rect 6328 32388 6960 32416
rect 6328 32376 6334 32388
rect 6932 32357 6960 32388
rect 7377 32385 7389 32419
rect 7423 32416 7435 32419
rect 7423 32388 7512 32416
rect 7423 32385 7435 32388
rect 7377 32379 7435 32385
rect 6917 32351 6975 32357
rect 6196 32320 6592 32348
rect 6365 32283 6423 32289
rect 6365 32280 6377 32283
rect 6104 32252 6377 32280
rect 6365 32249 6377 32252
rect 6411 32249 6423 32283
rect 6564 32280 6592 32320
rect 6917 32317 6929 32351
rect 6963 32317 6975 32351
rect 6917 32311 6975 32317
rect 7374 32280 7380 32292
rect 6564 32252 7380 32280
rect 6365 32243 6423 32249
rect 7374 32240 7380 32252
rect 7432 32240 7438 32292
rect 7484 32289 7512 32388
rect 7650 32308 7656 32360
rect 7708 32348 7714 32360
rect 8036 32357 8064 32456
rect 9582 32444 9588 32496
rect 9640 32484 9646 32496
rect 12406 32484 12434 32524
rect 12710 32512 12716 32564
rect 12768 32512 12774 32564
rect 13170 32552 13176 32564
rect 12820 32524 13176 32552
rect 9640 32456 10447 32484
rect 9640 32444 9646 32456
rect 10042 32376 10048 32428
rect 10100 32376 10106 32428
rect 10226 32376 10232 32428
rect 10284 32376 10290 32428
rect 10321 32419 10379 32425
rect 10321 32385 10333 32419
rect 10367 32385 10379 32419
rect 10419 32416 10447 32456
rect 12360 32456 12572 32484
rect 10689 32419 10747 32425
rect 10689 32416 10701 32419
rect 10419 32388 10701 32416
rect 10321 32379 10379 32385
rect 10689 32385 10701 32388
rect 10735 32416 10747 32419
rect 10781 32419 10839 32425
rect 10781 32416 10793 32419
rect 10735 32388 10793 32416
rect 10735 32385 10747 32388
rect 10689 32379 10747 32385
rect 10781 32385 10793 32388
rect 10827 32385 10839 32419
rect 10781 32379 10839 32385
rect 10965 32419 11023 32425
rect 10965 32385 10977 32419
rect 11011 32416 11023 32419
rect 12158 32416 12164 32428
rect 11011 32388 12164 32416
rect 11011 32385 11023 32388
rect 10965 32379 11023 32385
rect 7929 32351 7987 32357
rect 7929 32348 7941 32351
rect 7708 32320 7941 32348
rect 7708 32308 7714 32320
rect 7929 32317 7941 32320
rect 7975 32317 7987 32351
rect 7929 32311 7987 32317
rect 8021 32351 8079 32357
rect 8021 32317 8033 32351
rect 8067 32317 8079 32351
rect 10060 32348 10088 32376
rect 10336 32348 10364 32379
rect 10060 32320 10364 32348
rect 10597 32351 10655 32357
rect 8021 32311 8079 32317
rect 10597 32317 10609 32351
rect 10643 32348 10655 32351
rect 10980 32348 11008 32379
rect 12158 32376 12164 32388
rect 12216 32376 12222 32428
rect 10643 32320 11008 32348
rect 10643 32317 10655 32320
rect 10597 32311 10655 32317
rect 12250 32308 12256 32360
rect 12308 32308 12314 32360
rect 7469 32283 7527 32289
rect 7469 32249 7481 32283
rect 7515 32249 7527 32283
rect 7469 32243 7527 32249
rect 10134 32240 10140 32292
rect 10192 32280 10198 32292
rect 10781 32283 10839 32289
rect 10781 32280 10793 32283
rect 10192 32252 10793 32280
rect 10192 32240 10198 32252
rect 10781 32249 10793 32252
rect 10827 32249 10839 32283
rect 12360 32280 12388 32456
rect 12434 32376 12440 32428
rect 12492 32376 12498 32428
rect 12544 32425 12572 32456
rect 12728 32425 12756 32512
rect 12529 32419 12587 32425
rect 12529 32385 12541 32419
rect 12575 32385 12587 32419
rect 12529 32379 12587 32385
rect 12713 32419 12771 32425
rect 12713 32385 12725 32419
rect 12759 32385 12771 32419
rect 12713 32379 12771 32385
rect 12452 32348 12480 32376
rect 12820 32348 12848 32524
rect 13170 32512 13176 32524
rect 13228 32512 13234 32564
rect 15102 32512 15108 32564
rect 15160 32512 15166 32564
rect 15194 32512 15200 32564
rect 15252 32552 15258 32564
rect 15657 32555 15715 32561
rect 15657 32552 15669 32555
rect 15252 32524 15669 32552
rect 15252 32512 15258 32524
rect 15657 32521 15669 32524
rect 15703 32521 15715 32555
rect 15657 32515 15715 32521
rect 15930 32512 15936 32564
rect 15988 32552 15994 32564
rect 15988 32524 16160 32552
rect 15988 32512 15994 32524
rect 13541 32487 13599 32493
rect 13541 32484 13553 32487
rect 12452 32320 12848 32348
rect 12912 32456 13553 32484
rect 12912 32280 12940 32456
rect 13541 32453 13553 32456
rect 13587 32484 13599 32487
rect 15120 32484 15148 32512
rect 13587 32456 15148 32484
rect 13587 32453 13599 32456
rect 13541 32447 13599 32453
rect 15286 32444 15292 32496
rect 15344 32484 15350 32496
rect 15344 32456 15976 32484
rect 15344 32444 15350 32456
rect 13170 32376 13176 32428
rect 13228 32416 13234 32428
rect 13403 32419 13461 32425
rect 13403 32416 13415 32419
rect 13228 32388 13415 32416
rect 13228 32376 13234 32388
rect 13403 32385 13415 32388
rect 13449 32385 13461 32419
rect 13403 32379 13461 32385
rect 13630 32376 13636 32428
rect 13688 32376 13694 32428
rect 13761 32419 13819 32425
rect 13761 32416 13773 32419
rect 13740 32385 13773 32416
rect 13807 32385 13819 32419
rect 13740 32379 13819 32385
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32416 13967 32419
rect 15654 32416 15660 32428
rect 13955 32388 15660 32416
rect 13955 32385 13967 32388
rect 13909 32379 13967 32385
rect 12986 32308 12992 32360
rect 13044 32348 13050 32360
rect 13740 32348 13768 32379
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15746 32376 15752 32428
rect 15804 32416 15810 32428
rect 15948 32425 15976 32456
rect 16132 32425 16160 32524
rect 16298 32512 16304 32564
rect 16356 32552 16362 32564
rect 16393 32555 16451 32561
rect 16393 32552 16405 32555
rect 16356 32524 16405 32552
rect 16356 32512 16362 32524
rect 16393 32521 16405 32524
rect 16439 32521 16451 32555
rect 16393 32515 16451 32521
rect 16408 32484 16436 32515
rect 17034 32512 17040 32564
rect 17092 32552 17098 32564
rect 17218 32552 17224 32564
rect 17092 32524 17224 32552
rect 17092 32512 17098 32524
rect 17218 32512 17224 32524
rect 17276 32512 17282 32564
rect 17402 32512 17408 32564
rect 17460 32512 17466 32564
rect 17862 32552 17868 32564
rect 17512 32524 17868 32552
rect 16761 32487 16819 32493
rect 16761 32484 16773 32487
rect 16408 32456 16773 32484
rect 16761 32453 16773 32456
rect 16807 32453 16819 32487
rect 17420 32484 17448 32512
rect 17512 32493 17540 32524
rect 17862 32512 17868 32524
rect 17920 32512 17926 32564
rect 18230 32512 18236 32564
rect 18288 32512 18294 32564
rect 18966 32512 18972 32564
rect 19024 32512 19030 32564
rect 19058 32512 19064 32564
rect 19116 32552 19122 32564
rect 21361 32555 21419 32561
rect 21361 32552 21373 32555
rect 19116 32524 21373 32552
rect 19116 32512 19122 32524
rect 21361 32521 21373 32524
rect 21407 32521 21419 32555
rect 21361 32515 21419 32521
rect 22833 32555 22891 32561
rect 22833 32521 22845 32555
rect 22879 32521 22891 32555
rect 22833 32515 22891 32521
rect 16761 32447 16819 32453
rect 16868 32456 17448 32484
rect 17497 32487 17555 32493
rect 15841 32419 15899 32425
rect 15841 32416 15853 32419
rect 15804 32388 15853 32416
rect 15804 32376 15810 32388
rect 15841 32385 15853 32388
rect 15887 32385 15899 32419
rect 15841 32379 15899 32385
rect 15933 32419 15991 32425
rect 15933 32385 15945 32419
rect 15979 32385 15991 32419
rect 15933 32379 15991 32385
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 13044 32320 13768 32348
rect 13044 32308 13050 32320
rect 12360 32252 12940 32280
rect 10781 32243 10839 32249
rect 5997 32215 6055 32221
rect 5997 32181 6009 32215
rect 6043 32212 6055 32215
rect 6822 32212 6828 32224
rect 6043 32184 6828 32212
rect 6043 32181 6055 32184
rect 5997 32175 6055 32181
rect 6822 32172 6828 32184
rect 6880 32172 6886 32224
rect 9490 32172 9496 32224
rect 9548 32212 9554 32224
rect 10045 32215 10103 32221
rect 10045 32212 10057 32215
rect 9548 32184 10057 32212
rect 9548 32172 9554 32184
rect 10045 32181 10057 32184
rect 10091 32212 10103 32215
rect 10318 32212 10324 32224
rect 10091 32184 10324 32212
rect 10091 32181 10103 32184
rect 10045 32175 10103 32181
rect 10318 32172 10324 32184
rect 10376 32172 10382 32224
rect 12710 32172 12716 32224
rect 12768 32172 12774 32224
rect 13265 32215 13323 32221
rect 13265 32181 13277 32215
rect 13311 32212 13323 32215
rect 13906 32212 13912 32224
rect 13311 32184 13912 32212
rect 13311 32181 13323 32184
rect 13265 32175 13323 32181
rect 13906 32172 13912 32184
rect 13964 32172 13970 32224
rect 15948 32212 15976 32379
rect 16206 32376 16212 32428
rect 16264 32416 16270 32428
rect 16301 32419 16359 32425
rect 16301 32416 16313 32419
rect 16264 32388 16313 32416
rect 16264 32376 16270 32388
rect 16301 32385 16313 32388
rect 16347 32385 16359 32419
rect 16301 32379 16359 32385
rect 16485 32419 16543 32425
rect 16485 32385 16497 32419
rect 16531 32416 16543 32419
rect 16868 32416 16896 32456
rect 17497 32453 17509 32487
rect 17543 32453 17555 32487
rect 18248 32484 18276 32512
rect 17497 32447 17555 32453
rect 17788 32456 18276 32484
rect 16531 32388 16896 32416
rect 16945 32419 17003 32425
rect 16531 32385 16543 32388
rect 16485 32379 16543 32385
rect 16945 32385 16957 32419
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 16025 32351 16083 32357
rect 16025 32317 16037 32351
rect 16071 32317 16083 32351
rect 16025 32311 16083 32317
rect 16040 32280 16068 32311
rect 16666 32308 16672 32360
rect 16724 32308 16730 32360
rect 16960 32348 16988 32379
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 17126 32376 17132 32428
rect 17184 32416 17190 32428
rect 17788 32425 17816 32456
rect 17313 32419 17371 32425
rect 17313 32416 17325 32419
rect 17184 32388 17325 32416
rect 17184 32376 17190 32388
rect 17313 32385 17325 32388
rect 17359 32385 17371 32419
rect 17313 32379 17371 32385
rect 17773 32419 17831 32425
rect 17773 32385 17785 32419
rect 17819 32385 17831 32419
rect 17773 32379 17831 32385
rect 18141 32419 18199 32425
rect 18141 32385 18153 32419
rect 18187 32416 18199 32419
rect 18322 32416 18328 32428
rect 18187 32388 18328 32416
rect 18187 32385 18199 32388
rect 18141 32379 18199 32385
rect 18322 32376 18328 32388
rect 18380 32376 18386 32428
rect 18414 32376 18420 32428
rect 18472 32416 18478 32428
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 18472 32388 18705 32416
rect 18472 32376 18478 32388
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18693 32379 18751 32385
rect 18782 32376 18788 32428
rect 18840 32376 18846 32428
rect 17865 32351 17923 32357
rect 17865 32348 17877 32351
rect 16960 32320 17877 32348
rect 17865 32317 17877 32320
rect 17911 32348 17923 32351
rect 18233 32351 18291 32357
rect 18233 32348 18245 32351
rect 17911 32320 18245 32348
rect 17911 32317 17923 32320
rect 17865 32311 17923 32317
rect 18233 32317 18245 32320
rect 18279 32317 18291 32351
rect 18233 32311 18291 32317
rect 16684 32280 16712 32308
rect 16040 32252 16712 32280
rect 16761 32283 16819 32289
rect 16761 32249 16773 32283
rect 16807 32280 16819 32283
rect 17586 32280 17592 32292
rect 16807 32252 17592 32280
rect 16807 32249 16819 32252
rect 16761 32243 16819 32249
rect 17586 32240 17592 32252
rect 17644 32240 17650 32292
rect 18049 32283 18107 32289
rect 18049 32249 18061 32283
rect 18095 32280 18107 32283
rect 18800 32280 18828 32376
rect 18095 32252 18828 32280
rect 18095 32249 18107 32252
rect 18049 32243 18107 32249
rect 17129 32215 17187 32221
rect 17129 32212 17141 32215
rect 15948 32184 17141 32212
rect 17129 32181 17141 32184
rect 17175 32181 17187 32215
rect 17129 32175 17187 32181
rect 17218 32172 17224 32224
rect 17276 32212 17282 32224
rect 17681 32215 17739 32221
rect 17681 32212 17693 32215
rect 17276 32184 17693 32212
rect 17276 32172 17282 32184
rect 17681 32181 17693 32184
rect 17727 32181 17739 32215
rect 17681 32175 17739 32181
rect 18601 32215 18659 32221
rect 18601 32181 18613 32215
rect 18647 32212 18659 32215
rect 18984 32212 19012 32512
rect 22848 32484 22876 32515
rect 23106 32512 23112 32564
rect 23164 32552 23170 32564
rect 23164 32524 24900 32552
rect 23164 32512 23170 32524
rect 23201 32487 23259 32493
rect 23201 32484 23213 32487
rect 22848 32456 23213 32484
rect 23201 32453 23213 32456
rect 23247 32453 23259 32487
rect 24762 32484 24768 32496
rect 24426 32456 24768 32484
rect 23201 32447 23259 32453
rect 24762 32444 24768 32456
rect 24820 32444 24826 32496
rect 24872 32484 24900 32524
rect 26050 32512 26056 32564
rect 26108 32552 26114 32564
rect 26973 32555 27031 32561
rect 26973 32552 26985 32555
rect 26108 32524 26985 32552
rect 26108 32512 26114 32524
rect 26973 32521 26985 32524
rect 27019 32521 27031 32555
rect 26973 32515 27031 32521
rect 27338 32512 27344 32564
rect 27396 32512 27402 32564
rect 28626 32512 28632 32564
rect 28684 32512 28690 32564
rect 29638 32512 29644 32564
rect 29696 32552 29702 32564
rect 29733 32555 29791 32561
rect 29733 32552 29745 32555
rect 29696 32524 29745 32552
rect 29696 32512 29702 32524
rect 29733 32521 29745 32524
rect 29779 32521 29791 32555
rect 29733 32515 29791 32521
rect 30926 32512 30932 32564
rect 30984 32512 30990 32564
rect 31386 32512 31392 32564
rect 31444 32552 31450 32564
rect 32125 32555 32183 32561
rect 32125 32552 32137 32555
rect 31444 32524 32137 32552
rect 31444 32512 31450 32524
rect 32125 32521 32137 32524
rect 32171 32521 32183 32555
rect 32125 32515 32183 32521
rect 33229 32555 33287 32561
rect 33229 32521 33241 32555
rect 33275 32552 33287 32555
rect 33778 32552 33784 32564
rect 33275 32524 33784 32552
rect 33275 32521 33287 32524
rect 33229 32515 33287 32521
rect 33778 32512 33784 32524
rect 33836 32512 33842 32564
rect 40313 32555 40371 32561
rect 40313 32521 40325 32555
rect 40359 32521 40371 32555
rect 40313 32515 40371 32521
rect 28644 32484 28672 32512
rect 24872 32456 28672 32484
rect 30944 32484 30972 32512
rect 31573 32487 31631 32493
rect 31573 32484 31585 32487
rect 30944 32456 31585 32484
rect 31573 32453 31585 32456
rect 31619 32453 31631 32487
rect 31573 32447 31631 32453
rect 31754 32444 31760 32496
rect 31812 32444 31818 32496
rect 31941 32487 31999 32493
rect 31941 32453 31953 32487
rect 31987 32484 31999 32487
rect 32214 32484 32220 32496
rect 31987 32456 32220 32484
rect 31987 32453 31999 32456
rect 31941 32447 31999 32453
rect 32214 32444 32220 32456
rect 32272 32484 32278 32496
rect 33594 32484 33600 32496
rect 32272 32456 33600 32484
rect 32272 32444 32278 32456
rect 33594 32444 33600 32456
rect 33652 32444 33658 32496
rect 40328 32484 40356 32515
rect 43898 32512 43904 32564
rect 43956 32512 43962 32564
rect 40681 32487 40739 32493
rect 40681 32484 40693 32487
rect 40328 32456 40693 32484
rect 40681 32453 40693 32456
rect 40727 32453 40739 32487
rect 40681 32447 40739 32453
rect 41138 32444 41144 32496
rect 41196 32444 41202 32496
rect 21266 32376 21272 32428
rect 21324 32376 21330 32428
rect 22649 32419 22707 32425
rect 22649 32385 22661 32419
rect 22695 32416 22707 32419
rect 22830 32416 22836 32428
rect 22695 32388 22836 32416
rect 22695 32385 22707 32388
rect 22649 32379 22707 32385
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 28902 32376 28908 32428
rect 28960 32416 28966 32428
rect 29273 32419 29331 32425
rect 29273 32416 29285 32419
rect 28960 32388 29285 32416
rect 28960 32376 28966 32388
rect 29273 32385 29285 32388
rect 29319 32385 29331 32419
rect 29273 32379 29331 32385
rect 29549 32419 29607 32425
rect 29549 32385 29561 32419
rect 29595 32416 29607 32419
rect 29914 32416 29920 32428
rect 29595 32388 29920 32416
rect 29595 32385 29607 32388
rect 29549 32379 29607 32385
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 30190 32376 30196 32428
rect 30248 32376 30254 32428
rect 30834 32376 30840 32428
rect 30892 32376 30898 32428
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 32398 32416 32404 32428
rect 32355 32388 32404 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 32493 32419 32551 32425
rect 32493 32385 32505 32419
rect 32539 32416 32551 32419
rect 32582 32416 32588 32428
rect 32539 32388 32588 32416
rect 32539 32385 32551 32388
rect 32493 32379 32551 32385
rect 32582 32376 32588 32388
rect 32640 32376 32646 32428
rect 32861 32419 32919 32425
rect 32861 32385 32873 32419
rect 32907 32416 32919 32419
rect 33042 32416 33048 32428
rect 32907 32388 33048 32416
rect 32907 32385 32919 32388
rect 32861 32379 32919 32385
rect 33042 32376 33048 32388
rect 33100 32416 33106 32428
rect 33410 32416 33416 32428
rect 33100 32388 33416 32416
rect 33100 32376 33106 32388
rect 33410 32376 33416 32388
rect 33468 32376 33474 32428
rect 40126 32376 40132 32428
rect 40184 32376 40190 32428
rect 43916 32416 43944 32512
rect 43993 32419 44051 32425
rect 43993 32416 44005 32419
rect 43916 32388 44005 32416
rect 43993 32385 44005 32388
rect 44039 32385 44051 32419
rect 43993 32379 44051 32385
rect 21082 32308 21088 32360
rect 21140 32308 21146 32360
rect 21818 32308 21824 32360
rect 21876 32348 21882 32360
rect 22925 32351 22983 32357
rect 22925 32348 22937 32351
rect 21876 32320 22937 32348
rect 21876 32308 21882 32320
rect 22925 32317 22937 32320
rect 22971 32317 22983 32351
rect 22925 32311 22983 32317
rect 25958 32308 25964 32360
rect 26016 32308 26022 32360
rect 27430 32308 27436 32360
rect 27488 32308 27494 32360
rect 27522 32308 27528 32360
rect 27580 32348 27586 32360
rect 27617 32351 27675 32357
rect 27617 32348 27629 32351
rect 27580 32320 27629 32348
rect 27580 32308 27586 32320
rect 27617 32317 27629 32320
rect 27663 32348 27675 32351
rect 27663 32320 28856 32348
rect 27663 32317 27675 32320
rect 27617 32311 27675 32317
rect 28828 32292 28856 32320
rect 29362 32308 29368 32360
rect 29420 32348 29426 32360
rect 30208 32348 30236 32376
rect 29420 32320 30236 32348
rect 32953 32351 33011 32357
rect 29420 32308 29426 32320
rect 32953 32317 32965 32351
rect 32999 32348 33011 32351
rect 33134 32348 33140 32360
rect 32999 32320 33140 32348
rect 32999 32317 33011 32320
rect 32953 32311 33011 32317
rect 33134 32308 33140 32320
rect 33192 32308 33198 32360
rect 40402 32308 40408 32360
rect 40460 32308 40466 32360
rect 28810 32240 28816 32292
rect 28868 32280 28874 32292
rect 28868 32252 36676 32280
rect 28868 32240 28874 32252
rect 36648 32224 36676 32252
rect 18647 32184 19012 32212
rect 18647 32181 18659 32184
rect 18601 32175 18659 32181
rect 20530 32172 20536 32224
rect 20588 32172 20594 32224
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 23566 32212 23572 32224
rect 22796 32184 23572 32212
rect 22796 32172 22802 32184
rect 23566 32172 23572 32184
rect 23624 32212 23630 32224
rect 24673 32215 24731 32221
rect 24673 32212 24685 32215
rect 23624 32184 24685 32212
rect 23624 32172 23630 32184
rect 24673 32181 24685 32184
rect 24719 32181 24731 32215
rect 24673 32175 24731 32181
rect 26510 32172 26516 32224
rect 26568 32172 26574 32224
rect 32674 32172 32680 32224
rect 32732 32212 32738 32224
rect 33778 32212 33784 32224
rect 32732 32184 33784 32212
rect 32732 32172 32738 32184
rect 33778 32172 33784 32184
rect 33836 32172 33842 32224
rect 36630 32172 36636 32224
rect 36688 32172 36694 32224
rect 36814 32172 36820 32224
rect 36872 32212 36878 32224
rect 40678 32212 40684 32224
rect 36872 32184 40684 32212
rect 36872 32172 36878 32184
rect 40678 32172 40684 32184
rect 40736 32172 40742 32224
rect 41230 32172 41236 32224
rect 41288 32212 41294 32224
rect 42153 32215 42211 32221
rect 42153 32212 42165 32215
rect 41288 32184 42165 32212
rect 41288 32172 41294 32184
rect 42153 32181 42165 32184
rect 42199 32181 42211 32215
rect 42153 32175 42211 32181
rect 43806 32172 43812 32224
rect 43864 32172 43870 32224
rect 1104 32122 45172 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 45172 32122
rect 1104 32048 45172 32070
rect 4614 31968 4620 32020
rect 4672 32008 4678 32020
rect 6178 32008 6184 32020
rect 4672 31980 6184 32008
rect 4672 31968 4678 31980
rect 6178 31968 6184 31980
rect 6236 31968 6242 32020
rect 6730 31968 6736 32020
rect 6788 31968 6794 32020
rect 7098 31968 7104 32020
rect 7156 32008 7162 32020
rect 7156 31980 10272 32008
rect 7156 31968 7162 31980
rect 2406 31832 2412 31884
rect 2464 31872 2470 31884
rect 2869 31875 2927 31881
rect 2869 31872 2881 31875
rect 2464 31844 2881 31872
rect 2464 31832 2470 31844
rect 2869 31841 2881 31844
rect 2915 31841 2927 31875
rect 2869 31835 2927 31841
rect 3053 31875 3111 31881
rect 3053 31841 3065 31875
rect 3099 31872 3111 31875
rect 4632 31872 4660 31968
rect 6748 31940 6776 31968
rect 7009 31943 7067 31949
rect 7009 31940 7021 31943
rect 6748 31912 7021 31940
rect 7009 31909 7021 31912
rect 7055 31909 7067 31943
rect 7009 31903 7067 31909
rect 9309 31943 9367 31949
rect 9309 31909 9321 31943
rect 9355 31940 9367 31943
rect 9861 31943 9919 31949
rect 9861 31940 9873 31943
rect 9355 31912 9873 31940
rect 9355 31909 9367 31912
rect 9309 31903 9367 31909
rect 9861 31909 9873 31912
rect 9907 31909 9919 31943
rect 9861 31903 9919 31909
rect 9953 31943 10011 31949
rect 9953 31909 9965 31943
rect 9999 31940 10011 31943
rect 10134 31940 10140 31952
rect 9999 31912 10140 31940
rect 9999 31909 10011 31912
rect 9953 31903 10011 31909
rect 10134 31900 10140 31912
rect 10192 31900 10198 31952
rect 10244 31940 10272 31980
rect 10318 31968 10324 32020
rect 10376 31968 10382 32020
rect 10781 32011 10839 32017
rect 10781 31977 10793 32011
rect 10827 32008 10839 32011
rect 11606 32008 11612 32020
rect 10827 31980 11612 32008
rect 10827 31977 10839 31980
rect 10781 31971 10839 31977
rect 11606 31968 11612 31980
rect 11664 31968 11670 32020
rect 12342 31968 12348 32020
rect 12400 32008 12406 32020
rect 14090 32008 14096 32020
rect 12400 31980 14096 32008
rect 12400 31968 12406 31980
rect 14090 31968 14096 31980
rect 14148 32008 14154 32020
rect 14185 32011 14243 32017
rect 14185 32008 14197 32011
rect 14148 31980 14197 32008
rect 14148 31968 14154 31980
rect 14185 31977 14197 31980
rect 14231 31977 14243 32011
rect 14185 31971 14243 31977
rect 14277 32011 14335 32017
rect 14277 31977 14289 32011
rect 14323 32008 14335 32011
rect 14826 32008 14832 32020
rect 14323 31980 14832 32008
rect 14323 31977 14335 31980
rect 14277 31971 14335 31977
rect 14826 31968 14832 31980
rect 14884 31968 14890 32020
rect 15654 31968 15660 32020
rect 15712 32008 15718 32020
rect 17313 32011 17371 32017
rect 17313 32008 17325 32011
rect 15712 31980 17325 32008
rect 15712 31968 15718 31980
rect 17313 31977 17325 31980
rect 17359 31977 17371 32011
rect 17770 32008 17776 32020
rect 17313 31971 17371 31977
rect 17420 31980 17776 32008
rect 12802 31940 12808 31952
rect 10244 31912 12808 31940
rect 12802 31900 12808 31912
rect 12860 31900 12866 31952
rect 13170 31940 13176 31952
rect 13096 31912 13176 31940
rect 3099 31844 4660 31872
rect 5445 31875 5503 31881
rect 3099 31841 3111 31844
rect 3053 31835 3111 31841
rect 5445 31841 5457 31875
rect 5491 31872 5503 31875
rect 5902 31872 5908 31884
rect 5491 31844 5908 31872
rect 5491 31841 5503 31844
rect 5445 31835 5503 31841
rect 5902 31832 5908 31844
rect 5960 31832 5966 31884
rect 6454 31832 6460 31884
rect 6512 31872 6518 31884
rect 6917 31875 6975 31881
rect 6512 31844 6868 31872
rect 6512 31832 6518 31844
rect 5166 31764 5172 31816
rect 5224 31764 5230 31816
rect 6840 31804 6868 31844
rect 6917 31841 6929 31875
rect 6963 31872 6975 31875
rect 7561 31875 7619 31881
rect 7561 31872 7573 31875
rect 6963 31844 7573 31872
rect 6963 31841 6975 31844
rect 6917 31835 6975 31841
rect 7561 31841 7573 31844
rect 7607 31841 7619 31875
rect 7561 31835 7619 31841
rect 9125 31875 9183 31881
rect 9125 31841 9137 31875
rect 9171 31872 9183 31875
rect 10413 31875 10471 31881
rect 10413 31872 10425 31875
rect 9171 31844 9812 31872
rect 9171 31841 9183 31844
rect 9125 31835 9183 31841
rect 7006 31804 7012 31816
rect 6578 31776 6776 31804
rect 6840 31776 7012 31804
rect 6748 31736 6776 31776
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 7576 31804 7604 31835
rect 7745 31807 7803 31813
rect 7745 31804 7757 31807
rect 7576 31776 7757 31804
rect 7745 31773 7757 31776
rect 7791 31773 7803 31807
rect 7745 31767 7803 31773
rect 7837 31807 7895 31813
rect 7837 31773 7849 31807
rect 7883 31804 7895 31807
rect 8294 31804 8300 31816
rect 7883 31776 8300 31804
rect 7883 31773 7895 31776
rect 7837 31767 7895 31773
rect 8294 31764 8300 31776
rect 8352 31764 8358 31816
rect 8386 31764 8392 31816
rect 8444 31764 8450 31816
rect 9217 31807 9275 31813
rect 9217 31773 9229 31807
rect 9263 31804 9275 31807
rect 9490 31804 9496 31816
rect 9263 31776 9496 31804
rect 9263 31773 9275 31776
rect 9217 31767 9275 31773
rect 9490 31764 9496 31776
rect 9548 31764 9554 31816
rect 9585 31807 9643 31813
rect 9585 31773 9597 31807
rect 9631 31804 9643 31807
rect 9674 31804 9680 31816
rect 9631 31776 9680 31804
rect 9631 31773 9643 31776
rect 9585 31767 9643 31773
rect 9674 31764 9680 31776
rect 9732 31764 9738 31816
rect 9784 31813 9812 31844
rect 9876 31844 10425 31872
rect 9769 31807 9827 31813
rect 9769 31773 9781 31807
rect 9815 31773 9827 31807
rect 9769 31767 9827 31773
rect 6822 31736 6828 31748
rect 6748 31708 6828 31736
rect 6822 31696 6828 31708
rect 6880 31736 6886 31748
rect 8404 31736 8432 31764
rect 6880 31708 8432 31736
rect 6880 31696 6886 31708
rect 9306 31696 9312 31748
rect 9364 31736 9370 31748
rect 9876 31736 9904 31844
rect 10413 31841 10425 31844
rect 10459 31841 10471 31875
rect 10413 31835 10471 31841
rect 12250 31832 12256 31884
rect 12308 31872 12314 31884
rect 12989 31875 13047 31881
rect 12989 31872 13001 31875
rect 12308 31844 13001 31872
rect 12308 31832 12314 31844
rect 12989 31841 13001 31844
rect 13035 31841 13047 31875
rect 12989 31835 13047 31841
rect 10042 31764 10048 31816
rect 10100 31764 10106 31816
rect 10226 31764 10232 31816
rect 10284 31804 10290 31816
rect 10597 31807 10655 31813
rect 10597 31804 10609 31807
rect 10284 31776 10609 31804
rect 10284 31764 10290 31776
rect 10597 31773 10609 31776
rect 10643 31773 10655 31807
rect 11974 31804 11980 31816
rect 10597 31767 10655 31773
rect 10704 31776 11980 31804
rect 9364 31708 9904 31736
rect 9364 31696 9370 31708
rect 10318 31696 10324 31748
rect 10376 31696 10382 31748
rect 2406 31628 2412 31680
rect 2464 31628 2470 31680
rect 2777 31671 2835 31677
rect 2777 31637 2789 31671
rect 2823 31668 2835 31671
rect 3234 31668 3240 31680
rect 2823 31640 3240 31668
rect 2823 31637 2835 31640
rect 2777 31631 2835 31637
rect 3234 31628 3240 31640
rect 3292 31628 3298 31680
rect 9398 31628 9404 31680
rect 9456 31668 9462 31680
rect 9493 31671 9551 31677
rect 9493 31668 9505 31671
rect 9456 31640 9505 31668
rect 9456 31628 9462 31640
rect 9493 31637 9505 31640
rect 9539 31637 9551 31671
rect 9493 31631 9551 31637
rect 9858 31628 9864 31680
rect 9916 31668 9922 31680
rect 10042 31668 10048 31680
rect 9916 31640 10048 31668
rect 9916 31628 9922 31640
rect 10042 31628 10048 31640
rect 10100 31628 10106 31680
rect 10229 31671 10287 31677
rect 10229 31637 10241 31671
rect 10275 31668 10287 31671
rect 10704 31668 10732 31776
rect 11974 31764 11980 31776
rect 12032 31764 12038 31816
rect 12158 31764 12164 31816
rect 12216 31804 12222 31816
rect 12897 31807 12955 31813
rect 12897 31804 12909 31807
rect 12216 31776 12909 31804
rect 12216 31764 12222 31776
rect 12897 31773 12909 31776
rect 12943 31804 12955 31807
rect 13096 31804 13124 31912
rect 13170 31900 13176 31912
rect 13228 31900 13234 31952
rect 17420 31940 17448 31980
rect 17770 31968 17776 31980
rect 17828 31968 17834 32020
rect 18046 31968 18052 32020
rect 18104 32008 18110 32020
rect 18104 31980 20024 32008
rect 18104 31968 18110 31980
rect 18138 31940 18144 31952
rect 14200 31912 17448 31940
rect 17604 31912 18144 31940
rect 13357 31875 13415 31881
rect 13357 31841 13369 31875
rect 13403 31872 13415 31875
rect 14200 31872 14228 31912
rect 13403 31844 14228 31872
rect 13403 31841 13415 31844
rect 13357 31835 13415 31841
rect 13556 31816 13584 31844
rect 14274 31832 14280 31884
rect 14332 31872 14338 31884
rect 14734 31872 14740 31884
rect 14332 31844 14740 31872
rect 14332 31832 14338 31844
rect 14734 31832 14740 31844
rect 14792 31832 14798 31884
rect 12943 31776 13124 31804
rect 13265 31807 13323 31813
rect 12943 31773 12955 31776
rect 12897 31767 12955 31773
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 13265 31767 13323 31773
rect 12250 31696 12256 31748
rect 12308 31736 12314 31748
rect 13280 31736 13308 31767
rect 13538 31764 13544 31816
rect 13596 31764 13602 31816
rect 13909 31807 13967 31813
rect 13909 31773 13921 31807
rect 13955 31773 13967 31807
rect 13909 31767 13967 31773
rect 14093 31807 14151 31813
rect 14093 31773 14105 31807
rect 14139 31804 14151 31807
rect 14366 31804 14372 31816
rect 14139 31776 14372 31804
rect 14139 31773 14151 31776
rect 14093 31767 14151 31773
rect 13630 31736 13636 31748
rect 12308 31708 13308 31736
rect 13556 31708 13636 31736
rect 12308 31696 12314 31708
rect 13556 31677 13584 31708
rect 13630 31696 13636 31708
rect 13688 31696 13694 31748
rect 13814 31696 13820 31748
rect 13872 31696 13878 31748
rect 13924 31736 13952 31767
rect 14366 31764 14372 31776
rect 14424 31764 14430 31816
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14642 31804 14648 31816
rect 14507 31776 14648 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 14642 31764 14648 31776
rect 14700 31804 14706 31816
rect 17604 31804 17632 31912
rect 18138 31900 18144 31912
rect 18196 31900 18202 31952
rect 19996 31884 20024 31980
rect 20530 31968 20536 32020
rect 20588 31968 20594 32020
rect 20625 32011 20683 32017
rect 20625 31977 20637 32011
rect 20671 32008 20683 32011
rect 21082 32008 21088 32020
rect 20671 31980 21088 32008
rect 20671 31977 20683 31980
rect 20625 31971 20683 31977
rect 21082 31968 21088 31980
rect 21140 31968 21146 32020
rect 22738 32008 22744 32020
rect 22572 31980 22744 32008
rect 17773 31875 17831 31881
rect 17773 31841 17785 31875
rect 17819 31872 17831 31875
rect 18230 31872 18236 31884
rect 17819 31844 18236 31872
rect 17819 31841 17831 31844
rect 17773 31835 17831 31841
rect 18230 31832 18236 31844
rect 18288 31872 18294 31884
rect 19150 31872 19156 31884
rect 18288 31844 19156 31872
rect 18288 31832 18294 31844
rect 19150 31832 19156 31844
rect 19208 31832 19214 31884
rect 19978 31832 19984 31884
rect 20036 31832 20042 31884
rect 14700 31776 17632 31804
rect 17681 31807 17739 31813
rect 14700 31764 14706 31776
rect 17681 31773 17693 31807
rect 17727 31804 17739 31807
rect 18414 31804 18420 31816
rect 17727 31776 18420 31804
rect 17727 31773 17739 31776
rect 17681 31767 17739 31773
rect 18414 31764 18420 31776
rect 18472 31764 18478 31816
rect 20349 31807 20407 31813
rect 19306 31776 20300 31804
rect 14182 31736 14188 31748
rect 13924 31708 14188 31736
rect 14182 31696 14188 31708
rect 14240 31736 14246 31748
rect 19306 31736 19334 31776
rect 14240 31708 19334 31736
rect 20272 31736 20300 31776
rect 20349 31773 20361 31807
rect 20395 31804 20407 31807
rect 20548 31804 20576 31968
rect 22186 31940 22192 31952
rect 21100 31912 22192 31940
rect 21100 31881 21128 31912
rect 22186 31900 22192 31912
rect 22244 31900 22250 31952
rect 21085 31875 21143 31881
rect 21085 31841 21097 31875
rect 21131 31841 21143 31875
rect 21085 31835 21143 31841
rect 21174 31832 21180 31884
rect 21232 31832 21238 31884
rect 22572 31872 22600 31980
rect 22738 31968 22744 31980
rect 22796 31968 22802 32020
rect 22830 31968 22836 32020
rect 22888 32008 22894 32020
rect 23477 32011 23535 32017
rect 23477 32008 23489 32011
rect 22888 31980 23489 32008
rect 22888 31968 22894 31980
rect 23477 31977 23489 31980
rect 23523 31977 23535 32011
rect 23477 31971 23535 31977
rect 23584 31980 25452 32008
rect 22649 31943 22707 31949
rect 22649 31909 22661 31943
rect 22695 31909 22707 31943
rect 22649 31903 22707 31909
rect 22848 31912 23336 31940
rect 21376 31844 22600 31872
rect 20395 31776 20576 31804
rect 20993 31807 21051 31813
rect 20395 31773 20407 31776
rect 20349 31767 20407 31773
rect 20993 31773 21005 31807
rect 21039 31804 21051 31807
rect 21266 31804 21272 31816
rect 21039 31776 21272 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21266 31764 21272 31776
rect 21324 31764 21330 31816
rect 21376 31736 21404 31844
rect 22189 31807 22247 31813
rect 22189 31773 22201 31807
rect 22235 31804 22247 31807
rect 22373 31807 22431 31813
rect 22235 31776 22324 31804
rect 22235 31773 22247 31776
rect 22189 31767 22247 31773
rect 20272 31708 21404 31736
rect 22296 31736 22324 31776
rect 22373 31773 22385 31807
rect 22419 31804 22431 31807
rect 22664 31804 22692 31903
rect 22848 31804 22876 31912
rect 23106 31832 23112 31884
rect 23164 31832 23170 31884
rect 23198 31832 23204 31884
rect 23256 31832 23262 31884
rect 22419 31776 22692 31804
rect 22756 31776 22876 31804
rect 23308 31804 23336 31912
rect 23382 31900 23388 31952
rect 23440 31940 23446 31952
rect 23584 31940 23612 31980
rect 23440 31912 23612 31940
rect 23440 31900 23446 31912
rect 24486 31900 24492 31952
rect 24544 31900 24550 31952
rect 24765 31943 24823 31949
rect 24765 31909 24777 31943
rect 24811 31909 24823 31943
rect 24765 31903 24823 31909
rect 25424 31940 25452 31980
rect 28626 31968 28632 32020
rect 28684 32008 28690 32020
rect 28721 32011 28779 32017
rect 28721 32008 28733 32011
rect 28684 31980 28733 32008
rect 28684 31968 28690 31980
rect 28721 31977 28733 31980
rect 28767 32008 28779 32011
rect 28902 32008 28908 32020
rect 28767 31980 28908 32008
rect 28767 31977 28779 31980
rect 28721 31971 28779 31977
rect 28902 31968 28908 31980
rect 28960 31968 28966 32020
rect 30101 32011 30159 32017
rect 30101 31977 30113 32011
rect 30147 32008 30159 32011
rect 30834 32008 30840 32020
rect 30147 31980 30840 32008
rect 30147 31977 30159 31980
rect 30101 31971 30159 31977
rect 30834 31968 30840 31980
rect 30892 31968 30898 32020
rect 32398 31968 32404 32020
rect 32456 32008 32462 32020
rect 33226 32008 33232 32020
rect 32456 31980 33232 32008
rect 32456 31968 32462 31980
rect 33226 31968 33232 31980
rect 33284 31968 33290 32020
rect 40126 31968 40132 32020
rect 40184 32008 40190 32020
rect 40865 32011 40923 32017
rect 40865 32008 40877 32011
rect 40184 31980 40877 32008
rect 40184 31968 40190 31980
rect 40865 31977 40877 31980
rect 40911 31977 40923 32011
rect 40865 31971 40923 31977
rect 26418 31940 26424 31952
rect 25424 31912 26424 31940
rect 24121 31875 24179 31881
rect 24121 31841 24133 31875
rect 24167 31872 24179 31875
rect 24210 31872 24216 31884
rect 24167 31844 24216 31872
rect 24167 31841 24179 31844
rect 24121 31835 24179 31841
rect 24210 31832 24216 31844
rect 24268 31872 24274 31884
rect 24504 31872 24532 31900
rect 24268 31844 24532 31872
rect 24268 31832 24274 31844
rect 23658 31804 23664 31816
rect 23308 31776 23664 31804
rect 22419 31773 22431 31776
rect 22373 31767 22431 31773
rect 22756 31736 22784 31776
rect 23658 31764 23664 31776
rect 23716 31764 23722 31816
rect 23937 31807 23995 31813
rect 23937 31773 23949 31807
rect 23983 31804 23995 31807
rect 24489 31807 24547 31813
rect 23983 31776 24440 31804
rect 23983 31773 23995 31776
rect 23937 31767 23995 31773
rect 22296 31708 22784 31736
rect 14240 31696 14246 31708
rect 23566 31696 23572 31748
rect 23624 31736 23630 31748
rect 23845 31739 23903 31745
rect 23845 31736 23857 31739
rect 23624 31708 23857 31736
rect 23624 31696 23630 31708
rect 23845 31705 23857 31708
rect 23891 31705 23903 31739
rect 24412 31736 24440 31776
rect 24489 31773 24501 31807
rect 24535 31804 24547 31807
rect 24780 31804 24808 31903
rect 25424 31881 25452 31912
rect 26418 31900 26424 31912
rect 26476 31900 26482 31952
rect 26881 31943 26939 31949
rect 26881 31909 26893 31943
rect 26927 31940 26939 31943
rect 26927 31912 27108 31940
rect 26927 31909 26939 31912
rect 26881 31903 26939 31909
rect 25409 31875 25467 31881
rect 25409 31841 25421 31875
rect 25455 31841 25467 31875
rect 25409 31835 25467 31841
rect 26326 31832 26332 31884
rect 26384 31872 26390 31884
rect 26973 31875 27031 31881
rect 26973 31872 26985 31875
rect 26384 31844 26985 31872
rect 26384 31832 26390 31844
rect 26973 31841 26985 31844
rect 27019 31841 27031 31875
rect 27080 31872 27108 31912
rect 28534 31900 28540 31952
rect 28592 31940 28598 31952
rect 28810 31940 28816 31952
rect 28592 31912 28816 31940
rect 28592 31900 28598 31912
rect 28810 31900 28816 31912
rect 28868 31900 28874 31952
rect 27249 31875 27307 31881
rect 27249 31872 27261 31875
rect 27080 31844 27261 31872
rect 26973 31835 27031 31841
rect 27249 31841 27261 31844
rect 27295 31841 27307 31875
rect 27249 31835 27307 31841
rect 27706 31832 27712 31884
rect 27764 31872 27770 31884
rect 28920 31872 28948 31968
rect 32490 31900 32496 31952
rect 32548 31900 32554 31952
rect 35805 31943 35863 31949
rect 35805 31909 35817 31943
rect 35851 31940 35863 31943
rect 35894 31940 35900 31952
rect 35851 31912 35900 31940
rect 35851 31909 35863 31912
rect 35805 31903 35863 31909
rect 35894 31900 35900 31912
rect 35952 31900 35958 31952
rect 36081 31943 36139 31949
rect 36081 31909 36093 31943
rect 36127 31909 36139 31943
rect 36081 31903 36139 31909
rect 38473 31943 38531 31949
rect 38473 31909 38485 31943
rect 38519 31909 38531 31943
rect 38473 31903 38531 31909
rect 42705 31943 42763 31949
rect 42705 31909 42717 31943
rect 42751 31909 42763 31943
rect 42705 31903 42763 31909
rect 27764 31844 28304 31872
rect 28920 31844 29776 31872
rect 27764 31832 27770 31844
rect 24535 31776 24808 31804
rect 25225 31807 25283 31813
rect 24535 31773 24547 31776
rect 24489 31767 24547 31773
rect 25225 31773 25237 31807
rect 25271 31804 25283 31807
rect 25498 31804 25504 31816
rect 25271 31776 25504 31804
rect 25271 31773 25283 31776
rect 25225 31767 25283 31773
rect 25498 31764 25504 31776
rect 25556 31764 25562 31816
rect 26234 31764 26240 31816
rect 26292 31764 26298 31816
rect 26510 31764 26516 31816
rect 26568 31764 26574 31816
rect 26694 31764 26700 31816
rect 26752 31764 26758 31816
rect 28276 31804 28304 31844
rect 28813 31807 28871 31813
rect 28813 31804 28825 31807
rect 28276 31776 28825 31804
rect 28813 31773 28825 31776
rect 28859 31773 28871 31807
rect 28813 31767 28871 31773
rect 29181 31807 29239 31813
rect 29181 31773 29193 31807
rect 29227 31804 29239 31807
rect 29270 31804 29276 31816
rect 29227 31776 29276 31804
rect 29227 31773 29239 31776
rect 29181 31767 29239 31773
rect 29270 31764 29276 31776
rect 29328 31764 29334 31816
rect 29748 31813 29776 31844
rect 29822 31832 29828 31884
rect 29880 31832 29886 31884
rect 32508 31872 32536 31900
rect 32324 31844 32536 31872
rect 32324 31816 32352 31844
rect 29733 31807 29791 31813
rect 29733 31773 29745 31807
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 32306 31764 32312 31816
rect 32364 31764 32370 31816
rect 32490 31764 32496 31816
rect 32548 31764 32554 31816
rect 34790 31764 34796 31816
rect 34848 31804 34854 31816
rect 35253 31807 35311 31813
rect 35253 31804 35265 31807
rect 34848 31776 35265 31804
rect 34848 31764 34854 31776
rect 35253 31773 35265 31776
rect 35299 31773 35311 31807
rect 35253 31767 35311 31773
rect 35989 31807 36047 31813
rect 35989 31773 36001 31807
rect 36035 31804 36047 31807
rect 36096 31804 36124 31903
rect 36538 31832 36544 31884
rect 36596 31832 36602 31884
rect 36630 31832 36636 31884
rect 36688 31832 36694 31884
rect 36035 31776 36124 31804
rect 38381 31807 38439 31813
rect 36035 31773 36047 31776
rect 35989 31767 36047 31773
rect 38381 31773 38393 31807
rect 38427 31804 38439 31807
rect 38488 31804 38516 31903
rect 38654 31832 38660 31884
rect 38712 31832 38718 31884
rect 38746 31832 38752 31884
rect 38804 31872 38810 31884
rect 38933 31875 38991 31881
rect 38933 31872 38945 31875
rect 38804 31844 38945 31872
rect 38804 31832 38810 31844
rect 38933 31841 38945 31844
rect 38979 31841 38991 31875
rect 38933 31835 38991 31841
rect 39025 31875 39083 31881
rect 39025 31841 39037 31875
rect 39071 31872 39083 31875
rect 40494 31872 40500 31884
rect 39071 31844 40500 31872
rect 39071 31841 39083 31844
rect 39025 31835 39083 31841
rect 38427 31776 38516 31804
rect 38672 31804 38700 31832
rect 39040 31804 39068 31835
rect 40494 31832 40500 31844
rect 40552 31872 40558 31884
rect 41417 31875 41475 31881
rect 41417 31872 41429 31875
rect 40552 31844 41429 31872
rect 40552 31832 40558 31844
rect 41417 31841 41429 31844
rect 41463 31841 41475 31875
rect 41417 31835 41475 31841
rect 41506 31832 41512 31884
rect 41564 31832 41570 31884
rect 42720 31872 42748 31903
rect 43073 31875 43131 31881
rect 43073 31872 43085 31875
rect 42720 31844 43085 31872
rect 43073 31841 43085 31844
rect 43119 31841 43131 31875
rect 43073 31835 43131 31841
rect 38672 31776 39068 31804
rect 38427 31773 38439 31776
rect 38381 31767 38439 31773
rect 41230 31764 41236 31816
rect 41288 31764 41294 31816
rect 41325 31807 41383 31813
rect 41325 31773 41337 31807
rect 41371 31804 41383 31807
rect 41524 31804 41552 31832
rect 41371 31776 41552 31804
rect 41371 31773 41383 31776
rect 41325 31767 41383 31773
rect 42518 31764 42524 31816
rect 42576 31764 42582 31816
rect 42794 31764 42800 31816
rect 42852 31764 42858 31816
rect 25133 31739 25191 31745
rect 25133 31736 25145 31739
rect 24412 31708 25145 31736
rect 23845 31699 23903 31705
rect 25133 31705 25145 31708
rect 25179 31736 25191 31739
rect 25593 31739 25651 31745
rect 25593 31736 25605 31739
rect 25179 31708 25605 31736
rect 25179 31705 25191 31708
rect 25133 31699 25191 31705
rect 25593 31705 25605 31708
rect 25639 31705 25651 31739
rect 25593 31699 25651 31705
rect 27706 31696 27712 31748
rect 27764 31696 27770 31748
rect 43530 31696 43536 31748
rect 43588 31696 43594 31748
rect 10275 31640 10732 31668
rect 13541 31671 13599 31677
rect 10275 31637 10287 31640
rect 10229 31631 10287 31637
rect 13541 31637 13553 31671
rect 13587 31637 13599 31671
rect 13541 31631 13599 31637
rect 20070 31628 20076 31680
rect 20128 31668 20134 31680
rect 20165 31671 20223 31677
rect 20165 31668 20177 31671
rect 20128 31640 20177 31668
rect 20128 31628 20134 31640
rect 20165 31637 20177 31640
rect 20211 31637 20223 31671
rect 20165 31631 20223 31637
rect 22005 31671 22063 31677
rect 22005 31637 22017 31671
rect 22051 31668 22063 31671
rect 22094 31668 22100 31680
rect 22051 31640 22100 31668
rect 22051 31637 22063 31640
rect 22005 31631 22063 31637
rect 22094 31628 22100 31640
rect 22152 31628 22158 31680
rect 22554 31628 22560 31680
rect 22612 31628 22618 31680
rect 23017 31671 23075 31677
rect 23017 31637 23029 31671
rect 23063 31668 23075 31671
rect 24118 31668 24124 31680
rect 23063 31640 24124 31668
rect 23063 31637 23075 31640
rect 23017 31631 23075 31637
rect 24118 31628 24124 31640
rect 24176 31628 24182 31680
rect 24673 31671 24731 31677
rect 24673 31637 24685 31671
rect 24719 31668 24731 31671
rect 24762 31668 24768 31680
rect 24719 31640 24768 31668
rect 24719 31637 24731 31640
rect 24673 31631 24731 31637
rect 24762 31628 24768 31640
rect 24820 31628 24826 31680
rect 26326 31628 26332 31680
rect 26384 31628 26390 31680
rect 33962 31628 33968 31680
rect 34020 31668 34026 31680
rect 34701 31671 34759 31677
rect 34701 31668 34713 31671
rect 34020 31640 34713 31668
rect 34020 31628 34026 31640
rect 34701 31637 34713 31640
rect 34747 31637 34759 31671
rect 34701 31631 34759 31637
rect 36446 31628 36452 31680
rect 36504 31628 36510 31680
rect 38010 31628 38016 31680
rect 38068 31668 38074 31680
rect 38197 31671 38255 31677
rect 38197 31668 38209 31671
rect 38068 31640 38209 31668
rect 38068 31628 38074 31640
rect 38197 31637 38209 31640
rect 38243 31637 38255 31671
rect 38197 31631 38255 31637
rect 38841 31671 38899 31677
rect 38841 31637 38853 31671
rect 38887 31668 38899 31671
rect 39482 31668 39488 31680
rect 38887 31640 39488 31668
rect 38887 31637 38899 31640
rect 38841 31631 38899 31637
rect 39482 31628 39488 31640
rect 39540 31628 39546 31680
rect 44542 31628 44548 31680
rect 44600 31628 44606 31680
rect 1104 31578 45172 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 45172 31578
rect 1104 31504 45172 31526
rect 2406 31424 2412 31476
rect 2464 31424 2470 31476
rect 4062 31424 4068 31476
rect 4120 31464 4126 31476
rect 9217 31467 9275 31473
rect 4120 31436 9076 31464
rect 4120 31424 4126 31436
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 2424 31328 2452 31424
rect 4890 31396 4896 31408
rect 4002 31368 4896 31396
rect 4890 31356 4896 31368
rect 4948 31356 4954 31408
rect 8849 31399 8907 31405
rect 8849 31396 8861 31399
rect 8404 31368 8861 31396
rect 2179 31300 2452 31328
rect 7929 31331 7987 31337
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 7929 31297 7941 31331
rect 7975 31297 7987 31331
rect 7929 31291 7987 31297
rect 1486 31220 1492 31272
rect 1544 31260 1550 31272
rect 2498 31260 2504 31272
rect 1544 31232 2504 31260
rect 1544 31220 1550 31232
rect 2498 31220 2504 31232
rect 2556 31220 2562 31272
rect 2774 31220 2780 31272
rect 2832 31220 2838 31272
rect 3418 31220 3424 31272
rect 3476 31260 3482 31272
rect 6454 31260 6460 31272
rect 3476 31232 6460 31260
rect 3476 31220 3482 31232
rect 6454 31220 6460 31232
rect 6512 31220 6518 31272
rect 7834 31220 7840 31272
rect 7892 31220 7898 31272
rect 7944 31260 7972 31291
rect 8294 31288 8300 31340
rect 8352 31328 8358 31340
rect 8404 31337 8432 31368
rect 8849 31365 8861 31368
rect 8895 31365 8907 31399
rect 8849 31359 8907 31365
rect 9048 31340 9076 31436
rect 9217 31433 9229 31467
rect 9263 31464 9275 31467
rect 9306 31464 9312 31476
rect 9263 31436 9312 31464
rect 9263 31433 9275 31436
rect 9217 31427 9275 31433
rect 9306 31424 9312 31436
rect 9364 31424 9370 31476
rect 9674 31424 9680 31476
rect 9732 31424 9738 31476
rect 9953 31467 10011 31473
rect 9953 31433 9965 31467
rect 9999 31464 10011 31467
rect 10226 31464 10232 31476
rect 9999 31436 10232 31464
rect 9999 31433 10011 31436
rect 9953 31427 10011 31433
rect 10226 31424 10232 31436
rect 10284 31424 10290 31476
rect 10318 31424 10324 31476
rect 10376 31464 10382 31476
rect 10505 31467 10563 31473
rect 10505 31464 10517 31467
rect 10376 31436 10517 31464
rect 10376 31424 10382 31436
rect 10505 31433 10517 31436
rect 10551 31433 10563 31467
rect 13354 31464 13360 31476
rect 10505 31427 10563 31433
rect 12452 31436 13360 31464
rect 9585 31399 9643 31405
rect 9585 31365 9597 31399
rect 9631 31365 9643 31399
rect 9692 31396 9720 31424
rect 9692 31368 9996 31396
rect 9585 31359 9643 31365
rect 8389 31331 8447 31337
rect 8389 31328 8401 31331
rect 8352 31300 8401 31328
rect 8352 31288 8358 31300
rect 8389 31297 8401 31300
rect 8435 31297 8447 31331
rect 8389 31291 8447 31297
rect 8573 31331 8631 31337
rect 8573 31297 8585 31331
rect 8619 31328 8631 31331
rect 8662 31328 8668 31340
rect 8619 31300 8668 31328
rect 8619 31297 8631 31300
rect 8573 31291 8631 31297
rect 8662 31288 8668 31300
rect 8720 31288 8726 31340
rect 8938 31288 8944 31340
rect 8996 31288 9002 31340
rect 9030 31288 9036 31340
rect 9088 31288 9094 31340
rect 9490 31328 9496 31340
rect 9140 31300 9496 31328
rect 8956 31260 8984 31288
rect 7944 31232 8984 31260
rect 9140 31192 9168 31300
rect 9490 31288 9496 31300
rect 9548 31288 9554 31340
rect 9600 31272 9628 31359
rect 9769 31331 9827 31337
rect 9769 31297 9781 31331
rect 9815 31297 9827 31331
rect 9968 31328 9996 31368
rect 10042 31356 10048 31408
rect 10100 31356 10106 31408
rect 12452 31405 12480 31436
rect 13354 31424 13360 31436
rect 13412 31464 13418 31476
rect 14642 31464 14648 31476
rect 13412 31436 14648 31464
rect 13412 31424 13418 31436
rect 14642 31424 14648 31436
rect 14700 31424 14706 31476
rect 17770 31424 17776 31476
rect 17828 31464 17834 31476
rect 18233 31467 18291 31473
rect 18233 31464 18245 31467
rect 17828 31436 18245 31464
rect 17828 31424 17834 31436
rect 18233 31433 18245 31436
rect 18279 31433 18291 31467
rect 18233 31427 18291 31433
rect 21266 31424 21272 31476
rect 21324 31424 21330 31476
rect 21542 31424 21548 31476
rect 21600 31424 21606 31476
rect 22278 31464 22284 31476
rect 21652 31436 22284 31464
rect 10689 31399 10747 31405
rect 10689 31396 10701 31399
rect 10152 31368 10701 31396
rect 10152 31328 10180 31368
rect 10689 31365 10701 31368
rect 10735 31365 10747 31399
rect 10689 31359 10747 31365
rect 12437 31399 12495 31405
rect 12437 31365 12449 31399
rect 12483 31365 12495 31399
rect 13814 31396 13820 31408
rect 12437 31359 12495 31365
rect 13096 31368 13820 31396
rect 13096 31340 13124 31368
rect 13814 31356 13820 31368
rect 13872 31396 13878 31408
rect 15105 31399 15163 31405
rect 15105 31396 15117 31399
rect 13872 31368 15117 31396
rect 13872 31356 13878 31368
rect 15105 31365 15117 31368
rect 15151 31365 15163 31399
rect 15105 31359 15163 31365
rect 15197 31399 15255 31405
rect 15197 31365 15209 31399
rect 15243 31396 15255 31399
rect 15657 31399 15715 31405
rect 15657 31396 15669 31399
rect 15243 31368 15669 31396
rect 15243 31365 15255 31368
rect 15197 31359 15255 31365
rect 15657 31365 15669 31368
rect 15703 31365 15715 31399
rect 15657 31359 15715 31365
rect 19797 31399 19855 31405
rect 19797 31365 19809 31399
rect 19843 31396 19855 31399
rect 20070 31396 20076 31408
rect 19843 31368 20076 31396
rect 19843 31365 19855 31368
rect 19797 31359 19855 31365
rect 20070 31356 20076 31368
rect 20128 31356 20134 31408
rect 21652 31396 21680 31436
rect 22278 31424 22284 31436
rect 22336 31464 22342 31476
rect 22336 31436 22508 31464
rect 22336 31424 22342 31436
rect 21560 31368 21680 31396
rect 9968 31300 10180 31328
rect 9769 31291 9827 31297
rect 9582 31220 9588 31272
rect 9640 31220 9646 31272
rect 4264 31164 9168 31192
rect 1854 31084 1860 31136
rect 1912 31124 1918 31136
rect 1949 31127 2007 31133
rect 1949 31124 1961 31127
rect 1912 31096 1961 31124
rect 1912 31084 1918 31096
rect 1949 31093 1961 31096
rect 1995 31093 2007 31127
rect 1949 31087 2007 31093
rect 4062 31084 4068 31136
rect 4120 31124 4126 31136
rect 4264 31133 4292 31164
rect 9398 31152 9404 31204
rect 9456 31192 9462 31204
rect 9784 31192 9812 31291
rect 10226 31288 10232 31340
rect 10284 31328 10290 31340
rect 10321 31331 10379 31337
rect 10321 31328 10333 31331
rect 10284 31300 10333 31328
rect 10284 31288 10290 31300
rect 10321 31297 10333 31300
rect 10367 31328 10379 31331
rect 10502 31328 10508 31340
rect 10367 31300 10508 31328
rect 10367 31297 10379 31300
rect 10321 31291 10379 31297
rect 10502 31288 10508 31300
rect 10560 31288 10566 31340
rect 10597 31331 10655 31337
rect 10597 31297 10609 31331
rect 10643 31297 10655 31331
rect 10597 31291 10655 31297
rect 10781 31331 10839 31337
rect 10781 31297 10793 31331
rect 10827 31297 10839 31331
rect 10781 31291 10839 31297
rect 9858 31220 9864 31272
rect 9916 31260 9922 31272
rect 10137 31263 10195 31269
rect 10137 31260 10149 31263
rect 9916 31232 10149 31260
rect 9916 31220 9922 31232
rect 10137 31229 10149 31232
rect 10183 31229 10195 31263
rect 10612 31260 10640 31291
rect 10137 31223 10195 31229
rect 10419 31232 10640 31260
rect 9456 31164 9812 31192
rect 9456 31152 9462 31164
rect 4249 31127 4307 31133
rect 4249 31124 4261 31127
rect 4120 31096 4261 31124
rect 4120 31084 4126 31096
rect 4249 31093 4261 31096
rect 4295 31093 4307 31127
rect 4249 31087 4307 31093
rect 8294 31084 8300 31136
rect 8352 31084 8358 31136
rect 8389 31127 8447 31133
rect 8389 31093 8401 31127
rect 8435 31124 8447 31127
rect 10321 31127 10379 31133
rect 10321 31124 10333 31127
rect 8435 31096 10333 31124
rect 8435 31093 8447 31096
rect 8389 31087 8447 31093
rect 10321 31093 10333 31096
rect 10367 31124 10379 31127
rect 10419 31124 10447 31232
rect 10367 31096 10447 31124
rect 10367 31093 10379 31096
rect 10321 31087 10379 31093
rect 10502 31084 10508 31136
rect 10560 31124 10566 31136
rect 10796 31124 10824 31291
rect 10870 31288 10876 31340
rect 10928 31328 10934 31340
rect 12342 31337 12348 31340
rect 12161 31331 12219 31337
rect 12161 31328 12173 31331
rect 10928 31300 12173 31328
rect 10928 31288 10934 31300
rect 12161 31297 12173 31300
rect 12207 31297 12219 31331
rect 12161 31291 12219 31297
rect 12309 31331 12348 31337
rect 12309 31297 12321 31331
rect 12309 31291 12348 31297
rect 12342 31288 12348 31291
rect 12400 31288 12406 31340
rect 12526 31288 12532 31340
rect 12584 31288 12590 31340
rect 12626 31331 12684 31337
rect 12626 31297 12638 31331
rect 12672 31297 12684 31331
rect 12626 31291 12684 31297
rect 12434 31152 12440 31204
rect 12492 31192 12498 31204
rect 12636 31192 12664 31291
rect 13078 31288 13084 31340
rect 13136 31288 13142 31340
rect 14734 31288 14740 31340
rect 14792 31288 14798 31340
rect 14826 31288 14832 31340
rect 14884 31288 14890 31340
rect 14922 31331 14980 31337
rect 14922 31297 14934 31331
rect 14968 31297 14980 31331
rect 14922 31291 14980 31297
rect 15335 31331 15393 31337
rect 15335 31297 15347 31331
rect 15381 31328 15393 31331
rect 15562 31328 15568 31340
rect 15381 31300 15568 31328
rect 15381 31297 15393 31300
rect 15335 31291 15393 31297
rect 12802 31220 12808 31272
rect 12860 31220 12866 31272
rect 12986 31220 12992 31272
rect 13044 31260 13050 31272
rect 14936 31260 14964 31291
rect 15562 31288 15568 31300
rect 15620 31288 15626 31340
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 15672 31300 15761 31328
rect 13044 31232 14964 31260
rect 13044 31220 13050 31232
rect 15470 31220 15476 31272
rect 15528 31220 15534 31272
rect 12492 31164 12664 31192
rect 12820 31192 12848 31220
rect 12820 31164 13492 31192
rect 12492 31152 12498 31164
rect 10560 31096 10824 31124
rect 10560 31084 10566 31096
rect 12802 31084 12808 31136
rect 12860 31084 12866 31136
rect 12894 31084 12900 31136
rect 12952 31124 12958 31136
rect 13170 31124 13176 31136
rect 12952 31096 13176 31124
rect 12952 31084 12958 31096
rect 13170 31084 13176 31096
rect 13228 31084 13234 31136
rect 13464 31133 13492 31164
rect 13814 31152 13820 31204
rect 13872 31192 13878 31204
rect 14090 31192 14096 31204
rect 13872 31164 14096 31192
rect 13872 31152 13878 31164
rect 14090 31152 14096 31164
rect 14148 31152 14154 31204
rect 15488 31192 15516 31220
rect 15304 31164 15516 31192
rect 13449 31127 13507 31133
rect 13449 31093 13461 31127
rect 13495 31124 13507 31127
rect 14734 31124 14740 31136
rect 13495 31096 14740 31124
rect 13495 31093 13507 31096
rect 13449 31087 13507 31093
rect 14734 31084 14740 31096
rect 14792 31124 14798 31136
rect 15304 31124 15332 31164
rect 15672 31136 15700 31300
rect 15749 31297 15761 31300
rect 15795 31328 15807 31331
rect 16206 31328 16212 31340
rect 15795 31300 16212 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 16206 31288 16212 31300
rect 16264 31288 16270 31340
rect 18322 31288 18328 31340
rect 18380 31288 18386 31340
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 21560 31328 21588 31368
rect 22094 31356 22100 31408
rect 22152 31356 22158 31408
rect 22480 31396 22508 31436
rect 23658 31424 23664 31476
rect 23716 31424 23722 31476
rect 24118 31424 24124 31476
rect 24176 31424 24182 31476
rect 25958 31424 25964 31476
rect 26016 31424 26022 31476
rect 26694 31424 26700 31476
rect 26752 31464 26758 31476
rect 27157 31467 27215 31473
rect 27157 31464 27169 31467
rect 26752 31436 27169 31464
rect 26752 31424 26758 31436
rect 27157 31433 27169 31436
rect 27203 31433 27215 31467
rect 27157 31427 27215 31433
rect 27525 31467 27583 31473
rect 27525 31433 27537 31467
rect 27571 31464 27583 31467
rect 28626 31464 28632 31476
rect 27571 31436 28632 31464
rect 27571 31433 27583 31436
rect 27525 31427 27583 31433
rect 28626 31424 28632 31436
rect 28684 31424 28690 31476
rect 29822 31424 29828 31476
rect 29880 31424 29886 31476
rect 32306 31424 32312 31476
rect 32364 31424 32370 31476
rect 32490 31424 32496 31476
rect 32548 31464 32554 31476
rect 32861 31467 32919 31473
rect 32861 31464 32873 31467
rect 32548 31436 32873 31464
rect 32548 31424 32554 31436
rect 32861 31433 32873 31436
rect 32907 31433 32919 31467
rect 33870 31464 33876 31476
rect 32861 31427 32919 31433
rect 33704 31436 33876 31464
rect 24762 31405 24768 31408
rect 22480 31368 22586 31396
rect 24756 31359 24768 31405
rect 24762 31356 24768 31359
rect 24820 31356 24826 31408
rect 29914 31356 29920 31408
rect 29972 31356 29978 31408
rect 32508 31368 32996 31396
rect 20864 31300 21588 31328
rect 21637 31331 21695 31337
rect 20864 31288 20870 31300
rect 21637 31297 21649 31331
rect 21683 31297 21695 31331
rect 21637 31291 21695 31297
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 26786 31328 26792 31340
rect 26375 31300 26792 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 19150 31220 19156 31272
rect 19208 31260 19214 31272
rect 19521 31263 19579 31269
rect 19521 31260 19533 31263
rect 19208 31232 19533 31260
rect 19208 31220 19214 31232
rect 19521 31229 19533 31232
rect 19567 31229 19579 31263
rect 19521 31223 19579 31229
rect 14792 31096 15332 31124
rect 14792 31084 14798 31096
rect 15470 31084 15476 31136
rect 15528 31084 15534 31136
rect 15654 31084 15660 31136
rect 15712 31084 15718 31136
rect 21652 31124 21680 31291
rect 21818 31220 21824 31272
rect 21876 31220 21882 31272
rect 23569 31263 23627 31269
rect 23569 31260 23581 31263
rect 21928 31232 23581 31260
rect 21928 31124 21956 31232
rect 23569 31229 23581 31232
rect 23615 31260 23627 31263
rect 24044 31260 24072 31291
rect 26786 31288 26792 31300
rect 26844 31288 26850 31340
rect 29362 31288 29368 31340
rect 29420 31328 29426 31340
rect 29641 31331 29699 31337
rect 29641 31328 29653 31331
rect 29420 31300 29653 31328
rect 29420 31288 29426 31300
rect 29641 31297 29653 31300
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 29825 31331 29883 31337
rect 29825 31297 29837 31331
rect 29871 31328 29883 31331
rect 29932 31328 29960 31356
rect 32508 31337 32536 31368
rect 32968 31337 32996 31368
rect 29871 31300 29960 31328
rect 32493 31331 32551 31337
rect 29871 31297 29883 31300
rect 29825 31291 29883 31297
rect 32493 31297 32505 31331
rect 32539 31297 32551 31331
rect 32493 31291 32551 31297
rect 32677 31331 32735 31337
rect 32677 31297 32689 31331
rect 32723 31328 32735 31331
rect 32769 31331 32827 31337
rect 32769 31328 32781 31331
rect 32723 31300 32781 31328
rect 32723 31297 32735 31300
rect 32677 31291 32735 31297
rect 32769 31297 32781 31300
rect 32815 31297 32827 31331
rect 32769 31291 32827 31297
rect 32953 31331 33011 31337
rect 32953 31297 32965 31331
rect 32999 31297 33011 31331
rect 32953 31291 33011 31297
rect 23615 31232 24072 31260
rect 23615 31229 23627 31232
rect 23569 31223 23627 31229
rect 24210 31220 24216 31272
rect 24268 31220 24274 31272
rect 24489 31263 24547 31269
rect 24489 31229 24501 31263
rect 24535 31229 24547 31263
rect 24489 31223 24547 31229
rect 21652 31096 21956 31124
rect 24504 31124 24532 31223
rect 26234 31220 26240 31272
rect 26292 31220 26298 31272
rect 26418 31220 26424 31272
rect 26476 31220 26482 31272
rect 26510 31220 26516 31272
rect 26568 31220 26574 31272
rect 27062 31220 27068 31272
rect 27120 31260 27126 31272
rect 27617 31263 27675 31269
rect 27617 31260 27629 31263
rect 27120 31232 27629 31260
rect 27120 31220 27126 31232
rect 27617 31229 27629 31232
rect 27663 31229 27675 31263
rect 27617 31223 27675 31229
rect 27709 31263 27767 31269
rect 27709 31229 27721 31263
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 25869 31195 25927 31201
rect 25869 31161 25881 31195
rect 25915 31192 25927 31195
rect 26252 31192 26280 31220
rect 25915 31164 26280 31192
rect 25915 31161 25927 31164
rect 25869 31155 25927 31161
rect 27522 31152 27528 31204
rect 27580 31192 27586 31204
rect 27724 31192 27752 31223
rect 30098 31220 30104 31272
rect 30156 31260 30162 31272
rect 32692 31260 32720 31291
rect 30156 31232 32720 31260
rect 30156 31220 30162 31232
rect 27580 31164 27752 31192
rect 27580 31152 27586 31164
rect 24762 31124 24768 31136
rect 24504 31096 24768 31124
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 32968 31124 32996 31291
rect 33502 31288 33508 31340
rect 33560 31288 33566 31340
rect 33594 31288 33600 31340
rect 33652 31328 33658 31340
rect 33704 31337 33732 31436
rect 33870 31424 33876 31436
rect 33928 31424 33934 31476
rect 33962 31424 33968 31476
rect 34020 31424 34026 31476
rect 34057 31467 34115 31473
rect 34057 31433 34069 31467
rect 34103 31433 34115 31467
rect 34057 31427 34115 31433
rect 33781 31399 33839 31405
rect 33781 31365 33793 31399
rect 33827 31396 33839 31399
rect 33980 31396 34008 31424
rect 33827 31368 34008 31396
rect 34072 31396 34100 31427
rect 39482 31424 39488 31476
rect 39540 31424 39546 31476
rect 42518 31424 42524 31476
rect 42576 31464 42582 31476
rect 42613 31467 42671 31473
rect 42613 31464 42625 31467
rect 42576 31436 42625 31464
rect 42576 31424 42582 31436
rect 42613 31433 42625 31436
rect 42659 31433 42671 31467
rect 42613 31427 42671 31433
rect 43073 31467 43131 31473
rect 43073 31433 43085 31467
rect 43119 31464 43131 31467
rect 43254 31464 43260 31476
rect 43119 31436 43260 31464
rect 43119 31433 43131 31436
rect 43073 31427 43131 31433
rect 43254 31424 43260 31436
rect 43312 31424 43318 31476
rect 34425 31399 34483 31405
rect 34425 31396 34437 31399
rect 34072 31368 34437 31396
rect 33827 31365 33839 31368
rect 33781 31359 33839 31365
rect 34425 31365 34437 31368
rect 34471 31365 34483 31399
rect 34425 31359 34483 31365
rect 38010 31356 38016 31408
rect 38068 31356 38074 31408
rect 43346 31356 43352 31408
rect 43404 31396 43410 31408
rect 43404 31368 43668 31396
rect 43404 31356 43410 31368
rect 33689 31331 33747 31337
rect 33689 31328 33701 31331
rect 33652 31300 33701 31328
rect 33652 31288 33658 31300
rect 33689 31297 33701 31300
rect 33735 31297 33747 31331
rect 33689 31291 33747 31297
rect 33873 31331 33931 31337
rect 33873 31297 33885 31331
rect 33919 31328 33931 31331
rect 34054 31328 34060 31340
rect 33919 31300 34060 31328
rect 33919 31297 33931 31300
rect 33873 31291 33931 31297
rect 34054 31288 34060 31300
rect 34112 31288 34118 31340
rect 35526 31288 35532 31340
rect 35584 31328 35590 31340
rect 36354 31328 36360 31340
rect 35584 31300 36360 31328
rect 35584 31288 35590 31300
rect 36354 31288 36360 31300
rect 36412 31288 36418 31340
rect 37734 31288 37740 31340
rect 37792 31288 37798 31340
rect 39114 31288 39120 31340
rect 39172 31288 39178 31340
rect 43640 31337 43668 31368
rect 42981 31331 43039 31337
rect 42981 31297 42993 31331
rect 43027 31328 43039 31331
rect 43625 31331 43683 31337
rect 43027 31300 43576 31328
rect 43027 31297 43039 31300
rect 42981 31291 43039 31297
rect 43548 31272 43576 31300
rect 43625 31297 43637 31331
rect 43671 31297 43683 31331
rect 43625 31291 43683 31297
rect 43898 31288 43904 31340
rect 43956 31288 43962 31340
rect 44542 31288 44548 31340
rect 44600 31288 44606 31340
rect 34149 31263 34207 31269
rect 34149 31229 34161 31263
rect 34195 31229 34207 31263
rect 34149 31223 34207 31229
rect 33042 31152 33048 31204
rect 33100 31192 33106 31204
rect 34164 31192 34192 31223
rect 42886 31220 42892 31272
rect 42944 31260 42950 31272
rect 43165 31263 43223 31269
rect 43165 31260 43177 31263
rect 42944 31232 43177 31260
rect 42944 31220 42950 31232
rect 43165 31229 43177 31232
rect 43211 31229 43223 31263
rect 43165 31223 43223 31229
rect 43530 31220 43536 31272
rect 43588 31260 43594 31272
rect 43588 31232 43852 31260
rect 43588 31220 43594 31232
rect 33100 31164 34192 31192
rect 33100 31152 33106 31164
rect 33870 31124 33876 31136
rect 32968 31096 33876 31124
rect 33870 31084 33876 31096
rect 33928 31084 33934 31136
rect 34164 31124 34192 31164
rect 35434 31152 35440 31204
rect 35492 31192 35498 31204
rect 35897 31195 35955 31201
rect 35897 31192 35909 31195
rect 35492 31164 35909 31192
rect 35492 31152 35498 31164
rect 35897 31161 35909 31164
rect 35943 31161 35955 31195
rect 35897 31155 35955 31161
rect 43070 31152 43076 31204
rect 43128 31192 43134 31204
rect 43824 31201 43852 31232
rect 43717 31195 43775 31201
rect 43717 31192 43729 31195
rect 43128 31164 43729 31192
rect 43128 31152 43134 31164
rect 43717 31161 43729 31164
rect 43763 31161 43775 31195
rect 43717 31155 43775 31161
rect 43809 31195 43867 31201
rect 43809 31161 43821 31195
rect 43855 31192 43867 31195
rect 44560 31192 44588 31288
rect 43855 31164 44588 31192
rect 43855 31161 43867 31164
rect 43809 31155 43867 31161
rect 35618 31124 35624 31136
rect 34164 31096 35624 31124
rect 35618 31084 35624 31096
rect 35676 31084 35682 31136
rect 43438 31084 43444 31136
rect 43496 31084 43502 31136
rect 1104 31034 45172 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 45172 31034
rect 1104 30960 45172 30982
rect 2774 30880 2780 30932
rect 2832 30920 2838 30932
rect 3329 30923 3387 30929
rect 3329 30920 3341 30923
rect 2832 30892 3341 30920
rect 2832 30880 2838 30892
rect 3329 30889 3341 30892
rect 3375 30889 3387 30923
rect 3329 30883 3387 30889
rect 3712 30892 3924 30920
rect 3234 30812 3240 30864
rect 3292 30852 3298 30864
rect 3712 30852 3740 30892
rect 3292 30824 3740 30852
rect 3789 30855 3847 30861
rect 3292 30812 3298 30824
rect 3789 30821 3801 30855
rect 3835 30821 3847 30855
rect 3789 30815 3847 30821
rect 1486 30744 1492 30796
rect 1544 30744 1550 30796
rect 1765 30787 1823 30793
rect 1765 30753 1777 30787
rect 1811 30784 1823 30787
rect 1854 30784 1860 30796
rect 1811 30756 1860 30784
rect 1811 30753 1823 30756
rect 1765 30747 1823 30753
rect 1854 30744 1860 30756
rect 1912 30744 1918 30796
rect 3418 30716 3424 30728
rect 2898 30688 3424 30716
rect 3418 30676 3424 30688
rect 3476 30676 3482 30728
rect 3513 30719 3571 30725
rect 3513 30685 3525 30719
rect 3559 30716 3571 30719
rect 3804 30716 3832 30815
rect 3559 30688 3832 30716
rect 3896 30716 3924 30892
rect 4614 30880 4620 30932
rect 4672 30880 4678 30932
rect 8938 30880 8944 30932
rect 8996 30920 9002 30932
rect 9306 30920 9312 30932
rect 8996 30892 9312 30920
rect 8996 30880 9002 30892
rect 9306 30880 9312 30892
rect 9364 30880 9370 30932
rect 9398 30880 9404 30932
rect 9456 30880 9462 30932
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 12621 30923 12679 30929
rect 12621 30920 12633 30923
rect 11940 30892 12633 30920
rect 11940 30880 11946 30892
rect 12621 30889 12633 30892
rect 12667 30889 12679 30923
rect 12621 30883 12679 30889
rect 12802 30880 12808 30932
rect 12860 30920 12866 30932
rect 13357 30923 13415 30929
rect 13357 30920 13369 30923
rect 12860 30892 13369 30920
rect 12860 30880 12866 30892
rect 13357 30889 13369 30892
rect 13403 30889 13415 30923
rect 13357 30883 13415 30889
rect 13446 30880 13452 30932
rect 13504 30920 13510 30932
rect 13504 30892 13768 30920
rect 13504 30880 13510 30892
rect 4433 30787 4491 30793
rect 4433 30753 4445 30787
rect 4479 30784 4491 30787
rect 4632 30784 4660 30880
rect 8294 30812 8300 30864
rect 8352 30852 8358 30864
rect 10870 30852 10876 30864
rect 8352 30824 10876 30852
rect 8352 30812 8358 30824
rect 10870 30812 10876 30824
rect 10928 30812 10934 30864
rect 11238 30812 11244 30864
rect 11296 30812 11302 30864
rect 13538 30852 13544 30864
rect 12728 30824 13544 30852
rect 4479 30756 4660 30784
rect 4479 30753 4491 30756
rect 4433 30747 4491 30753
rect 9030 30744 9036 30796
rect 9088 30784 9094 30796
rect 9088 30756 9168 30784
rect 9088 30744 9094 30756
rect 4617 30719 4675 30725
rect 4617 30716 4629 30719
rect 3896 30688 4629 30716
rect 3559 30685 3571 30688
rect 3513 30679 3571 30685
rect 4617 30685 4629 30688
rect 4663 30685 4675 30719
rect 4617 30679 4675 30685
rect 5166 30676 5172 30728
rect 5224 30676 5230 30728
rect 8938 30676 8944 30728
rect 8996 30725 9002 30728
rect 9140 30725 9168 30756
rect 9490 30744 9496 30796
rect 9548 30784 9554 30796
rect 10045 30787 10103 30793
rect 10045 30784 10057 30787
rect 9548 30756 9720 30784
rect 9548 30744 9554 30756
rect 8996 30716 9005 30725
rect 9125 30719 9183 30725
rect 8996 30688 9041 30716
rect 8996 30679 9005 30688
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 8996 30676 9002 30679
rect 9582 30676 9588 30728
rect 9640 30676 9646 30728
rect 9692 30725 9720 30756
rect 9784 30756 10057 30784
rect 9784 30728 9812 30756
rect 10045 30753 10057 30756
rect 10091 30784 10103 30787
rect 11256 30784 11284 30812
rect 12069 30787 12127 30793
rect 12069 30784 12081 30787
rect 10091 30756 10364 30784
rect 11256 30756 11468 30784
rect 10091 30753 10103 30756
rect 10045 30747 10103 30753
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30685 9735 30719
rect 9677 30679 9735 30685
rect 9766 30676 9772 30728
rect 9824 30676 9830 30728
rect 10137 30719 10195 30725
rect 10137 30716 10149 30719
rect 9968 30688 10149 30716
rect 3786 30608 3792 30660
rect 3844 30648 3850 30660
rect 9968 30657 9996 30688
rect 10137 30685 10149 30688
rect 10183 30685 10195 30719
rect 10137 30679 10195 30685
rect 10226 30676 10232 30728
rect 10284 30676 10290 30728
rect 10336 30725 10364 30756
rect 10321 30719 10379 30725
rect 10321 30685 10333 30719
rect 10367 30716 10379 30719
rect 10873 30719 10931 30725
rect 10873 30716 10885 30719
rect 10367 30688 10885 30716
rect 10367 30685 10379 30688
rect 10321 30679 10379 30685
rect 10873 30685 10885 30688
rect 10919 30685 10931 30719
rect 10873 30679 10931 30685
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 11440 30725 11468 30756
rect 11532 30756 12081 30784
rect 11287 30719 11345 30725
rect 11287 30716 11299 30719
rect 11112 30688 11299 30716
rect 11112 30676 11118 30688
rect 11287 30685 11299 30688
rect 11333 30685 11345 30719
rect 11287 30679 11345 30685
rect 11425 30719 11483 30725
rect 11425 30685 11437 30719
rect 11471 30685 11483 30719
rect 11425 30679 11483 30685
rect 11532 30657 11560 30756
rect 12069 30753 12081 30756
rect 12115 30753 12127 30787
rect 12069 30747 12127 30753
rect 11645 30719 11703 30725
rect 11645 30716 11657 30719
rect 11624 30685 11657 30716
rect 11691 30685 11703 30719
rect 11624 30679 11703 30685
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30716 11851 30719
rect 11882 30716 11888 30728
rect 11839 30688 11888 30716
rect 11839 30685 11851 30688
rect 11793 30679 11851 30685
rect 4249 30651 4307 30657
rect 4249 30648 4261 30651
rect 3844 30620 4261 30648
rect 3844 30608 3850 30620
rect 4249 30617 4261 30620
rect 4295 30617 4307 30651
rect 4249 30611 4307 30617
rect 4709 30651 4767 30657
rect 4709 30617 4721 30651
rect 4755 30648 4767 30651
rect 9953 30651 10011 30657
rect 9953 30648 9965 30651
rect 4755 30620 9965 30648
rect 4755 30617 4767 30620
rect 4709 30611 4767 30617
rect 9953 30617 9965 30620
rect 9999 30617 10011 30651
rect 9953 30611 10011 30617
rect 10965 30651 11023 30657
rect 10965 30617 10977 30651
rect 11011 30648 11023 30651
rect 11517 30651 11575 30657
rect 11517 30648 11529 30651
rect 11011 30620 11529 30648
rect 11011 30617 11023 30620
rect 10965 30611 11023 30617
rect 11517 30617 11529 30620
rect 11563 30617 11575 30651
rect 11517 30611 11575 30617
rect 11624 30648 11652 30679
rect 11882 30676 11888 30688
rect 11940 30676 11946 30728
rect 12161 30718 12219 30724
rect 11992 30690 12173 30718
rect 11992 30648 12020 30690
rect 12161 30684 12173 30690
rect 12207 30684 12219 30718
rect 12161 30678 12219 30684
rect 12250 30676 12256 30728
rect 12308 30718 12314 30728
rect 12437 30719 12495 30725
rect 12308 30716 12388 30718
rect 12437 30716 12449 30719
rect 12308 30690 12449 30716
rect 12308 30676 12314 30690
rect 12360 30688 12449 30690
rect 12437 30685 12449 30688
rect 12483 30685 12495 30719
rect 12437 30679 12495 30685
rect 12529 30719 12587 30725
rect 12529 30685 12541 30719
rect 12575 30716 12587 30719
rect 12728 30716 12756 30824
rect 13538 30812 13544 30824
rect 13596 30812 13602 30864
rect 12802 30744 12808 30796
rect 12860 30744 12866 30796
rect 13170 30744 13176 30796
rect 13228 30744 13234 30796
rect 12575 30688 12756 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 12894 30676 12900 30728
rect 12952 30676 12958 30728
rect 13357 30719 13415 30725
rect 13357 30716 13369 30719
rect 13004 30688 13369 30716
rect 13004 30648 13032 30688
rect 13357 30685 13369 30688
rect 13403 30685 13415 30719
rect 13357 30679 13415 30685
rect 13541 30719 13599 30725
rect 13541 30685 13553 30719
rect 13587 30685 13599 30719
rect 13541 30679 13599 30685
rect 11624 30620 12020 30648
rect 12452 30620 13032 30648
rect 13265 30651 13323 30657
rect 4154 30540 4160 30592
rect 4212 30540 4218 30592
rect 4798 30540 4804 30592
rect 4856 30580 4862 30592
rect 4985 30583 5043 30589
rect 4985 30580 4997 30583
rect 4856 30552 4997 30580
rect 4856 30540 4862 30552
rect 4985 30549 4997 30552
rect 5031 30549 5043 30583
rect 4985 30543 5043 30549
rect 9033 30583 9091 30589
rect 9033 30549 9045 30583
rect 9079 30580 9091 30583
rect 9858 30580 9864 30592
rect 9079 30552 9864 30580
rect 9079 30549 9091 30552
rect 9033 30543 9091 30549
rect 9858 30540 9864 30552
rect 9916 30540 9922 30592
rect 11146 30540 11152 30592
rect 11204 30540 11210 30592
rect 11330 30540 11336 30592
rect 11388 30580 11394 30592
rect 11624 30580 11652 30620
rect 11388 30552 11652 30580
rect 11885 30583 11943 30589
rect 11388 30540 11394 30552
rect 11885 30549 11897 30583
rect 11931 30580 11943 30583
rect 12452 30580 12480 30620
rect 13265 30617 13277 30651
rect 13311 30617 13323 30651
rect 13556 30648 13584 30679
rect 13630 30676 13636 30728
rect 13688 30676 13694 30728
rect 13740 30716 13768 30892
rect 13906 30880 13912 30932
rect 13964 30920 13970 30932
rect 14231 30923 14289 30929
rect 14231 30920 14243 30923
rect 13964 30892 14243 30920
rect 13964 30880 13970 30892
rect 14231 30889 14243 30892
rect 14277 30889 14289 30923
rect 14231 30883 14289 30889
rect 14369 30923 14427 30929
rect 14369 30889 14381 30923
rect 14415 30920 14427 30923
rect 15470 30920 15476 30932
rect 14415 30892 15476 30920
rect 14415 30889 14427 30892
rect 14369 30883 14427 30889
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 16482 30880 16488 30932
rect 16540 30920 16546 30932
rect 18230 30920 18236 30932
rect 16540 30892 18236 30920
rect 16540 30880 16546 30892
rect 18230 30880 18236 30892
rect 18288 30920 18294 30932
rect 18417 30923 18475 30929
rect 18417 30920 18429 30923
rect 18288 30892 18429 30920
rect 18288 30880 18294 30892
rect 18417 30889 18429 30892
rect 18463 30889 18475 30923
rect 18417 30883 18475 30889
rect 19334 30880 19340 30932
rect 19392 30880 19398 30932
rect 21542 30880 21548 30932
rect 21600 30920 21606 30932
rect 21818 30920 21824 30932
rect 21600 30892 21824 30920
rect 21600 30880 21606 30892
rect 21818 30880 21824 30892
rect 21876 30920 21882 30932
rect 22281 30923 22339 30929
rect 22281 30920 22293 30923
rect 21876 30892 22293 30920
rect 21876 30880 21882 30892
rect 22281 30889 22293 30892
rect 22327 30889 22339 30923
rect 22281 30883 22339 30889
rect 13817 30855 13875 30861
rect 13817 30821 13829 30855
rect 13863 30821 13875 30855
rect 13817 30815 13875 30821
rect 16025 30855 16083 30861
rect 16025 30821 16037 30855
rect 16071 30852 16083 30855
rect 16071 30824 16804 30852
rect 16071 30821 16083 30824
rect 16025 30815 16083 30821
rect 13832 30784 13860 30815
rect 14461 30787 14519 30793
rect 14461 30784 14473 30787
rect 13832 30756 14473 30784
rect 14461 30753 14473 30756
rect 14507 30753 14519 30787
rect 14461 30747 14519 30753
rect 14553 30787 14611 30793
rect 14553 30753 14565 30787
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 14568 30716 14596 30747
rect 16666 30744 16672 30796
rect 16724 30744 16730 30796
rect 16776 30784 16804 30824
rect 16945 30787 17003 30793
rect 16945 30784 16957 30787
rect 16776 30756 16957 30784
rect 16945 30753 16957 30756
rect 16991 30753 17003 30787
rect 16945 30747 17003 30753
rect 15286 30716 15292 30728
rect 13740 30688 15292 30716
rect 15286 30676 15292 30688
rect 15344 30676 15350 30728
rect 15838 30676 15844 30728
rect 15896 30676 15902 30728
rect 16301 30719 16359 30725
rect 16301 30685 16313 30719
rect 16347 30716 16359 30719
rect 16482 30716 16488 30728
rect 16347 30688 16488 30716
rect 16347 30685 16359 30688
rect 16301 30679 16359 30685
rect 16482 30676 16488 30688
rect 16540 30676 16546 30728
rect 16577 30719 16635 30725
rect 16577 30685 16589 30719
rect 16623 30685 16635 30719
rect 16577 30679 16635 30685
rect 18877 30719 18935 30725
rect 18877 30685 18889 30719
rect 18923 30685 18935 30719
rect 19352 30716 19380 30880
rect 22296 30784 22324 30883
rect 26786 30880 26792 30932
rect 26844 30880 26850 30932
rect 30009 30923 30067 30929
rect 30009 30889 30021 30923
rect 30055 30920 30067 30923
rect 30098 30920 30104 30932
rect 30055 30892 30104 30920
rect 30055 30889 30067 30892
rect 30009 30883 30067 30889
rect 30098 30880 30104 30892
rect 30156 30880 30162 30932
rect 33502 30880 33508 30932
rect 33560 30880 33566 30932
rect 33870 30880 33876 30932
rect 33928 30880 33934 30932
rect 43438 30880 43444 30932
rect 43496 30880 43502 30932
rect 26053 30855 26111 30861
rect 26053 30821 26065 30855
rect 26099 30852 26111 30855
rect 43346 30852 43352 30864
rect 26099 30824 26188 30852
rect 26099 30821 26111 30824
rect 26053 30815 26111 30821
rect 26160 30793 26188 30824
rect 38626 30824 43352 30852
rect 22833 30787 22891 30793
rect 22833 30784 22845 30787
rect 22296 30756 22845 30784
rect 22833 30753 22845 30756
rect 22879 30753 22891 30787
rect 22833 30747 22891 30753
rect 26145 30787 26203 30793
rect 26145 30753 26157 30787
rect 26191 30753 26203 30787
rect 26145 30747 26203 30753
rect 27798 30744 27804 30796
rect 27856 30744 27862 30796
rect 29825 30787 29883 30793
rect 29825 30753 29837 30787
rect 29871 30784 29883 30787
rect 30190 30784 30196 30796
rect 29871 30756 30196 30784
rect 29871 30753 29883 30756
rect 29825 30747 29883 30753
rect 30190 30744 30196 30756
rect 30248 30744 30254 30796
rect 33318 30744 33324 30796
rect 33376 30744 33382 30796
rect 35894 30744 35900 30796
rect 35952 30744 35958 30796
rect 36446 30744 36452 30796
rect 36504 30784 36510 30796
rect 37645 30787 37703 30793
rect 37645 30784 37657 30787
rect 36504 30756 37657 30784
rect 36504 30744 36510 30756
rect 37645 30753 37657 30756
rect 37691 30784 37703 30787
rect 38626 30784 38654 30824
rect 43346 30812 43352 30824
rect 43404 30812 43410 30864
rect 37691 30756 38654 30784
rect 37691 30753 37703 30756
rect 37645 30747 37703 30753
rect 40310 30744 40316 30796
rect 40368 30744 40374 30796
rect 42150 30744 42156 30796
rect 42208 30784 42214 30796
rect 42797 30787 42855 30793
rect 42797 30784 42809 30787
rect 42208 30756 42809 30784
rect 42208 30744 42214 30756
rect 42797 30753 42809 30756
rect 42843 30753 42855 30787
rect 42797 30747 42855 30753
rect 43257 30787 43315 30793
rect 43257 30753 43269 30787
rect 43303 30784 43315 30787
rect 43456 30784 43484 30880
rect 43303 30756 43484 30784
rect 43303 30753 43315 30756
rect 43257 30747 43315 30753
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 19352 30688 21005 30716
rect 18877 30679 18935 30685
rect 20993 30685 21005 30688
rect 21039 30716 21051 30719
rect 24673 30719 24731 30725
rect 21039 30688 24348 30716
rect 21039 30685 21051 30688
rect 20993 30679 21051 30685
rect 13906 30648 13912 30660
rect 13556 30620 13912 30648
rect 13265 30611 13323 30617
rect 11931 30552 12480 30580
rect 13280 30580 13308 30611
rect 13906 30608 13912 30620
rect 13964 30608 13970 30660
rect 14090 30608 14096 30660
rect 14148 30608 14154 30660
rect 14826 30608 14832 30660
rect 14884 30648 14890 30660
rect 16592 30648 16620 30679
rect 16666 30648 16672 30660
rect 14884 30620 16672 30648
rect 14884 30608 14890 30620
rect 16666 30608 16672 30620
rect 16724 30608 16730 30660
rect 18230 30648 18236 30660
rect 18170 30620 18236 30648
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 18892 30648 18920 30679
rect 19334 30648 19340 30660
rect 18892 30620 19340 30648
rect 19334 30608 19340 30620
rect 19392 30608 19398 30660
rect 22554 30608 22560 30660
rect 22612 30648 22618 30660
rect 23078 30651 23136 30657
rect 23078 30648 23090 30651
rect 22612 30620 23090 30648
rect 22612 30608 22618 30620
rect 23078 30617 23090 30620
rect 23124 30617 23136 30651
rect 23078 30611 23136 30617
rect 13538 30580 13544 30592
rect 13280 30552 13544 30580
rect 11931 30549 11943 30552
rect 11885 30543 11943 30549
rect 13538 30540 13544 30552
rect 13596 30540 13602 30592
rect 16117 30583 16175 30589
rect 16117 30549 16129 30583
rect 16163 30580 16175 30583
rect 16206 30580 16212 30592
rect 16163 30552 16212 30580
rect 16163 30549 16175 30552
rect 16117 30543 16175 30549
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 16482 30540 16488 30592
rect 16540 30540 16546 30592
rect 19061 30583 19119 30589
rect 19061 30549 19073 30583
rect 19107 30580 19119 30583
rect 19426 30580 19432 30592
rect 19107 30552 19432 30580
rect 19107 30549 19119 30552
rect 19061 30543 19119 30549
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 24210 30540 24216 30592
rect 24268 30540 24274 30592
rect 24320 30580 24348 30688
rect 24673 30685 24685 30719
rect 24719 30716 24731 30719
rect 24762 30716 24768 30728
rect 24719 30688 24768 30716
rect 24719 30685 24731 30688
rect 24673 30679 24731 30685
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 24940 30719 24998 30725
rect 24940 30685 24952 30719
rect 24986 30716 24998 30719
rect 26326 30716 26332 30728
rect 24986 30688 26332 30716
rect 24986 30685 24998 30688
rect 24940 30679 24998 30685
rect 26326 30676 26332 30688
rect 26384 30676 26390 30728
rect 27154 30676 27160 30728
rect 27212 30676 27218 30728
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 29733 30719 29791 30725
rect 29733 30716 29745 30719
rect 29052 30688 29745 30716
rect 29052 30676 29058 30688
rect 29733 30685 29745 30688
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 32950 30676 32956 30728
rect 33008 30716 33014 30728
rect 33229 30719 33287 30725
rect 33229 30716 33241 30719
rect 33008 30688 33241 30716
rect 33008 30676 33014 30688
rect 33229 30685 33241 30688
rect 33275 30685 33287 30719
rect 33229 30679 33287 30685
rect 33965 30719 34023 30725
rect 33965 30685 33977 30719
rect 34011 30716 34023 30719
rect 34790 30716 34796 30728
rect 34011 30688 34796 30716
rect 34011 30685 34023 30688
rect 33965 30679 34023 30685
rect 34790 30676 34796 30688
rect 34848 30716 34854 30728
rect 35434 30716 35440 30728
rect 34848 30688 35440 30716
rect 34848 30676 34854 30688
rect 35434 30676 35440 30688
rect 35492 30676 35498 30728
rect 35618 30676 35624 30728
rect 35676 30676 35682 30728
rect 40218 30676 40224 30728
rect 40276 30676 40282 30728
rect 43162 30676 43168 30728
rect 43220 30676 43226 30728
rect 36354 30608 36360 30660
rect 36412 30608 36418 30660
rect 25038 30580 25044 30592
rect 24320 30552 25044 30580
rect 25038 30540 25044 30552
rect 25096 30540 25102 30592
rect 27338 30540 27344 30592
rect 27396 30540 27402 30592
rect 27890 30540 27896 30592
rect 27948 30580 27954 30592
rect 28445 30583 28503 30589
rect 28445 30580 28457 30583
rect 27948 30552 28457 30580
rect 27948 30540 27954 30552
rect 28445 30549 28457 30552
rect 28491 30549 28503 30583
rect 28445 30543 28503 30549
rect 40586 30540 40592 30592
rect 40644 30540 40650 30592
rect 1104 30490 45172 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 45172 30490
rect 1104 30416 45172 30438
rect 2498 30336 2504 30388
rect 2556 30376 2562 30388
rect 4798 30376 4804 30388
rect 2556 30348 2774 30376
rect 2556 30336 2562 30348
rect 2746 30308 2774 30348
rect 4448 30348 4804 30376
rect 4448 30317 4476 30348
rect 4798 30336 4804 30348
rect 4856 30336 4862 30388
rect 5905 30379 5963 30385
rect 5905 30345 5917 30379
rect 5951 30345 5963 30379
rect 5905 30339 5963 30345
rect 4433 30311 4491 30317
rect 2746 30280 4200 30308
rect 4172 30249 4200 30280
rect 4433 30277 4445 30311
rect 4479 30277 4491 30311
rect 4433 30271 4491 30277
rect 4890 30268 4896 30320
rect 4948 30268 4954 30320
rect 5920 30308 5948 30339
rect 8662 30336 8668 30388
rect 8720 30376 8726 30388
rect 8720 30348 9536 30376
rect 8720 30336 8726 30348
rect 6546 30308 6552 30320
rect 5920 30280 6552 30308
rect 4157 30243 4215 30249
rect 4157 30209 4169 30243
rect 4203 30209 4215 30243
rect 5920 30240 5948 30280
rect 6546 30268 6552 30280
rect 6604 30268 6610 30320
rect 6638 30268 6644 30320
rect 6696 30308 6702 30320
rect 6696 30280 6868 30308
rect 6696 30268 6702 30280
rect 4157 30203 4215 30209
rect 5644 30212 5948 30240
rect 5534 30064 5540 30116
rect 5592 30104 5598 30116
rect 5644 30104 5672 30212
rect 6730 30200 6736 30252
rect 6788 30200 6794 30252
rect 6840 30249 6868 30280
rect 6914 30268 6920 30320
rect 6972 30268 6978 30320
rect 9508 30308 9536 30348
rect 9582 30336 9588 30388
rect 9640 30376 9646 30388
rect 12526 30376 12532 30388
rect 9640 30348 12532 30376
rect 9640 30336 9646 30348
rect 12526 30336 12532 30348
rect 12584 30336 12590 30388
rect 15838 30336 15844 30388
rect 15896 30376 15902 30388
rect 16117 30379 16175 30385
rect 16117 30376 16129 30379
rect 15896 30348 16129 30376
rect 15896 30336 15902 30348
rect 16117 30345 16129 30348
rect 16163 30345 16175 30379
rect 16117 30339 16175 30345
rect 16224 30348 16528 30376
rect 10870 30308 10876 30320
rect 9508 30280 10876 30308
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 11146 30268 11152 30320
rect 11204 30308 11210 30320
rect 12345 30311 12403 30317
rect 12345 30308 12357 30311
rect 11204 30280 12357 30308
rect 11204 30268 11210 30280
rect 12345 30277 12357 30280
rect 12391 30277 12403 30311
rect 12345 30271 12403 30277
rect 15286 30268 15292 30320
rect 15344 30308 15350 30320
rect 16224 30308 16252 30348
rect 16500 30317 16528 30348
rect 16666 30336 16672 30388
rect 16724 30376 16730 30388
rect 17678 30376 17684 30388
rect 16724 30348 17684 30376
rect 16724 30336 16730 30348
rect 16776 30317 16804 30348
rect 17678 30336 17684 30348
rect 17736 30336 17742 30388
rect 23661 30379 23719 30385
rect 23661 30345 23673 30379
rect 23707 30376 23719 30379
rect 24118 30376 24124 30388
rect 23707 30348 24124 30376
rect 23707 30345 23719 30348
rect 23661 30339 23719 30345
rect 24118 30336 24124 30348
rect 24176 30336 24182 30388
rect 32309 30379 32367 30385
rect 32309 30345 32321 30379
rect 32355 30376 32367 30379
rect 32355 30348 33264 30376
rect 32355 30345 32367 30348
rect 32309 30339 32367 30345
rect 15344 30280 16252 30308
rect 16285 30311 16343 30317
rect 15344 30268 15350 30280
rect 16285 30277 16297 30311
rect 16331 30308 16343 30311
rect 16485 30311 16543 30317
rect 16331 30277 16344 30308
rect 16285 30271 16344 30277
rect 16485 30277 16497 30311
rect 16531 30277 16543 30311
rect 16485 30271 16543 30277
rect 16761 30311 16819 30317
rect 16761 30277 16773 30311
rect 16807 30277 16819 30311
rect 16761 30271 16819 30277
rect 16945 30311 17003 30317
rect 16945 30277 16957 30311
rect 16991 30308 17003 30311
rect 18138 30308 18144 30320
rect 16991 30280 18144 30308
rect 16991 30277 17003 30280
rect 16945 30271 17003 30277
rect 6825 30243 6883 30249
rect 6825 30209 6837 30243
rect 6871 30209 6883 30243
rect 6825 30203 6883 30209
rect 7009 30243 7067 30249
rect 7009 30209 7021 30243
rect 7055 30209 7067 30243
rect 7009 30203 7067 30209
rect 5902 30132 5908 30184
rect 5960 30172 5966 30184
rect 7024 30172 7052 30203
rect 11330 30200 11336 30252
rect 11388 30240 11394 30252
rect 12621 30243 12679 30249
rect 12621 30240 12633 30243
rect 11388 30212 12633 30240
rect 11388 30200 11394 30212
rect 12621 30209 12633 30212
rect 12667 30209 12679 30243
rect 12621 30203 12679 30209
rect 16316 30184 16344 30271
rect 18138 30268 18144 30280
rect 18196 30268 18202 30320
rect 19426 30268 19432 30320
rect 19484 30308 19490 30320
rect 19521 30311 19579 30317
rect 19521 30308 19533 30311
rect 19484 30280 19533 30308
rect 19484 30268 19490 30280
rect 19521 30277 19533 30280
rect 19567 30277 19579 30311
rect 20806 30308 20812 30320
rect 20746 30280 20812 30308
rect 19521 30271 19579 30277
rect 20806 30268 20812 30280
rect 20864 30268 20870 30320
rect 22186 30268 22192 30320
rect 22244 30268 22250 30320
rect 27249 30311 27307 30317
rect 27249 30277 27261 30311
rect 27295 30308 27307 30311
rect 27338 30308 27344 30320
rect 27295 30280 27344 30308
rect 27295 30277 27307 30280
rect 27249 30271 27307 30277
rect 27338 30268 27344 30280
rect 27396 30268 27402 30320
rect 27706 30268 27712 30320
rect 27764 30268 27770 30320
rect 32493 30311 32551 30317
rect 32493 30277 32505 30311
rect 32539 30308 32551 30311
rect 32582 30308 32588 30320
rect 32539 30280 32588 30308
rect 32539 30277 32551 30280
rect 32493 30271 32551 30277
rect 32582 30268 32588 30280
rect 32640 30268 32646 30320
rect 16574 30200 16580 30252
rect 16632 30240 16638 30252
rect 16669 30243 16727 30249
rect 16669 30240 16681 30243
rect 16632 30212 16681 30240
rect 16632 30200 16638 30212
rect 16669 30209 16681 30212
rect 16715 30240 16727 30243
rect 18782 30240 18788 30252
rect 16715 30212 18788 30240
rect 16715 30209 16727 30212
rect 16669 30203 16727 30209
rect 18782 30200 18788 30212
rect 18840 30200 18846 30252
rect 24210 30200 24216 30252
rect 24268 30200 24274 30252
rect 26602 30200 26608 30252
rect 26660 30200 26666 30252
rect 29457 30243 29515 30249
rect 29457 30240 29469 30243
rect 28460 30212 29469 30240
rect 28460 30184 28488 30212
rect 29457 30209 29469 30212
rect 29503 30209 29515 30243
rect 29457 30203 29515 30209
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30240 29791 30243
rect 29914 30240 29920 30252
rect 29779 30212 29920 30240
rect 29779 30209 29791 30212
rect 29733 30203 29791 30209
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 32217 30243 32275 30249
rect 32217 30209 32229 30243
rect 32263 30209 32275 30243
rect 32217 30203 32275 30209
rect 32677 30243 32735 30249
rect 32677 30209 32689 30243
rect 32723 30240 32735 30243
rect 32989 30243 33047 30249
rect 32723 30212 32904 30240
rect 32723 30209 32735 30212
rect 32677 30203 32735 30209
rect 5960 30144 7052 30172
rect 5960 30132 5966 30144
rect 12526 30132 12532 30184
rect 12584 30132 12590 30184
rect 14090 30132 14096 30184
rect 14148 30132 14154 30184
rect 16298 30132 16304 30184
rect 16356 30172 16362 30184
rect 16356 30144 16712 30172
rect 16356 30132 16362 30144
rect 7098 30104 7104 30116
rect 5592 30076 5672 30104
rect 6288 30076 7104 30104
rect 5592 30064 5598 30076
rect 4890 29996 4896 30048
rect 4948 30036 4954 30048
rect 6288 30036 6316 30076
rect 7098 30064 7104 30076
rect 7156 30064 7162 30116
rect 12805 30107 12863 30113
rect 12805 30073 12817 30107
rect 12851 30104 12863 30107
rect 14108 30104 14136 30132
rect 16684 30113 16712 30144
rect 19150 30132 19156 30184
rect 19208 30172 19214 30184
rect 19245 30175 19303 30181
rect 19245 30172 19257 30175
rect 19208 30144 19257 30172
rect 19208 30132 19214 30144
rect 19245 30141 19257 30144
rect 19291 30141 19303 30175
rect 19245 30135 19303 30141
rect 19978 30132 19984 30184
rect 20036 30172 20042 30184
rect 20993 30175 21051 30181
rect 20993 30172 21005 30175
rect 20036 30144 21005 30172
rect 20036 30132 20042 30144
rect 20993 30141 21005 30144
rect 21039 30141 21051 30175
rect 20993 30135 21051 30141
rect 22830 30132 22836 30184
rect 22888 30132 22894 30184
rect 26142 30132 26148 30184
rect 26200 30172 26206 30184
rect 26973 30175 27031 30181
rect 26973 30172 26985 30175
rect 26200 30144 26985 30172
rect 26200 30132 26206 30144
rect 26973 30141 26985 30144
rect 27019 30141 27031 30175
rect 26973 30135 27031 30141
rect 28442 30132 28448 30184
rect 28500 30132 28506 30184
rect 28721 30175 28779 30181
rect 28721 30141 28733 30175
rect 28767 30172 28779 30175
rect 28994 30172 29000 30184
rect 28767 30144 29000 30172
rect 28767 30141 28779 30144
rect 28721 30135 28779 30141
rect 28994 30132 29000 30144
rect 29052 30132 29058 30184
rect 30282 30172 30288 30184
rect 29104 30144 30288 30172
rect 12851 30076 14136 30104
rect 16669 30107 16727 30113
rect 12851 30073 12863 30076
rect 12805 30067 12863 30073
rect 16669 30073 16681 30107
rect 16715 30073 16727 30107
rect 16669 30067 16727 30073
rect 24578 30064 24584 30116
rect 24636 30104 24642 30116
rect 24636 30076 26924 30104
rect 24636 30064 24642 30076
rect 4948 30008 6316 30036
rect 4948 29996 4954 30008
rect 6362 29996 6368 30048
rect 6420 29996 6426 30048
rect 12621 30039 12679 30045
rect 12621 30005 12633 30039
rect 12667 30036 12679 30039
rect 12710 30036 12716 30048
rect 12667 30008 12716 30036
rect 12667 30005 12679 30008
rect 12621 29999 12679 30005
rect 12710 29996 12716 30008
rect 12768 29996 12774 30048
rect 16206 29996 16212 30048
rect 16264 30036 16270 30048
rect 16301 30039 16359 30045
rect 16301 30036 16313 30039
rect 16264 30008 16313 30036
rect 16264 29996 16270 30008
rect 16301 30005 16313 30008
rect 16347 30005 16359 30039
rect 16301 29999 16359 30005
rect 26786 29996 26792 30048
rect 26844 29996 26850 30048
rect 26896 30036 26924 30076
rect 29104 30036 29132 30144
rect 30282 30132 30288 30144
rect 30340 30132 30346 30184
rect 29546 30064 29552 30116
rect 29604 30104 29610 30116
rect 29604 30076 30052 30104
rect 29604 30064 29610 30076
rect 30024 30048 30052 30076
rect 32232 30048 32260 30203
rect 32876 30172 32904 30212
rect 32989 30209 33001 30243
rect 33035 30240 33047 30243
rect 33137 30243 33195 30249
rect 33137 30240 33149 30243
rect 33035 30212 33149 30240
rect 33035 30209 33047 30212
rect 32989 30203 33047 30209
rect 33137 30209 33149 30212
rect 33183 30209 33195 30243
rect 33137 30203 33195 30209
rect 33236 30172 33264 30348
rect 33318 30336 33324 30388
rect 33376 30376 33382 30388
rect 33689 30379 33747 30385
rect 33689 30376 33701 30379
rect 33376 30348 33701 30376
rect 33376 30336 33382 30348
rect 33689 30345 33701 30348
rect 33735 30345 33747 30379
rect 33689 30339 33747 30345
rect 39482 30336 39488 30388
rect 39540 30336 39546 30388
rect 40310 30336 40316 30388
rect 40368 30376 40374 30388
rect 40681 30379 40739 30385
rect 40681 30376 40693 30379
rect 40368 30348 40693 30376
rect 40368 30336 40374 30348
rect 40681 30345 40693 30348
rect 40727 30345 40739 30379
rect 40681 30339 40739 30345
rect 33502 30268 33508 30320
rect 33560 30308 33566 30320
rect 38013 30311 38071 30317
rect 33560 30280 33732 30308
rect 33560 30268 33566 30280
rect 33318 30200 33324 30252
rect 33376 30200 33382 30252
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30209 33655 30243
rect 33597 30203 33655 30209
rect 33612 30172 33640 30203
rect 33704 30181 33732 30280
rect 38013 30277 38025 30311
rect 38059 30308 38071 30311
rect 38102 30308 38108 30320
rect 38059 30280 38108 30308
rect 38059 30277 38071 30280
rect 38013 30271 38071 30277
rect 38102 30268 38108 30280
rect 38160 30268 38166 30320
rect 39500 30308 39528 30336
rect 39669 30311 39727 30317
rect 39669 30308 39681 30311
rect 39500 30280 39681 30308
rect 39669 30277 39681 30280
rect 39715 30277 39727 30311
rect 39669 30271 39727 30277
rect 41230 30268 41236 30320
rect 41288 30268 41294 30320
rect 43530 30268 43536 30320
rect 43588 30308 43594 30320
rect 43625 30311 43683 30317
rect 43625 30308 43637 30311
rect 43588 30280 43637 30308
rect 43588 30268 43594 30280
rect 43625 30277 43637 30280
rect 43671 30277 43683 30311
rect 43625 30271 43683 30277
rect 33965 30243 34023 30249
rect 33965 30209 33977 30243
rect 34011 30240 34023 30243
rect 37277 30243 37335 30249
rect 34011 30212 34192 30240
rect 34011 30209 34023 30212
rect 33965 30203 34023 30209
rect 32876 30144 33088 30172
rect 33236 30144 33640 30172
rect 33689 30175 33747 30181
rect 32769 30107 32827 30113
rect 32769 30073 32781 30107
rect 32815 30073 32827 30107
rect 32769 30067 32827 30073
rect 32861 30107 32919 30113
rect 32861 30073 32873 30107
rect 32907 30104 32919 30107
rect 32950 30104 32956 30116
rect 32907 30076 32956 30104
rect 32907 30073 32919 30076
rect 32861 30067 32919 30073
rect 26896 30008 29132 30036
rect 29914 29996 29920 30048
rect 29972 29996 29978 30048
rect 30006 29996 30012 30048
rect 30064 29996 30070 30048
rect 32214 29996 32220 30048
rect 32272 29996 32278 30048
rect 32784 30036 32812 30067
rect 32950 30064 32956 30076
rect 33008 30064 33014 30116
rect 33060 30104 33088 30144
rect 33689 30141 33701 30175
rect 33735 30141 33747 30175
rect 33689 30135 33747 30141
rect 34164 30116 34192 30212
rect 37277 30209 37289 30243
rect 37323 30240 37335 30243
rect 37921 30243 37979 30249
rect 37323 30212 37596 30240
rect 37323 30209 37335 30212
rect 37277 30203 37335 30209
rect 34146 30104 34152 30116
rect 33060 30076 34152 30104
rect 34146 30064 34152 30076
rect 34204 30064 34210 30116
rect 37568 30113 37596 30212
rect 37921 30209 37933 30243
rect 37967 30240 37979 30243
rect 38565 30243 38623 30249
rect 38565 30240 38577 30243
rect 37967 30212 38577 30240
rect 37967 30209 37979 30212
rect 37921 30203 37979 30209
rect 38565 30209 38577 30212
rect 38611 30209 38623 30243
rect 38565 30203 38623 30209
rect 39114 30200 39120 30252
rect 39172 30240 39178 30252
rect 39301 30243 39359 30249
rect 39301 30240 39313 30243
rect 39172 30212 39313 30240
rect 39172 30200 39178 30212
rect 39301 30209 39313 30212
rect 39347 30209 39359 30243
rect 39301 30203 39359 30209
rect 39485 30243 39543 30249
rect 39485 30209 39497 30243
rect 39531 30209 39543 30243
rect 39485 30203 39543 30209
rect 38102 30132 38108 30184
rect 38160 30172 38166 30184
rect 38746 30172 38752 30184
rect 38160 30144 38752 30172
rect 38160 30132 38166 30144
rect 38746 30132 38752 30144
rect 38804 30132 38810 30184
rect 39206 30132 39212 30184
rect 39264 30172 39270 30184
rect 39500 30172 39528 30203
rect 39574 30200 39580 30252
rect 39632 30200 39638 30252
rect 39853 30243 39911 30249
rect 39853 30209 39865 30243
rect 39899 30209 39911 30243
rect 39853 30203 39911 30209
rect 39945 30243 40003 30249
rect 39945 30209 39957 30243
rect 39991 30240 40003 30243
rect 40126 30240 40132 30252
rect 39991 30212 40132 30240
rect 39991 30209 40003 30212
rect 39945 30203 40003 30209
rect 39264 30144 39528 30172
rect 39868 30172 39896 30203
rect 40126 30200 40132 30212
rect 40184 30200 40190 30252
rect 40957 30243 41015 30249
rect 40957 30209 40969 30243
rect 41003 30240 41015 30243
rect 41248 30240 41276 30268
rect 41506 30240 41512 30252
rect 41003 30212 41512 30240
rect 41003 30209 41015 30212
rect 40957 30203 41015 30209
rect 41506 30200 41512 30212
rect 41564 30200 41570 30252
rect 43162 30200 43168 30252
rect 43220 30200 43226 30252
rect 43346 30200 43352 30252
rect 43404 30200 43410 30252
rect 40034 30172 40040 30184
rect 39868 30144 40040 30172
rect 39264 30132 39270 30144
rect 40034 30132 40040 30144
rect 40092 30172 40098 30184
rect 40681 30175 40739 30181
rect 40681 30172 40693 30175
rect 40092 30144 40693 30172
rect 40092 30132 40098 30144
rect 40681 30141 40693 30144
rect 40727 30141 40739 30175
rect 43180 30172 43208 30200
rect 43441 30175 43499 30181
rect 43441 30172 43453 30175
rect 43180 30144 43453 30172
rect 40681 30135 40739 30141
rect 43441 30141 43453 30144
rect 43487 30141 43499 30175
rect 43441 30135 43499 30141
rect 37553 30107 37611 30113
rect 37553 30073 37565 30107
rect 37599 30073 37611 30107
rect 40696 30104 40724 30135
rect 41322 30104 41328 30116
rect 40696 30076 41328 30104
rect 37553 30067 37611 30073
rect 41322 30064 41328 30076
rect 41380 30064 41386 30116
rect 43070 30064 43076 30116
rect 43128 30104 43134 30116
rect 43128 30076 43392 30104
rect 43128 30064 43134 30076
rect 33134 30036 33140 30048
rect 32784 30008 33140 30036
rect 33134 29996 33140 30008
rect 33192 30036 33198 30048
rect 33873 30039 33931 30045
rect 33873 30036 33885 30039
rect 33192 30008 33885 30036
rect 33192 29996 33198 30008
rect 33873 30005 33885 30008
rect 33919 30036 33931 30039
rect 34330 30036 34336 30048
rect 33919 30008 34336 30036
rect 33919 30005 33931 30008
rect 33873 29999 33931 30005
rect 34330 29996 34336 30008
rect 34388 29996 34394 30048
rect 37458 29996 37464 30048
rect 37516 29996 37522 30048
rect 39298 29996 39304 30048
rect 39356 29996 39362 30048
rect 39666 29996 39672 30048
rect 39724 29996 39730 30048
rect 40494 29996 40500 30048
rect 40552 30036 40558 30048
rect 40865 30039 40923 30045
rect 40865 30036 40877 30039
rect 40552 30008 40877 30036
rect 40552 29996 40558 30008
rect 40865 30005 40877 30008
rect 40911 30036 40923 30039
rect 41414 30036 41420 30048
rect 40911 30008 41420 30036
rect 40911 30005 40923 30008
rect 40865 29999 40923 30005
rect 41414 29996 41420 30008
rect 41472 30036 41478 30048
rect 41966 30036 41972 30048
rect 41472 30008 41972 30036
rect 41472 29996 41478 30008
rect 41966 29996 41972 30008
rect 42024 30036 42030 30048
rect 43364 30045 43392 30076
rect 43165 30039 43223 30045
rect 43165 30036 43177 30039
rect 42024 30008 43177 30036
rect 42024 29996 42030 30008
rect 43165 30005 43177 30008
rect 43211 30005 43223 30039
rect 43165 29999 43223 30005
rect 43349 30039 43407 30045
rect 43349 30005 43361 30039
rect 43395 30005 43407 30039
rect 43349 29999 43407 30005
rect 1104 29946 45172 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 45172 29946
rect 1104 29872 45172 29894
rect 5166 29792 5172 29844
rect 5224 29792 5230 29844
rect 5353 29835 5411 29841
rect 5353 29801 5365 29835
rect 5399 29832 5411 29835
rect 6362 29832 6368 29844
rect 5399 29804 6368 29832
rect 5399 29801 5411 29804
rect 5353 29795 5411 29801
rect 6362 29792 6368 29804
rect 6420 29792 6426 29844
rect 11238 29792 11244 29844
rect 11296 29792 11302 29844
rect 12618 29792 12624 29844
rect 12676 29832 12682 29844
rect 14185 29835 14243 29841
rect 14185 29832 14197 29835
rect 12676 29804 14197 29832
rect 12676 29792 12682 29804
rect 14185 29801 14197 29804
rect 14231 29801 14243 29835
rect 14185 29795 14243 29801
rect 19334 29792 19340 29844
rect 19392 29832 19398 29844
rect 19705 29835 19763 29841
rect 19705 29832 19717 29835
rect 19392 29804 19717 29832
rect 19392 29792 19398 29804
rect 19705 29801 19717 29804
rect 19751 29801 19763 29835
rect 19705 29795 19763 29801
rect 27062 29792 27068 29844
rect 27120 29792 27126 29844
rect 27154 29792 27160 29844
rect 27212 29792 27218 29844
rect 28626 29792 28632 29844
rect 28684 29832 28690 29844
rect 28905 29835 28963 29841
rect 28905 29832 28917 29835
rect 28684 29804 28917 29832
rect 28684 29792 28690 29804
rect 28905 29801 28917 29804
rect 28951 29801 28963 29835
rect 28905 29795 28963 29801
rect 28994 29792 29000 29844
rect 29052 29792 29058 29844
rect 29362 29792 29368 29844
rect 29420 29792 29426 29844
rect 29914 29792 29920 29844
rect 29972 29792 29978 29844
rect 30190 29792 30196 29844
rect 30248 29792 30254 29844
rect 30282 29792 30288 29844
rect 30340 29832 30346 29844
rect 32306 29832 32312 29844
rect 30340 29804 32312 29832
rect 30340 29792 30346 29804
rect 32306 29792 32312 29804
rect 32364 29792 32370 29844
rect 32401 29835 32459 29841
rect 32401 29801 32413 29835
rect 32447 29832 32459 29835
rect 32447 29804 32904 29832
rect 32447 29801 32459 29804
rect 32401 29795 32459 29801
rect 6012 29736 6500 29764
rect 6012 29696 6040 29736
rect 6365 29699 6423 29705
rect 6365 29696 6377 29699
rect 5460 29668 6040 29696
rect 4982 29588 4988 29640
rect 5040 29588 5046 29640
rect 5000 29492 5028 29588
rect 5337 29563 5395 29569
rect 5337 29529 5349 29563
rect 5383 29560 5395 29563
rect 5460 29560 5488 29668
rect 5810 29628 5816 29640
rect 5552 29600 5816 29628
rect 5552 29569 5580 29600
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 5902 29588 5908 29640
rect 5960 29588 5966 29640
rect 6012 29637 6040 29668
rect 6196 29668 6377 29696
rect 6196 29640 6224 29668
rect 6365 29665 6377 29668
rect 6411 29665 6423 29699
rect 6472 29696 6500 29736
rect 27522 29724 27528 29776
rect 27580 29724 27586 29776
rect 29012 29764 29040 29792
rect 29012 29736 29224 29764
rect 6638 29696 6644 29708
rect 6472 29668 6644 29696
rect 6365 29659 6423 29665
rect 6638 29656 6644 29668
rect 6696 29656 6702 29708
rect 12250 29696 12256 29708
rect 10060 29668 12256 29696
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29597 6055 29631
rect 5997 29591 6055 29597
rect 6086 29588 6092 29640
rect 6144 29588 6150 29640
rect 6178 29588 6184 29640
rect 6236 29588 6242 29640
rect 6270 29588 6276 29640
rect 6328 29588 6334 29640
rect 10060 29637 10088 29668
rect 12250 29656 12256 29668
rect 12308 29656 12314 29708
rect 20349 29699 20407 29705
rect 15488 29668 16344 29696
rect 10045 29631 10103 29637
rect 10045 29628 10057 29631
rect 8128 29600 10057 29628
rect 5383 29532 5488 29560
rect 5537 29563 5595 29569
rect 5383 29529 5395 29532
rect 5337 29523 5395 29529
rect 5537 29529 5549 29563
rect 5583 29529 5595 29563
rect 5537 29523 5595 29529
rect 5629 29563 5687 29569
rect 5629 29529 5641 29563
rect 5675 29560 5687 29563
rect 6641 29563 6699 29569
rect 6641 29560 6653 29563
rect 5675 29532 6653 29560
rect 5675 29529 5687 29532
rect 5629 29523 5687 29529
rect 6641 29529 6653 29532
rect 6687 29529 6699 29563
rect 6641 29523 6699 29529
rect 7098 29520 7104 29572
rect 7156 29520 7162 29572
rect 8128 29501 8156 29600
rect 10045 29597 10057 29600
rect 10091 29597 10103 29631
rect 10045 29591 10103 29597
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29628 11207 29631
rect 14277 29631 14335 29637
rect 11195 29600 11468 29628
rect 11195 29597 11207 29600
rect 11149 29591 11207 29597
rect 11440 29504 11468 29600
rect 14277 29597 14289 29631
rect 14323 29628 14335 29631
rect 14918 29628 14924 29640
rect 14323 29600 14924 29628
rect 14323 29597 14335 29600
rect 14277 29591 14335 29597
rect 14918 29588 14924 29600
rect 14976 29588 14982 29640
rect 15488 29637 15516 29668
rect 16316 29640 16344 29668
rect 20349 29665 20361 29699
rect 20395 29696 20407 29699
rect 21174 29696 21180 29708
rect 20395 29668 21180 29696
rect 20395 29665 20407 29668
rect 20349 29659 20407 29665
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 27540 29696 27568 29724
rect 27709 29699 27767 29705
rect 27709 29696 27721 29699
rect 27540 29668 27721 29696
rect 27709 29665 27721 29668
rect 27755 29665 27767 29699
rect 27709 29659 27767 29665
rect 28442 29656 28448 29708
rect 28500 29696 28506 29708
rect 28997 29699 29055 29705
rect 28997 29696 29009 29699
rect 28500 29668 29009 29696
rect 28500 29656 28506 29668
rect 28997 29665 29009 29668
rect 29043 29665 29055 29699
rect 28997 29659 29055 29665
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 15212 29600 15301 29628
rect 15212 29560 15240 29600
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 15473 29631 15531 29637
rect 15473 29597 15485 29631
rect 15519 29597 15531 29631
rect 15473 29591 15531 29597
rect 15562 29588 15568 29640
rect 15620 29628 15626 29640
rect 15749 29631 15807 29637
rect 15749 29628 15761 29631
rect 15620 29600 15761 29628
rect 15620 29588 15626 29600
rect 15749 29597 15761 29600
rect 15795 29597 15807 29631
rect 15749 29591 15807 29597
rect 15657 29563 15715 29569
rect 15657 29560 15669 29563
rect 15212 29532 15669 29560
rect 15212 29504 15240 29532
rect 15657 29529 15669 29532
rect 15703 29529 15715 29563
rect 15764 29560 15792 29591
rect 16298 29588 16304 29640
rect 16356 29588 16362 29640
rect 18506 29588 18512 29640
rect 18564 29588 18570 29640
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20073 29631 20131 29637
rect 20073 29628 20085 29631
rect 20036 29600 20085 29628
rect 20036 29588 20042 29600
rect 20073 29597 20085 29600
rect 20119 29597 20131 29631
rect 20073 29591 20131 29597
rect 22281 29631 22339 29637
rect 22281 29597 22293 29631
rect 22327 29628 22339 29631
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22327 29600 22385 29628
rect 22327 29597 22339 29600
rect 22281 29591 22339 29597
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 22922 29588 22928 29640
rect 22980 29588 22986 29640
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 24949 29631 25007 29637
rect 24949 29628 24961 29631
rect 24912 29600 24961 29628
rect 24912 29588 24918 29600
rect 24949 29597 24961 29600
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 25774 29588 25780 29640
rect 25832 29628 25838 29640
rect 29196 29637 29224 29736
rect 29825 29699 29883 29705
rect 29825 29665 29837 29699
rect 29871 29696 29883 29699
rect 29932 29696 29960 29792
rect 30098 29724 30104 29776
rect 30156 29764 30162 29776
rect 31757 29767 31815 29773
rect 30156 29736 30696 29764
rect 30156 29724 30162 29736
rect 29871 29668 29960 29696
rect 29871 29665 29883 29668
rect 29825 29659 29883 29665
rect 30006 29656 30012 29708
rect 30064 29696 30070 29708
rect 30561 29699 30619 29705
rect 30561 29696 30573 29699
rect 30064 29668 30573 29696
rect 30064 29656 30070 29668
rect 30561 29665 30573 29668
rect 30607 29665 30619 29699
rect 30561 29659 30619 29665
rect 26053 29631 26111 29637
rect 26053 29628 26065 29631
rect 25832 29600 26065 29628
rect 25832 29588 25838 29600
rect 26053 29597 26065 29600
rect 26099 29628 26111 29631
rect 26421 29631 26479 29637
rect 26421 29628 26433 29631
rect 26099 29600 26433 29628
rect 26099 29597 26111 29600
rect 26053 29591 26111 29597
rect 26421 29597 26433 29600
rect 26467 29597 26479 29631
rect 26421 29591 26479 29597
rect 27525 29631 27583 29637
rect 27525 29597 27537 29631
rect 27571 29628 27583 29631
rect 29181 29631 29239 29637
rect 29181 29628 29193 29631
rect 27571 29600 29193 29628
rect 27571 29597 27583 29600
rect 27525 29591 27583 29597
rect 29181 29597 29193 29600
rect 29227 29597 29239 29631
rect 29181 29591 29239 29597
rect 29546 29588 29552 29640
rect 29604 29588 29610 29640
rect 29733 29631 29791 29637
rect 29733 29597 29745 29631
rect 29779 29628 29791 29631
rect 30377 29631 30435 29637
rect 30377 29628 30389 29631
rect 29779 29600 30389 29628
rect 29779 29597 29791 29600
rect 29733 29591 29791 29597
rect 30377 29597 30389 29600
rect 30423 29597 30435 29631
rect 30377 29591 30435 29597
rect 18524 29560 18552 29588
rect 15764 29532 18552 29560
rect 15657 29523 15715 29529
rect 24394 29520 24400 29572
rect 24452 29560 24458 29572
rect 27617 29563 27675 29569
rect 27617 29560 27629 29563
rect 24452 29532 27629 29560
rect 24452 29520 24458 29532
rect 27617 29529 27629 29532
rect 27663 29529 27675 29563
rect 27617 29523 27675 29529
rect 28626 29520 28632 29572
rect 28684 29520 28690 29572
rect 28905 29563 28963 29569
rect 28905 29529 28917 29563
rect 28951 29560 28963 29563
rect 29564 29560 29592 29588
rect 28951 29532 29592 29560
rect 28951 29529 28963 29532
rect 28905 29523 28963 29529
rect 8113 29495 8171 29501
rect 8113 29492 8125 29495
rect 5000 29464 8125 29492
rect 8113 29461 8125 29464
rect 8159 29461 8171 29495
rect 8113 29455 8171 29461
rect 10137 29495 10195 29501
rect 10137 29461 10149 29495
rect 10183 29492 10195 29495
rect 10778 29492 10784 29504
rect 10183 29464 10784 29492
rect 10183 29461 10195 29464
rect 10137 29455 10195 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11422 29452 11428 29504
rect 11480 29452 11486 29504
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 15378 29452 15384 29504
rect 15436 29452 15442 29504
rect 20165 29495 20223 29501
rect 20165 29461 20177 29495
rect 20211 29492 20223 29495
rect 21726 29492 21732 29504
rect 20211 29464 21732 29492
rect 20211 29461 20223 29464
rect 20165 29455 20223 29461
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 22094 29452 22100 29504
rect 22152 29452 22158 29504
rect 25498 29452 25504 29504
rect 25556 29452 25562 29504
rect 28644 29492 28672 29520
rect 29748 29492 29776 29591
rect 30466 29588 30472 29640
rect 30524 29588 30530 29640
rect 30668 29637 30696 29736
rect 31757 29733 31769 29767
rect 31803 29764 31815 29767
rect 32214 29764 32220 29776
rect 31803 29736 32220 29764
rect 31803 29733 31815 29736
rect 31757 29727 31815 29733
rect 32214 29724 32220 29736
rect 32272 29764 32278 29776
rect 32876 29764 32904 29804
rect 32950 29792 32956 29844
rect 33008 29792 33014 29844
rect 33318 29792 33324 29844
rect 33376 29792 33382 29844
rect 33502 29792 33508 29844
rect 33560 29792 33566 29844
rect 39298 29832 39304 29844
rect 39224 29804 39304 29832
rect 33336 29764 33364 29792
rect 32272 29736 32812 29764
rect 32272 29724 32278 29736
rect 31772 29668 32260 29696
rect 31772 29637 31800 29668
rect 32232 29637 32260 29668
rect 32784 29637 32812 29736
rect 32876 29736 33364 29764
rect 30653 29631 30711 29637
rect 30653 29597 30665 29631
rect 30699 29597 30711 29631
rect 30653 29591 30711 29597
rect 31757 29631 31815 29637
rect 31757 29597 31769 29631
rect 31803 29597 31815 29631
rect 31757 29591 31815 29597
rect 31941 29631 31999 29637
rect 31941 29597 31953 29631
rect 31987 29628 31999 29631
rect 32125 29631 32183 29637
rect 32125 29628 32137 29631
rect 31987 29600 32137 29628
rect 31987 29597 31999 29600
rect 31941 29591 31999 29597
rect 32125 29597 32137 29600
rect 32171 29597 32183 29631
rect 32125 29591 32183 29597
rect 32217 29631 32275 29637
rect 32217 29597 32229 29631
rect 32263 29597 32275 29631
rect 32217 29591 32275 29597
rect 32769 29631 32827 29637
rect 32769 29597 32781 29631
rect 32815 29597 32827 29631
rect 32769 29591 32827 29597
rect 28644 29464 29776 29492
rect 30101 29495 30159 29501
rect 30101 29461 30113 29495
rect 30147 29492 30159 29495
rect 31772 29492 31800 29591
rect 32140 29560 32168 29591
rect 32585 29563 32643 29569
rect 32140 29532 32260 29560
rect 32232 29504 32260 29532
rect 32585 29529 32597 29563
rect 32631 29560 32643 29563
rect 32876 29560 32904 29736
rect 33520 29696 33548 29792
rect 35345 29699 35403 29705
rect 33520 29668 33824 29696
rect 33594 29588 33600 29640
rect 33652 29588 33658 29640
rect 33796 29637 33824 29668
rect 35345 29665 35357 29699
rect 35391 29696 35403 29699
rect 35618 29696 35624 29708
rect 35391 29668 35624 29696
rect 35391 29665 35403 29668
rect 35345 29659 35403 29665
rect 35618 29656 35624 29668
rect 35676 29696 35682 29708
rect 35676 29668 37320 29696
rect 35676 29656 35682 29668
rect 33781 29631 33839 29637
rect 33781 29597 33793 29631
rect 33827 29597 33839 29631
rect 33781 29591 33839 29597
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 32631 29532 32904 29560
rect 33137 29563 33195 29569
rect 32631 29529 32643 29532
rect 32585 29523 32643 29529
rect 33137 29529 33149 29563
rect 33183 29560 33195 29563
rect 33183 29532 33272 29560
rect 33183 29529 33195 29532
rect 33137 29523 33195 29529
rect 33244 29504 33272 29532
rect 33318 29520 33324 29572
rect 33376 29560 33382 29572
rect 35069 29563 35127 29569
rect 35069 29560 35081 29563
rect 33376 29532 35081 29560
rect 33376 29520 33382 29532
rect 35069 29529 35081 29532
rect 35115 29529 35127 29563
rect 35069 29523 35127 29529
rect 30147 29464 31800 29492
rect 30147 29461 30159 29464
rect 30101 29455 30159 29461
rect 32214 29452 32220 29504
rect 32272 29452 32278 29504
rect 33226 29452 33232 29504
rect 33284 29452 33290 29504
rect 33781 29495 33839 29501
rect 33781 29461 33793 29495
rect 33827 29492 33839 29495
rect 34146 29492 34152 29504
rect 33827 29464 34152 29492
rect 33827 29461 33839 29464
rect 33781 29455 33839 29461
rect 34146 29452 34152 29464
rect 34204 29452 34210 29504
rect 35176 29492 35204 29591
rect 35618 29520 35624 29572
rect 35676 29520 35682 29572
rect 36354 29520 36360 29572
rect 36412 29520 36418 29572
rect 37292 29504 37320 29668
rect 39224 29637 39252 29804
rect 39298 29792 39304 29804
rect 39356 29792 39362 29844
rect 39666 29792 39672 29844
rect 39724 29792 39730 29844
rect 40126 29792 40132 29844
rect 40184 29792 40190 29844
rect 40497 29835 40555 29841
rect 40497 29801 40509 29835
rect 40543 29832 40555 29835
rect 41230 29832 41236 29844
rect 40543 29804 41236 29832
rect 40543 29801 40555 29804
rect 40497 29795 40555 29801
rect 41230 29792 41236 29804
rect 41288 29792 41294 29844
rect 41322 29792 41328 29844
rect 41380 29832 41386 29844
rect 41380 29804 42104 29832
rect 41380 29792 41386 29804
rect 39485 29699 39543 29705
rect 39485 29665 39497 29699
rect 39531 29696 39543 29699
rect 39684 29696 39712 29792
rect 41785 29767 41843 29773
rect 41785 29764 41797 29767
rect 41248 29736 41797 29764
rect 39531 29668 39712 29696
rect 39531 29665 39543 29668
rect 39485 29659 39543 29665
rect 40218 29656 40224 29708
rect 40276 29696 40282 29708
rect 40405 29699 40463 29705
rect 40405 29696 40417 29699
rect 40276 29668 40417 29696
rect 40276 29656 40282 29668
rect 40405 29665 40417 29668
rect 40451 29665 40463 29699
rect 40405 29659 40463 29665
rect 40957 29699 41015 29705
rect 40957 29665 40969 29699
rect 41003 29696 41015 29699
rect 41141 29699 41199 29705
rect 41141 29696 41153 29699
rect 41003 29668 41153 29696
rect 41003 29665 41015 29668
rect 40957 29659 41015 29665
rect 41141 29665 41153 29668
rect 41187 29665 41199 29699
rect 41141 29659 41199 29665
rect 39209 29631 39267 29637
rect 39209 29597 39221 29631
rect 39255 29597 39267 29631
rect 39209 29591 39267 29597
rect 39393 29631 39451 29637
rect 39393 29597 39405 29631
rect 39439 29628 39451 29631
rect 39850 29628 39856 29640
rect 39439 29600 39856 29628
rect 39439 29597 39451 29600
rect 39393 29591 39451 29597
rect 39850 29588 39856 29600
rect 39908 29588 39914 29640
rect 40494 29588 40500 29640
rect 40552 29588 40558 29640
rect 40770 29588 40776 29640
rect 40828 29588 40834 29640
rect 41049 29631 41107 29637
rect 41049 29597 41061 29631
rect 41095 29628 41107 29631
rect 41248 29628 41276 29736
rect 41785 29733 41797 29736
rect 41831 29733 41843 29767
rect 41785 29727 41843 29733
rect 41966 29724 41972 29776
rect 42024 29724 42030 29776
rect 42076 29764 42104 29804
rect 42978 29792 42984 29844
rect 43036 29792 43042 29844
rect 43070 29792 43076 29844
rect 43128 29832 43134 29844
rect 43625 29835 43683 29841
rect 43625 29832 43637 29835
rect 43128 29804 43637 29832
rect 43128 29792 43134 29804
rect 43625 29801 43637 29804
rect 43671 29832 43683 29835
rect 43990 29832 43996 29844
rect 43671 29804 43996 29832
rect 43671 29801 43683 29804
rect 43625 29795 43683 29801
rect 43990 29792 43996 29804
rect 44048 29792 44054 29844
rect 43530 29764 43536 29776
rect 42076 29736 43536 29764
rect 41414 29656 41420 29708
rect 41472 29656 41478 29708
rect 41506 29656 41512 29708
rect 41564 29696 41570 29708
rect 41564 29668 41828 29696
rect 41564 29656 41570 29668
rect 41095 29600 41276 29628
rect 41095 29597 41107 29600
rect 41049 29591 41107 29597
rect 41322 29588 41328 29640
rect 41380 29588 41386 29640
rect 41800 29637 41828 29668
rect 41984 29637 42012 29724
rect 42076 29637 42104 29736
rect 43530 29724 43536 29736
rect 43588 29764 43594 29776
rect 43898 29764 43904 29776
rect 43588 29736 43904 29764
rect 43588 29724 43594 29736
rect 43898 29724 43904 29736
rect 43956 29724 43962 29776
rect 43809 29699 43867 29705
rect 42923 29668 43760 29696
rect 41601 29631 41659 29637
rect 41601 29597 41613 29631
rect 41647 29597 41659 29631
rect 41601 29591 41659 29597
rect 41785 29631 41843 29637
rect 41785 29597 41797 29631
rect 41831 29628 41843 29631
rect 41969 29631 42027 29637
rect 41831 29600 41920 29628
rect 41831 29597 41843 29600
rect 41785 29591 41843 29597
rect 38933 29563 38991 29569
rect 38933 29529 38945 29563
rect 38979 29560 38991 29563
rect 39942 29560 39948 29572
rect 38979 29532 39948 29560
rect 38979 29529 38991 29532
rect 38933 29523 38991 29529
rect 39942 29520 39948 29532
rect 40000 29560 40006 29572
rect 41616 29560 41644 29591
rect 40000 29532 41092 29560
rect 41616 29532 41828 29560
rect 40000 29520 40006 29532
rect 37090 29492 37096 29504
rect 35176 29464 37096 29492
rect 37090 29452 37096 29464
rect 37148 29452 37154 29504
rect 37274 29452 37280 29504
rect 37332 29492 37338 29504
rect 37461 29495 37519 29501
rect 37461 29492 37473 29495
rect 37332 29464 37473 29492
rect 37332 29452 37338 29464
rect 37461 29461 37473 29464
rect 37507 29461 37519 29495
rect 37461 29455 37519 29461
rect 39025 29495 39083 29501
rect 39025 29461 39037 29495
rect 39071 29492 39083 29495
rect 39574 29492 39580 29504
rect 39071 29464 39580 29492
rect 39071 29461 39083 29464
rect 39025 29455 39083 29461
rect 39574 29452 39580 29464
rect 39632 29452 39638 29504
rect 40589 29495 40647 29501
rect 40589 29461 40601 29495
rect 40635 29492 40647 29495
rect 40954 29492 40960 29504
rect 40635 29464 40960 29492
rect 40635 29461 40647 29464
rect 40589 29455 40647 29461
rect 40954 29452 40960 29464
rect 41012 29452 41018 29504
rect 41064 29492 41092 29532
rect 41800 29504 41828 29532
rect 41690 29492 41696 29504
rect 41064 29464 41696 29492
rect 41690 29452 41696 29464
rect 41748 29452 41754 29504
rect 41782 29452 41788 29504
rect 41840 29452 41846 29504
rect 41892 29492 41920 29600
rect 41969 29597 41981 29631
rect 42015 29597 42027 29631
rect 41969 29591 42027 29597
rect 42061 29631 42119 29637
rect 42061 29597 42073 29631
rect 42107 29597 42119 29631
rect 42061 29591 42119 29597
rect 42702 29588 42708 29640
rect 42760 29588 42766 29640
rect 42797 29631 42855 29637
rect 42797 29597 42809 29631
rect 42843 29628 42855 29631
rect 42923 29628 42951 29668
rect 43456 29640 43484 29668
rect 42843 29600 42951 29628
rect 42843 29597 42855 29600
rect 42797 29591 42855 29597
rect 43438 29588 43444 29640
rect 43496 29588 43502 29640
rect 43533 29631 43591 29637
rect 43533 29597 43545 29631
rect 43579 29597 43591 29631
rect 43732 29628 43760 29668
rect 43809 29665 43821 29699
rect 43855 29696 43867 29699
rect 43916 29696 43944 29724
rect 44082 29696 44088 29708
rect 43855 29668 44088 29696
rect 43855 29665 43867 29668
rect 43809 29659 43867 29665
rect 44082 29656 44088 29668
rect 44140 29656 44146 29708
rect 43898 29628 43904 29640
rect 43732 29600 43904 29628
rect 43533 29591 43591 29597
rect 42886 29520 42892 29572
rect 42944 29560 42950 29572
rect 42981 29563 43039 29569
rect 42981 29560 42993 29563
rect 42944 29532 42993 29560
rect 42944 29520 42950 29532
rect 42981 29529 42993 29532
rect 43027 29529 43039 29563
rect 42981 29523 43039 29529
rect 43346 29520 43352 29572
rect 43404 29560 43410 29572
rect 43548 29560 43576 29591
rect 43898 29588 43904 29600
rect 43956 29588 43962 29640
rect 43404 29532 43576 29560
rect 43404 29520 43410 29532
rect 41966 29492 41972 29504
rect 41892 29464 41972 29492
rect 41966 29452 41972 29464
rect 42024 29452 42030 29504
rect 43806 29452 43812 29504
rect 43864 29452 43870 29504
rect 1104 29402 45172 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 45172 29402
rect 1104 29328 45172 29350
rect 5534 29248 5540 29300
rect 5592 29248 5598 29300
rect 5902 29248 5908 29300
rect 5960 29288 5966 29300
rect 5960 29260 6040 29288
rect 5960 29248 5966 29260
rect 5552 29152 5580 29248
rect 6012 29220 6040 29260
rect 6086 29248 6092 29300
rect 6144 29288 6150 29300
rect 6365 29291 6423 29297
rect 6365 29288 6377 29291
rect 6144 29260 6377 29288
rect 6144 29248 6150 29260
rect 6365 29257 6377 29260
rect 6411 29257 6423 29291
rect 6365 29251 6423 29257
rect 11330 29248 11336 29300
rect 11388 29248 11394 29300
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 12805 29291 12863 29297
rect 12805 29288 12817 29291
rect 12584 29260 12817 29288
rect 12584 29248 12590 29260
rect 12805 29257 12817 29260
rect 12851 29257 12863 29291
rect 12805 29251 12863 29257
rect 13906 29248 13912 29300
rect 13964 29288 13970 29300
rect 14553 29291 14611 29297
rect 14553 29288 14565 29291
rect 13964 29260 14565 29288
rect 13964 29248 13970 29260
rect 14553 29257 14565 29260
rect 14599 29257 14611 29291
rect 15194 29288 15200 29300
rect 14553 29251 14611 29257
rect 14752 29260 15200 29288
rect 6012 29192 10824 29220
rect 6380 29161 6408 29192
rect 10796 29164 10824 29192
rect 10870 29180 10876 29232
rect 10928 29220 10934 29232
rect 10965 29223 11023 29229
rect 10965 29220 10977 29223
rect 10928 29192 10977 29220
rect 10928 29180 10934 29192
rect 10965 29189 10977 29192
rect 11011 29189 11023 29223
rect 10965 29183 11023 29189
rect 11057 29223 11115 29229
rect 11057 29189 11069 29223
rect 11103 29220 11115 29223
rect 11793 29223 11851 29229
rect 11103 29192 11468 29220
rect 11103 29189 11115 29192
rect 11057 29183 11115 29189
rect 5721 29155 5779 29161
rect 5721 29152 5733 29155
rect 5552 29124 5733 29152
rect 5721 29121 5733 29124
rect 5767 29121 5779 29155
rect 5721 29115 5779 29121
rect 5905 29155 5963 29161
rect 5905 29121 5917 29155
rect 5951 29121 5963 29155
rect 5905 29115 5963 29121
rect 6365 29155 6423 29161
rect 6365 29121 6377 29155
rect 6411 29121 6423 29155
rect 6365 29115 6423 29121
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29152 6607 29155
rect 6638 29152 6644 29164
rect 6595 29124 6644 29152
rect 6595 29121 6607 29124
rect 6549 29115 6607 29121
rect 5920 29084 5948 29115
rect 6638 29112 6644 29124
rect 6696 29112 6702 29164
rect 6730 29112 6736 29164
rect 6788 29112 6794 29164
rect 10686 29112 10692 29164
rect 10744 29112 10750 29164
rect 10778 29112 10784 29164
rect 10836 29112 10842 29164
rect 6748 29084 6776 29112
rect 5920 29056 6776 29084
rect 10980 29084 11008 29183
rect 11440 29164 11468 29192
rect 11793 29189 11805 29223
rect 11839 29220 11851 29223
rect 12437 29223 12495 29229
rect 12437 29220 12449 29223
rect 11839 29192 12449 29220
rect 11839 29189 11851 29192
rect 11793 29183 11851 29189
rect 12437 29189 12449 29192
rect 12483 29189 12495 29223
rect 12437 29183 12495 29189
rect 12544 29192 13124 29220
rect 11238 29161 11244 29164
rect 11195 29155 11244 29161
rect 11195 29121 11207 29155
rect 11241 29121 11244 29155
rect 11195 29115 11244 29121
rect 11238 29112 11244 29115
rect 11296 29112 11302 29164
rect 11422 29112 11428 29164
rect 11480 29112 11486 29164
rect 11701 29155 11759 29161
rect 11701 29121 11713 29155
rect 11747 29121 11759 29155
rect 11701 29115 11759 29121
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29121 12219 29155
rect 12161 29115 12219 29121
rect 11716 29084 11744 29115
rect 10980 29056 11744 29084
rect 12176 29084 12204 29115
rect 12250 29112 12256 29164
rect 12308 29152 12314 29164
rect 12544 29161 12572 29192
rect 13096 29164 13124 29192
rect 12529 29155 12587 29161
rect 12308 29124 12353 29152
rect 12308 29112 12314 29124
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12667 29155 12725 29161
rect 12667 29121 12679 29155
rect 12713 29152 12725 29155
rect 12713 29124 13032 29152
rect 12713 29121 12725 29124
rect 12667 29115 12725 29121
rect 12894 29084 12900 29096
rect 12176 29056 12900 29084
rect 12894 29044 12900 29056
rect 12952 29044 12958 29096
rect 13004 29084 13032 29124
rect 13078 29112 13084 29164
rect 13136 29112 13142 29164
rect 13170 29112 13176 29164
rect 13228 29112 13234 29164
rect 14752 29161 14780 29260
rect 15194 29248 15200 29260
rect 15252 29288 15258 29300
rect 15499 29291 15557 29297
rect 15252 29260 15424 29288
rect 15252 29248 15258 29260
rect 14918 29180 14924 29232
rect 14976 29180 14982 29232
rect 15286 29180 15292 29232
rect 15344 29180 15350 29232
rect 15396 29220 15424 29260
rect 15499 29257 15511 29291
rect 15545 29288 15557 29291
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15545 29260 16037 29288
rect 15545 29257 15557 29260
rect 15499 29251 15557 29257
rect 16025 29257 16037 29260
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 16298 29248 16304 29300
rect 16356 29248 16362 29300
rect 16485 29291 16543 29297
rect 16485 29257 16497 29291
rect 16531 29288 16543 29291
rect 18417 29291 18475 29297
rect 16531 29260 16988 29288
rect 16531 29257 16543 29260
rect 16485 29251 16543 29257
rect 16316 29220 16344 29248
rect 16960 29229 16988 29260
rect 18417 29257 18429 29291
rect 18463 29288 18475 29291
rect 18506 29288 18512 29300
rect 18463 29260 18512 29288
rect 18463 29257 18475 29260
rect 18417 29251 18475 29257
rect 18506 29248 18512 29260
rect 18564 29248 18570 29300
rect 22830 29248 22836 29300
rect 22888 29288 22894 29300
rect 23201 29291 23259 29297
rect 23201 29288 23213 29291
rect 22888 29260 23213 29288
rect 22888 29248 22894 29260
rect 23201 29257 23213 29260
rect 23247 29257 23259 29291
rect 23201 29251 23259 29257
rect 24854 29248 24860 29300
rect 24912 29248 24918 29300
rect 30006 29248 30012 29300
rect 30064 29288 30070 29300
rect 30064 29260 30604 29288
rect 30064 29248 30070 29260
rect 15396 29192 16068 29220
rect 14732 29155 14790 29161
rect 14732 29121 14744 29155
rect 14778 29121 14790 29155
rect 14732 29115 14790 29121
rect 14829 29155 14887 29161
rect 14829 29121 14841 29155
rect 14875 29121 14887 29155
rect 14829 29115 14887 29121
rect 13188 29084 13216 29112
rect 13004 29056 13216 29084
rect 14844 29084 14872 29115
rect 15010 29112 15016 29164
rect 15068 29161 15074 29164
rect 15068 29155 15107 29161
rect 15095 29121 15107 29155
rect 15068 29115 15107 29121
rect 15068 29112 15074 29115
rect 15194 29112 15200 29164
rect 15252 29112 15258 29164
rect 15378 29112 15384 29164
rect 15436 29152 15442 29164
rect 16040 29161 16068 29192
rect 16224 29192 16344 29220
rect 16945 29223 17003 29229
rect 16224 29161 16252 29192
rect 16945 29189 16957 29223
rect 16991 29189 17003 29223
rect 18230 29220 18236 29232
rect 18170 29192 18236 29220
rect 16945 29183 17003 29189
rect 18230 29180 18236 29192
rect 18288 29220 18294 29232
rect 22094 29229 22100 29232
rect 22077 29223 22100 29229
rect 18288 29192 19288 29220
rect 18288 29180 18294 29192
rect 19260 29164 19288 29192
rect 22077 29189 22089 29223
rect 22077 29183 22100 29189
rect 22094 29180 22100 29183
rect 22152 29180 22158 29232
rect 24949 29223 25007 29229
rect 23492 29192 24808 29220
rect 15749 29155 15807 29161
rect 15749 29152 15761 29155
rect 15436 29124 15761 29152
rect 15436 29112 15442 29124
rect 15749 29121 15761 29124
rect 15795 29121 15807 29155
rect 15749 29115 15807 29121
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29121 16083 29155
rect 16025 29115 16083 29121
rect 16209 29155 16267 29161
rect 16209 29121 16221 29155
rect 16255 29121 16267 29155
rect 16209 29115 16267 29121
rect 16301 29155 16359 29161
rect 16301 29121 16313 29155
rect 16347 29121 16359 29155
rect 16301 29115 16359 29121
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29152 18751 29155
rect 18782 29152 18788 29164
rect 18739 29124 18788 29152
rect 18739 29121 18751 29124
rect 18693 29115 18751 29121
rect 15654 29084 15660 29096
rect 14844 29056 15660 29084
rect 15654 29044 15660 29056
rect 15712 29044 15718 29096
rect 16316 29084 16344 29115
rect 18782 29112 18788 29124
rect 18840 29112 18846 29164
rect 18877 29155 18935 29161
rect 18877 29121 18889 29155
rect 18923 29121 18935 29155
rect 18877 29115 18935 29121
rect 15948 29056 16344 29084
rect 5813 29019 5871 29025
rect 5813 28985 5825 29019
rect 5859 29016 5871 29019
rect 6638 29016 6644 29028
rect 5859 28988 6644 29016
rect 5859 28985 5871 28988
rect 5813 28979 5871 28985
rect 6638 28976 6644 28988
rect 6696 28976 6702 29028
rect 9490 29016 9496 29028
rect 7852 28988 9496 29016
rect 5994 28908 6000 28960
rect 6052 28948 6058 28960
rect 7852 28948 7880 28988
rect 9490 28976 9496 28988
rect 9548 28976 9554 29028
rect 15841 29019 15899 29025
rect 15841 29016 15853 29019
rect 15488 28988 15853 29016
rect 6052 28920 7880 28948
rect 6052 28908 6058 28920
rect 7926 28908 7932 28960
rect 7984 28948 7990 28960
rect 11054 28948 11060 28960
rect 7984 28920 11060 28948
rect 7984 28908 7990 28920
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 13262 28908 13268 28960
rect 13320 28948 13326 28960
rect 14458 28948 14464 28960
rect 13320 28920 14464 28948
rect 13320 28908 13326 28920
rect 14458 28908 14464 28920
rect 14516 28908 14522 28960
rect 15488 28957 15516 28988
rect 15841 28985 15853 28988
rect 15887 28985 15899 29019
rect 15841 28979 15899 28985
rect 15473 28951 15531 28957
rect 15473 28917 15485 28951
rect 15519 28917 15531 28951
rect 15473 28911 15531 28917
rect 15657 28951 15715 28957
rect 15657 28917 15669 28951
rect 15703 28948 15715 28951
rect 15948 28948 15976 29056
rect 16666 29044 16672 29096
rect 16724 29044 16730 29096
rect 17678 29044 17684 29096
rect 17736 29084 17742 29096
rect 18892 29084 18920 29115
rect 18966 29112 18972 29164
rect 19024 29112 19030 29164
rect 19242 29112 19248 29164
rect 19300 29112 19306 29164
rect 20625 29155 20683 29161
rect 20625 29121 20637 29155
rect 20671 29152 20683 29155
rect 21358 29152 21364 29164
rect 20671 29124 21364 29152
rect 20671 29121 20683 29124
rect 20625 29115 20683 29121
rect 21358 29112 21364 29124
rect 21416 29112 21422 29164
rect 23492 29161 23520 29192
rect 23750 29161 23756 29164
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23744 29115 23756 29161
rect 23750 29112 23756 29115
rect 23808 29112 23814 29164
rect 24780 29096 24808 29192
rect 24949 29189 24961 29223
rect 24995 29220 25007 29223
rect 25038 29220 25044 29232
rect 24995 29192 25044 29220
rect 24995 29189 25007 29192
rect 24949 29183 25007 29189
rect 25038 29180 25044 29192
rect 25096 29180 25102 29232
rect 26786 29180 26792 29232
rect 26844 29220 26850 29232
rect 27249 29223 27307 29229
rect 27249 29220 27261 29223
rect 26844 29192 27261 29220
rect 26844 29180 26850 29192
rect 27249 29189 27261 29192
rect 27295 29189 27307 29223
rect 27249 29183 27307 29189
rect 27706 29180 27712 29232
rect 27764 29180 27770 29232
rect 30466 29220 30472 29232
rect 29932 29192 30472 29220
rect 29932 29161 29960 29192
rect 30466 29180 30472 29192
rect 30524 29180 30530 29232
rect 29917 29155 29975 29161
rect 29917 29152 29929 29155
rect 28460 29124 29929 29152
rect 28460 29096 28488 29124
rect 29917 29121 29929 29124
rect 29963 29121 29975 29155
rect 29917 29115 29975 29121
rect 30098 29112 30104 29164
rect 30156 29152 30162 29164
rect 30576 29161 30604 29260
rect 32214 29248 32220 29300
rect 32272 29248 32278 29300
rect 33134 29288 33140 29300
rect 32784 29260 33140 29288
rect 32784 29229 32812 29260
rect 33134 29248 33140 29260
rect 33192 29248 33198 29300
rect 33413 29291 33471 29297
rect 33413 29257 33425 29291
rect 33459 29288 33471 29291
rect 33594 29288 33600 29300
rect 33459 29260 33600 29288
rect 33459 29257 33471 29260
rect 33413 29251 33471 29257
rect 33594 29248 33600 29260
rect 33652 29248 33658 29300
rect 35437 29291 35495 29297
rect 35437 29257 35449 29291
rect 35483 29288 35495 29291
rect 35618 29288 35624 29300
rect 35483 29260 35624 29288
rect 35483 29257 35495 29260
rect 35437 29251 35495 29257
rect 35618 29248 35624 29260
rect 35676 29248 35682 29300
rect 37090 29248 37096 29300
rect 37148 29248 37154 29300
rect 39025 29291 39083 29297
rect 39025 29257 39037 29291
rect 39071 29288 39083 29291
rect 39206 29288 39212 29300
rect 39071 29260 39212 29288
rect 39071 29257 39083 29260
rect 39025 29251 39083 29257
rect 32769 29223 32827 29229
rect 32769 29189 32781 29223
rect 32815 29189 32827 29223
rect 32769 29183 32827 29189
rect 32953 29223 33011 29229
rect 32953 29189 32965 29223
rect 32999 29220 33011 29223
rect 34146 29220 34152 29232
rect 32999 29192 34152 29220
rect 32999 29189 33011 29192
rect 32953 29183 33011 29189
rect 34146 29180 34152 29192
rect 34204 29180 34210 29232
rect 35069 29223 35127 29229
rect 35069 29220 35081 29223
rect 34256 29192 35081 29220
rect 30377 29155 30435 29161
rect 30377 29152 30389 29155
rect 30156 29124 30389 29152
rect 30156 29112 30162 29124
rect 30377 29121 30389 29124
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 30561 29155 30619 29161
rect 30561 29121 30573 29155
rect 30607 29121 30619 29155
rect 30561 29115 30619 29121
rect 32309 29155 32367 29161
rect 32309 29121 32321 29155
rect 32355 29152 32367 29155
rect 32674 29152 32680 29164
rect 32355 29124 32680 29152
rect 32355 29121 32367 29124
rect 32309 29115 32367 29121
rect 32674 29112 32680 29124
rect 32732 29112 32738 29164
rect 33226 29112 33232 29164
rect 33284 29112 33290 29164
rect 33318 29112 33324 29164
rect 33376 29152 33382 29164
rect 33413 29155 33471 29161
rect 33413 29152 33425 29155
rect 33376 29124 33425 29152
rect 33376 29112 33382 29124
rect 33413 29121 33425 29124
rect 33459 29121 33471 29155
rect 33413 29115 33471 29121
rect 33502 29112 33508 29164
rect 33560 29152 33566 29164
rect 34256 29152 34284 29192
rect 35069 29189 35081 29192
rect 35115 29189 35127 29223
rect 35069 29183 35127 29189
rect 35161 29223 35219 29229
rect 35161 29189 35173 29223
rect 35207 29220 35219 29223
rect 35529 29223 35587 29229
rect 35529 29220 35541 29223
rect 35207 29192 35541 29220
rect 35207 29189 35219 29192
rect 35161 29183 35219 29189
rect 35529 29189 35541 29192
rect 35575 29189 35587 29223
rect 35529 29183 35587 29189
rect 33560 29124 34284 29152
rect 33560 29112 33566 29124
rect 34790 29112 34796 29164
rect 34848 29152 34854 29164
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34848 29124 34897 29152
rect 34848 29112 34854 29124
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 35253 29155 35311 29161
rect 35253 29121 35265 29155
rect 35299 29121 35311 29155
rect 35253 29115 35311 29121
rect 36173 29155 36231 29161
rect 36173 29121 36185 29155
rect 36219 29152 36231 29155
rect 37108 29152 37136 29248
rect 37458 29180 37464 29232
rect 37516 29220 37522 29232
rect 37553 29223 37611 29229
rect 37553 29220 37565 29223
rect 37516 29192 37565 29220
rect 37516 29180 37522 29192
rect 37553 29189 37565 29192
rect 37599 29189 37611 29223
rect 37553 29183 37611 29189
rect 39022 29152 39028 29164
rect 36219 29124 37136 29152
rect 38686 29124 39028 29152
rect 36219 29121 36231 29124
rect 36173 29115 36231 29121
rect 17736 29056 18957 29084
rect 17736 29044 17742 29056
rect 15703 28920 15976 28948
rect 15703 28917 15715 28920
rect 15657 28911 15715 28917
rect 18506 28908 18512 28960
rect 18564 28908 18570 28960
rect 18892 28948 18920 29056
rect 21542 29044 21548 29096
rect 21600 29084 21606 29096
rect 21821 29087 21879 29093
rect 21821 29084 21833 29087
rect 21600 29056 21833 29084
rect 21600 29044 21606 29056
rect 21821 29053 21833 29056
rect 21867 29053 21879 29087
rect 21821 29047 21879 29053
rect 24762 29044 24768 29096
rect 24820 29044 24826 29096
rect 26973 29087 27031 29093
rect 26973 29053 26985 29087
rect 27019 29053 27031 29087
rect 26973 29047 27031 29053
rect 19153 29019 19211 29025
rect 19153 28985 19165 29019
rect 19199 29016 19211 29019
rect 19426 29016 19432 29028
rect 19199 28988 19432 29016
rect 19199 28985 19211 28988
rect 19153 28979 19211 28985
rect 19426 28976 19432 28988
rect 19484 28976 19490 29028
rect 24780 29016 24808 29044
rect 26142 29016 26148 29028
rect 20180 28988 20576 29016
rect 24780 28988 26148 29016
rect 20180 28948 20208 28988
rect 18892 28920 20208 28948
rect 20254 28908 20260 28960
rect 20312 28948 20318 28960
rect 20441 28951 20499 28957
rect 20441 28948 20453 28951
rect 20312 28920 20453 28948
rect 20312 28908 20318 28920
rect 20441 28917 20453 28920
rect 20487 28917 20499 28951
rect 20548 28948 20576 28988
rect 26142 28976 26148 28988
rect 26200 29016 26206 29028
rect 26237 29019 26295 29025
rect 26237 29016 26249 29019
rect 26200 28988 26249 29016
rect 26200 28976 26206 28988
rect 26237 28985 26249 28988
rect 26283 29016 26295 29019
rect 26988 29016 27016 29047
rect 28442 29044 28448 29096
rect 28500 29044 28506 29096
rect 30009 29087 30067 29093
rect 30009 29053 30021 29087
rect 30055 29084 30067 29087
rect 30469 29087 30527 29093
rect 30469 29084 30481 29087
rect 30055 29056 30481 29084
rect 30055 29053 30067 29056
rect 30009 29047 30067 29053
rect 30469 29053 30481 29056
rect 30515 29053 30527 29087
rect 33244 29084 33272 29112
rect 30469 29047 30527 29053
rect 31726 29056 33272 29084
rect 28721 29019 28779 29025
rect 28721 29016 28733 29019
rect 26283 28988 27016 29016
rect 28644 28988 28733 29016
rect 26283 28985 26295 28988
rect 26237 28979 26295 28985
rect 28644 28960 28672 28988
rect 28721 28985 28733 28988
rect 28767 28985 28779 29019
rect 28721 28979 28779 28985
rect 30285 29019 30343 29025
rect 30285 28985 30297 29019
rect 30331 29016 30343 29019
rect 31726 29016 31754 29056
rect 34054 29044 34060 29096
rect 34112 29084 34118 29096
rect 35268 29084 35296 29115
rect 39022 29112 39028 29124
rect 39080 29112 39086 29164
rect 39132 29161 39160 29260
rect 39206 29248 39212 29260
rect 39264 29248 39270 29300
rect 39301 29291 39359 29297
rect 39301 29257 39313 29291
rect 39347 29288 39359 29291
rect 39390 29288 39396 29300
rect 39347 29260 39396 29288
rect 39347 29257 39359 29260
rect 39301 29251 39359 29257
rect 39390 29248 39396 29260
rect 39448 29248 39454 29300
rect 39850 29248 39856 29300
rect 39908 29248 39914 29300
rect 40126 29248 40132 29300
rect 40184 29248 40190 29300
rect 40218 29248 40224 29300
rect 40276 29248 40282 29300
rect 40770 29297 40776 29300
rect 40766 29288 40776 29297
rect 40731 29260 40776 29288
rect 40766 29251 40776 29260
rect 40770 29248 40776 29251
rect 40828 29248 40834 29300
rect 41049 29291 41107 29297
rect 41049 29257 41061 29291
rect 41095 29288 41107 29291
rect 41782 29288 41788 29300
rect 41095 29260 41788 29288
rect 41095 29257 41107 29260
rect 41049 29251 41107 29257
rect 39942 29220 39948 29232
rect 39224 29192 39948 29220
rect 39117 29155 39175 29161
rect 39117 29121 39129 29155
rect 39163 29121 39175 29155
rect 39117 29115 39175 29121
rect 34112 29056 35296 29084
rect 34112 29044 34118 29056
rect 37274 29044 37280 29096
rect 37332 29044 37338 29096
rect 38746 29084 38752 29096
rect 37384 29056 38752 29084
rect 30331 28988 31754 29016
rect 30331 28985 30343 28988
rect 30285 28979 30343 28985
rect 32306 28976 32312 29028
rect 32364 29016 32370 29028
rect 37384 29016 37412 29056
rect 38746 29044 38752 29056
rect 38804 29084 38810 29096
rect 39224 29084 39252 29192
rect 39942 29180 39948 29192
rect 40000 29180 40006 29232
rect 39482 29112 39488 29164
rect 39540 29112 39546 29164
rect 39761 29155 39819 29161
rect 39761 29121 39773 29155
rect 39807 29152 39819 29155
rect 40037 29155 40095 29161
rect 40037 29152 40049 29155
rect 39807 29124 40049 29152
rect 39807 29121 39819 29124
rect 39761 29115 39819 29121
rect 40037 29121 40049 29124
rect 40083 29152 40095 29155
rect 40144 29152 40172 29248
rect 40236 29220 40264 29248
rect 40681 29223 40739 29229
rect 40681 29220 40693 29223
rect 40236 29192 40693 29220
rect 40681 29189 40693 29192
rect 40727 29189 40739 29223
rect 40681 29183 40739 29189
rect 40083 29124 40172 29152
rect 40083 29121 40095 29124
rect 40037 29115 40095 29121
rect 40402 29112 40408 29164
rect 40460 29152 40466 29164
rect 40589 29155 40647 29161
rect 40589 29152 40601 29155
rect 40460 29124 40601 29152
rect 40460 29112 40466 29124
rect 40589 29121 40601 29124
rect 40635 29121 40647 29155
rect 40589 29115 40647 29121
rect 40862 29112 40868 29164
rect 40920 29112 40926 29164
rect 38804 29056 39252 29084
rect 38804 29044 38810 29056
rect 32364 28988 37412 29016
rect 39500 29016 39528 29112
rect 39942 29044 39948 29096
rect 40000 29084 40006 29096
rect 40129 29087 40187 29093
rect 40129 29084 40141 29087
rect 40000 29056 40141 29084
rect 40000 29044 40006 29056
rect 40129 29053 40141 29056
rect 40175 29053 40187 29087
rect 40129 29047 40187 29053
rect 40221 29087 40279 29093
rect 40221 29053 40233 29087
rect 40267 29053 40279 29087
rect 40221 29047 40279 29053
rect 40313 29087 40371 29093
rect 40313 29053 40325 29087
rect 40359 29084 40371 29087
rect 41064 29084 41092 29251
rect 41782 29248 41788 29260
rect 41840 29248 41846 29300
rect 42978 29248 42984 29300
rect 43036 29288 43042 29300
rect 43254 29288 43260 29300
rect 43036 29260 43260 29288
rect 43036 29248 43042 29260
rect 43254 29248 43260 29260
rect 43312 29248 43318 29300
rect 43346 29248 43352 29300
rect 43404 29248 43410 29300
rect 43806 29248 43812 29300
rect 43864 29248 43870 29300
rect 43898 29248 43904 29300
rect 43956 29248 43962 29300
rect 41417 29223 41475 29229
rect 41417 29189 41429 29223
rect 41463 29220 41475 29223
rect 41506 29220 41512 29232
rect 41463 29192 41512 29220
rect 41463 29189 41475 29192
rect 41417 29183 41475 29189
rect 41506 29180 41512 29192
rect 41564 29180 41570 29232
rect 41708 29192 42196 29220
rect 41141 29155 41199 29161
rect 41141 29121 41153 29155
rect 41187 29152 41199 29155
rect 41322 29152 41328 29164
rect 41187 29124 41328 29152
rect 41187 29121 41199 29124
rect 41141 29115 41199 29121
rect 41322 29112 41328 29124
rect 41380 29152 41386 29164
rect 41708 29161 41736 29192
rect 42168 29164 42196 29192
rect 42702 29180 42708 29232
rect 42760 29220 42766 29232
rect 43364 29220 43392 29248
rect 42760 29192 43116 29220
rect 43364 29192 43484 29220
rect 42760 29180 42766 29192
rect 41693 29155 41751 29161
rect 41380 29124 41644 29152
rect 41380 29112 41386 29124
rect 40359 29056 41092 29084
rect 40359 29053 40371 29056
rect 40313 29047 40371 29053
rect 40034 29016 40040 29028
rect 39500 28988 40040 29016
rect 32364 28976 32370 28988
rect 40034 28976 40040 28988
rect 40092 29016 40098 29028
rect 40236 29016 40264 29047
rect 40092 28988 40264 29016
rect 40092 28976 40098 28988
rect 21266 28948 21272 28960
rect 20548 28920 21272 28948
rect 20441 28911 20499 28917
rect 21266 28908 21272 28920
rect 21324 28908 21330 28960
rect 28626 28908 28632 28960
rect 28684 28908 28690 28960
rect 33134 28908 33140 28960
rect 33192 28908 33198 28960
rect 39577 28951 39635 28957
rect 39577 28917 39589 28951
rect 39623 28948 39635 28951
rect 40328 28948 40356 29047
rect 41230 29044 41236 29096
rect 41288 29044 41294 29096
rect 41616 29093 41644 29124
rect 41693 29121 41705 29155
rect 41739 29121 41751 29155
rect 41693 29115 41751 29121
rect 41966 29112 41972 29164
rect 42024 29152 42030 29164
rect 42061 29155 42119 29161
rect 42061 29152 42073 29155
rect 42024 29124 42073 29152
rect 42024 29112 42030 29124
rect 42061 29121 42073 29124
rect 42107 29121 42119 29155
rect 42061 29115 42119 29121
rect 42150 29112 42156 29164
rect 42208 29112 42214 29164
rect 42242 29112 42248 29164
rect 42300 29112 42306 29164
rect 42797 29155 42855 29161
rect 42797 29152 42809 29155
rect 42444 29124 42809 29152
rect 41601 29087 41659 29093
rect 41601 29053 41613 29087
rect 41647 29084 41659 29087
rect 42444 29084 42472 29124
rect 42797 29121 42809 29124
rect 42843 29121 42855 29155
rect 42797 29115 42855 29121
rect 42886 29112 42892 29164
rect 42944 29112 42950 29164
rect 42981 29155 43039 29161
rect 42981 29121 42993 29155
rect 43027 29121 43039 29155
rect 42981 29115 43039 29121
rect 41647 29056 42472 29084
rect 42521 29087 42579 29093
rect 41647 29053 41659 29056
rect 41601 29047 41659 29053
rect 42521 29053 42533 29087
rect 42567 29084 42579 29087
rect 42904 29084 42932 29112
rect 42567 29056 42932 29084
rect 42567 29053 42579 29056
rect 42521 29047 42579 29053
rect 40862 28976 40868 29028
rect 40920 28976 40926 29028
rect 42536 29016 42564 29047
rect 42260 28988 42564 29016
rect 39623 28920 40356 28948
rect 40880 28948 40908 28976
rect 41230 28948 41236 28960
rect 40880 28920 41236 28948
rect 39623 28917 39635 28920
rect 39577 28911 39635 28917
rect 41230 28908 41236 28920
rect 41288 28948 41294 28960
rect 42260 28948 42288 28988
rect 42610 28976 42616 29028
rect 42668 28976 42674 29028
rect 42996 29016 43024 29115
rect 43088 29084 43116 29192
rect 43162 29112 43168 29164
rect 43220 29152 43226 29164
rect 43349 29155 43407 29161
rect 43349 29152 43361 29155
rect 43220 29124 43361 29152
rect 43220 29112 43226 29124
rect 43349 29121 43361 29124
rect 43395 29121 43407 29155
rect 43456 29152 43484 29192
rect 43456 29124 43576 29152
rect 43349 29115 43407 29121
rect 43257 29087 43315 29093
rect 43257 29084 43269 29087
rect 43088 29056 43269 29084
rect 43257 29053 43269 29056
rect 43303 29084 43315 29087
rect 43438 29084 43444 29096
rect 43303 29056 43444 29084
rect 43303 29053 43315 29056
rect 43257 29047 43315 29053
rect 43438 29044 43444 29056
rect 43496 29044 43502 29096
rect 43548 29084 43576 29124
rect 43714 29112 43720 29164
rect 43772 29112 43778 29164
rect 43824 29152 43852 29248
rect 43916 29220 43944 29248
rect 43916 29192 44680 29220
rect 44652 29161 44680 29192
rect 44637 29155 44695 29161
rect 43824 29124 44588 29152
rect 43806 29084 43812 29096
rect 43548 29056 43812 29084
rect 43806 29044 43812 29056
rect 43864 29044 43870 29096
rect 43898 29044 43904 29096
rect 43956 29044 43962 29096
rect 43993 29087 44051 29093
rect 43993 29053 44005 29087
rect 44039 29084 44051 29087
rect 44082 29084 44088 29096
rect 44039 29056 44088 29084
rect 44039 29053 44051 29056
rect 43993 29047 44051 29053
rect 44082 29044 44088 29056
rect 44140 29044 44146 29096
rect 44560 29093 44588 29124
rect 44637 29121 44649 29155
rect 44683 29121 44695 29155
rect 44637 29115 44695 29121
rect 44545 29087 44603 29093
rect 44545 29053 44557 29087
rect 44591 29053 44603 29087
rect 44545 29047 44603 29053
rect 44269 29019 44327 29025
rect 44269 29016 44281 29019
rect 42996 28988 44281 29016
rect 44269 28985 44281 28988
rect 44315 28985 44327 29019
rect 44269 28979 44327 28985
rect 41288 28920 42288 28948
rect 41288 28908 41294 28920
rect 43898 28908 43904 28960
rect 43956 28948 43962 28960
rect 44177 28951 44235 28957
rect 44177 28948 44189 28951
rect 43956 28920 44189 28948
rect 43956 28908 43962 28920
rect 44177 28917 44189 28920
rect 44223 28917 44235 28951
rect 44177 28911 44235 28917
rect 1104 28858 45172 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 45172 28858
rect 1104 28784 45172 28806
rect 6549 28747 6607 28753
rect 6549 28713 6561 28747
rect 6595 28744 6607 28747
rect 6730 28744 6736 28756
rect 6595 28716 6736 28744
rect 6595 28713 6607 28716
rect 6549 28707 6607 28713
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 7926 28704 7932 28756
rect 7984 28744 7990 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 7984 28716 8493 28744
rect 7984 28704 7990 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 8481 28707 8539 28713
rect 8588 28716 8984 28744
rect 8294 28676 8300 28688
rect 6196 28648 8300 28676
rect 5258 28568 5264 28620
rect 5316 28608 5322 28620
rect 5994 28608 6000 28620
rect 5316 28580 6000 28608
rect 5316 28568 5322 28580
rect 5994 28568 6000 28580
rect 6052 28568 6058 28620
rect 6196 28608 6224 28648
rect 8294 28636 8300 28648
rect 8352 28636 8358 28688
rect 8205 28611 8263 28617
rect 8205 28608 8217 28611
rect 6104 28580 6224 28608
rect 7852 28580 8217 28608
rect 6104 28549 6132 28580
rect 5445 28543 5503 28549
rect 5445 28509 5457 28543
rect 5491 28540 5503 28543
rect 6089 28543 6147 28549
rect 6089 28540 6101 28543
rect 5491 28512 6101 28540
rect 5491 28509 5503 28512
rect 5445 28503 5503 28509
rect 6089 28509 6101 28512
rect 6135 28509 6147 28543
rect 6089 28503 6147 28509
rect 6181 28543 6239 28549
rect 6181 28509 6193 28543
rect 6227 28509 6239 28543
rect 6181 28503 6239 28509
rect 5721 28475 5779 28481
rect 5721 28472 5733 28475
rect 5460 28444 5733 28472
rect 5460 28416 5488 28444
rect 5721 28441 5733 28444
rect 5767 28441 5779 28475
rect 5721 28435 5779 28441
rect 5810 28432 5816 28484
rect 5868 28432 5874 28484
rect 5905 28475 5963 28481
rect 5905 28441 5917 28475
rect 5951 28472 5963 28475
rect 5994 28472 6000 28484
rect 5951 28444 6000 28472
rect 5951 28441 5963 28444
rect 5905 28435 5963 28441
rect 5994 28432 6000 28444
rect 6052 28432 6058 28484
rect 5442 28364 5448 28416
rect 5500 28364 5506 28416
rect 5626 28364 5632 28416
rect 5684 28364 5690 28416
rect 5828 28404 5856 28432
rect 6196 28404 6224 28503
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 6733 28543 6791 28549
rect 6733 28509 6745 28543
rect 6779 28540 6791 28543
rect 6822 28540 6828 28552
rect 6779 28512 6828 28540
rect 6779 28509 6791 28512
rect 6733 28503 6791 28509
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 5828 28376 6224 28404
rect 6362 28364 6368 28416
rect 6420 28404 6426 28416
rect 7852 28404 7880 28580
rect 8205 28577 8217 28580
rect 8251 28608 8263 28611
rect 8588 28608 8616 28716
rect 8956 28676 8984 28716
rect 9122 28704 9128 28756
rect 9180 28704 9186 28756
rect 10505 28747 10563 28753
rect 10505 28713 10517 28747
rect 10551 28744 10563 28747
rect 10686 28744 10692 28756
rect 10551 28716 10692 28744
rect 10551 28713 10563 28716
rect 10505 28707 10563 28713
rect 10686 28704 10692 28716
rect 10744 28704 10750 28756
rect 11238 28704 11244 28756
rect 11296 28704 11302 28756
rect 12894 28704 12900 28756
rect 12952 28704 12958 28756
rect 13538 28704 13544 28756
rect 13596 28744 13602 28756
rect 13725 28747 13783 28753
rect 13725 28744 13737 28747
rect 13596 28716 13737 28744
rect 13596 28704 13602 28716
rect 13725 28713 13737 28716
rect 13771 28713 13783 28747
rect 13725 28707 13783 28713
rect 15194 28704 15200 28756
rect 15252 28744 15258 28756
rect 15289 28747 15347 28753
rect 15289 28744 15301 28747
rect 15252 28716 15301 28744
rect 15252 28704 15258 28716
rect 15289 28713 15301 28716
rect 15335 28713 15347 28747
rect 18141 28747 18199 28753
rect 15289 28707 15347 28713
rect 17604 28716 18000 28744
rect 12710 28676 12716 28688
rect 8956 28648 12716 28676
rect 12710 28636 12716 28648
rect 12768 28676 12774 28688
rect 13262 28676 13268 28688
rect 12768 28648 13268 28676
rect 12768 28636 12774 28648
rect 13262 28636 13268 28648
rect 13320 28636 13326 28688
rect 13814 28636 13820 28688
rect 13872 28636 13878 28688
rect 8251 28580 8616 28608
rect 8251 28577 8263 28580
rect 8205 28571 8263 28577
rect 8662 28568 8668 28620
rect 8720 28608 8726 28620
rect 9214 28608 9220 28620
rect 8720 28580 9220 28608
rect 8720 28568 8726 28580
rect 9214 28568 9220 28580
rect 9272 28568 9278 28620
rect 9490 28568 9496 28620
rect 9548 28608 9554 28620
rect 10045 28611 10103 28617
rect 10045 28608 10057 28611
rect 9548 28580 10057 28608
rect 9548 28568 9554 28580
rect 10045 28577 10057 28580
rect 10091 28577 10103 28611
rect 10045 28571 10103 28577
rect 11054 28568 11060 28620
rect 11112 28608 11118 28620
rect 11112 28580 11192 28608
rect 11112 28568 11118 28580
rect 7926 28500 7932 28552
rect 7984 28500 7990 28552
rect 8021 28543 8079 28549
rect 8021 28509 8033 28543
rect 8067 28540 8079 28543
rect 8478 28540 8484 28552
rect 8067 28512 8484 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 8478 28500 8484 28512
rect 8536 28540 8542 28552
rect 9401 28543 9459 28549
rect 9401 28540 9413 28543
rect 8536 28512 9413 28540
rect 8536 28500 8542 28512
rect 9401 28509 9413 28512
rect 9447 28509 9459 28543
rect 9401 28503 9459 28509
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28540 10195 28543
rect 10594 28540 10600 28552
rect 10183 28512 10600 28540
rect 10183 28509 10195 28512
rect 10137 28503 10195 28509
rect 10594 28500 10600 28512
rect 10652 28500 10658 28552
rect 11164 28549 11192 28580
rect 13446 28568 13452 28620
rect 13504 28608 13510 28620
rect 13832 28608 13860 28636
rect 13504 28580 13860 28608
rect 15749 28611 15807 28617
rect 13504 28568 13510 28580
rect 15749 28577 15761 28611
rect 15795 28608 15807 28611
rect 16022 28608 16028 28620
rect 15795 28580 16028 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 16022 28568 16028 28580
rect 16080 28608 16086 28620
rect 16390 28608 16396 28620
rect 16080 28580 16396 28608
rect 16080 28568 16086 28580
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28509 11207 28543
rect 11149 28503 11207 28509
rect 13078 28500 13084 28552
rect 13136 28500 13142 28552
rect 13170 28500 13176 28552
rect 13228 28500 13234 28552
rect 13817 28543 13875 28549
rect 13817 28509 13829 28543
rect 13863 28509 13875 28543
rect 13817 28503 13875 28509
rect 8205 28475 8263 28481
rect 8205 28441 8217 28475
rect 8251 28472 8263 28475
rect 8570 28472 8576 28484
rect 8251 28444 8576 28472
rect 8251 28441 8263 28444
rect 8205 28435 8263 28441
rect 8570 28432 8576 28444
rect 8628 28432 8634 28484
rect 8662 28432 8668 28484
rect 8720 28432 8726 28484
rect 8938 28432 8944 28484
rect 8996 28432 9002 28484
rect 9157 28475 9215 28481
rect 9157 28441 9169 28475
rect 9203 28472 9215 28475
rect 9493 28475 9551 28481
rect 9493 28472 9505 28475
rect 9203 28444 9505 28472
rect 9203 28441 9215 28444
rect 9157 28435 9215 28441
rect 9493 28441 9505 28444
rect 9539 28441 9551 28475
rect 9493 28435 9551 28441
rect 13538 28432 13544 28484
rect 13596 28432 13602 28484
rect 13832 28416 13860 28503
rect 14458 28500 14464 28552
rect 14516 28500 14522 28552
rect 15657 28543 15715 28549
rect 15657 28509 15669 28543
rect 15703 28540 15715 28543
rect 15930 28540 15936 28552
rect 15703 28512 15936 28540
rect 15703 28509 15715 28512
rect 15657 28503 15715 28509
rect 15930 28500 15936 28512
rect 15988 28540 15994 28552
rect 17126 28540 17132 28552
rect 15988 28512 17132 28540
rect 15988 28500 15994 28512
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 17604 28549 17632 28716
rect 17972 28608 18000 28716
rect 18141 28713 18153 28747
rect 18187 28744 18199 28747
rect 18506 28744 18512 28756
rect 18187 28716 18512 28744
rect 18187 28713 18199 28716
rect 18141 28707 18199 28713
rect 18506 28704 18512 28716
rect 18564 28704 18570 28756
rect 18966 28704 18972 28756
rect 19024 28704 19030 28756
rect 21358 28704 21364 28756
rect 21416 28704 21422 28756
rect 21450 28704 21456 28756
rect 21508 28704 21514 28756
rect 22465 28747 22523 28753
rect 22465 28713 22477 28747
rect 22511 28744 22523 28747
rect 22922 28744 22928 28756
rect 22511 28716 22928 28744
rect 22511 28713 22523 28716
rect 22465 28707 22523 28713
rect 22922 28704 22928 28716
rect 22980 28704 22986 28756
rect 26329 28747 26387 28753
rect 26329 28713 26341 28747
rect 26375 28744 26387 28747
rect 26418 28744 26424 28756
rect 26375 28716 26424 28744
rect 26375 28713 26387 28716
rect 26329 28707 26387 28713
rect 26418 28704 26424 28716
rect 26476 28704 26482 28756
rect 26602 28704 26608 28756
rect 26660 28744 26666 28756
rect 26697 28747 26755 28753
rect 26697 28744 26709 28747
rect 26660 28716 26709 28744
rect 26660 28704 26666 28716
rect 26697 28713 26709 28716
rect 26743 28713 26755 28747
rect 26697 28707 26755 28713
rect 34790 28704 34796 28756
rect 34848 28744 34854 28756
rect 35069 28747 35127 28753
rect 35069 28744 35081 28747
rect 34848 28716 35081 28744
rect 34848 28704 34854 28716
rect 35069 28713 35081 28716
rect 35115 28713 35127 28747
rect 35069 28707 35127 28713
rect 40420 28716 41414 28744
rect 18325 28679 18383 28685
rect 18325 28645 18337 28679
rect 18371 28676 18383 28679
rect 18984 28676 19012 28704
rect 21468 28676 21496 28704
rect 40420 28688 40448 28716
rect 18371 28648 19012 28676
rect 20548 28648 21496 28676
rect 18371 28645 18383 28648
rect 18325 28639 18383 28645
rect 18417 28611 18475 28617
rect 18417 28608 18429 28611
rect 17972 28580 18429 28608
rect 18417 28577 18429 28580
rect 18463 28577 18475 28611
rect 19058 28608 19064 28620
rect 18417 28571 18475 28577
rect 18984 28580 19064 28608
rect 17405 28543 17463 28549
rect 17405 28509 17417 28543
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28509 17647 28543
rect 17589 28503 17647 28509
rect 14476 28472 14504 28500
rect 17420 28472 17448 28503
rect 17678 28500 17684 28552
rect 17736 28500 17742 28552
rect 17865 28543 17923 28549
rect 17865 28509 17877 28543
rect 17911 28540 17923 28543
rect 18782 28540 18788 28552
rect 17911 28512 18788 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 18782 28500 18788 28512
rect 18840 28540 18846 28552
rect 18984 28549 19012 28580
rect 19058 28568 19064 28580
rect 19116 28608 19122 28620
rect 20548 28608 20576 28648
rect 24210 28636 24216 28688
rect 24268 28636 24274 28688
rect 33410 28636 33416 28688
rect 33468 28676 33474 28688
rect 33870 28676 33876 28688
rect 33468 28648 33876 28676
rect 33468 28636 33474 28648
rect 33870 28636 33876 28648
rect 33928 28676 33934 28688
rect 35618 28676 35624 28688
rect 33928 28648 35624 28676
rect 33928 28636 33934 28648
rect 35618 28636 35624 28648
rect 35676 28636 35682 28688
rect 39114 28636 39120 28688
rect 39172 28676 39178 28688
rect 39393 28679 39451 28685
rect 39393 28676 39405 28679
rect 39172 28648 39405 28676
rect 39172 28636 39178 28648
rect 39393 28645 39405 28648
rect 39439 28645 39451 28679
rect 40402 28676 40408 28688
rect 39393 28639 39451 28645
rect 39776 28648 40408 28676
rect 19116 28580 20576 28608
rect 19116 28568 19122 28580
rect 21266 28568 21272 28620
rect 21324 28568 21330 28620
rect 22002 28568 22008 28620
rect 22060 28608 22066 28620
rect 23109 28611 23167 28617
rect 23109 28608 23121 28611
rect 22060 28580 23121 28608
rect 22060 28568 22066 28580
rect 23109 28577 23121 28580
rect 23155 28608 23167 28611
rect 23290 28608 23296 28620
rect 23155 28580 23296 28608
rect 23155 28577 23167 28580
rect 23109 28571 23167 28577
rect 23290 28568 23296 28580
rect 23348 28568 23354 28620
rect 23474 28568 23480 28620
rect 23532 28608 23538 28620
rect 23569 28611 23627 28617
rect 23569 28608 23581 28611
rect 23532 28580 23581 28608
rect 23532 28568 23538 28580
rect 23569 28577 23581 28580
rect 23615 28577 23627 28611
rect 23569 28571 23627 28577
rect 27341 28611 27399 28617
rect 27341 28577 27353 28611
rect 27387 28608 27399 28611
rect 27522 28608 27528 28620
rect 27387 28580 27528 28608
rect 27387 28577 27399 28580
rect 27341 28571 27399 28577
rect 27522 28568 27528 28580
rect 27580 28568 27586 28620
rect 32585 28611 32643 28617
rect 32585 28577 32597 28611
rect 32631 28608 32643 28611
rect 33042 28608 33048 28620
rect 32631 28580 33048 28608
rect 32631 28577 32643 28580
rect 32585 28571 32643 28577
rect 33042 28568 33048 28580
rect 33100 28568 33106 28620
rect 33321 28611 33379 28617
rect 33321 28577 33333 28611
rect 33367 28608 33379 28611
rect 34057 28611 34115 28617
rect 34057 28608 34069 28611
rect 33367 28580 34069 28608
rect 33367 28577 33379 28580
rect 33321 28571 33379 28577
rect 34057 28577 34069 28580
rect 34103 28577 34115 28611
rect 34057 28571 34115 28577
rect 34514 28568 34520 28620
rect 34572 28608 34578 28620
rect 35253 28611 35311 28617
rect 35253 28608 35265 28611
rect 34572 28580 35265 28608
rect 34572 28568 34578 28580
rect 35253 28577 35265 28580
rect 35299 28577 35311 28611
rect 35253 28571 35311 28577
rect 36078 28568 36084 28620
rect 36136 28568 36142 28620
rect 38746 28568 38752 28620
rect 38804 28568 38810 28620
rect 39408 28608 39436 28639
rect 39776 28620 39804 28648
rect 40402 28636 40408 28648
rect 40460 28636 40466 28688
rect 39408 28580 39712 28608
rect 18969 28543 19027 28549
rect 18969 28540 18981 28543
rect 18840 28512 18981 28540
rect 18840 28500 18846 28512
rect 18969 28509 18981 28512
rect 19015 28509 19027 28543
rect 18969 28503 19027 28509
rect 19150 28500 19156 28552
rect 19208 28540 19214 28552
rect 19245 28543 19303 28549
rect 19245 28540 19257 28543
rect 19208 28512 19257 28540
rect 19208 28500 19214 28512
rect 19245 28509 19257 28512
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 21726 28500 21732 28552
rect 21784 28500 21790 28552
rect 22830 28500 22836 28552
rect 22888 28500 22894 28552
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28540 23811 28543
rect 23934 28540 23940 28552
rect 23799 28512 23940 28540
rect 23799 28509 23811 28512
rect 23753 28503 23811 28509
rect 23934 28500 23940 28512
rect 23992 28500 23998 28552
rect 24394 28500 24400 28552
rect 24452 28500 24458 28552
rect 24854 28500 24860 28552
rect 24912 28540 24918 28552
rect 24949 28543 25007 28549
rect 24949 28540 24961 28543
rect 24912 28512 24961 28540
rect 24912 28500 24918 28512
rect 24949 28509 24961 28512
rect 24995 28509 25007 28543
rect 24949 28503 25007 28509
rect 27065 28543 27123 28549
rect 27065 28509 27077 28543
rect 27111 28540 27123 28543
rect 28626 28540 28632 28552
rect 27111 28512 28632 28540
rect 27111 28509 27123 28512
rect 27065 28503 27123 28509
rect 28626 28500 28632 28512
rect 28684 28500 28690 28552
rect 32674 28500 32680 28552
rect 32732 28500 32738 28552
rect 33134 28500 33140 28552
rect 33192 28540 33198 28552
rect 33597 28543 33655 28549
rect 33597 28540 33609 28543
rect 33192 28512 33609 28540
rect 33192 28500 33198 28512
rect 33597 28509 33609 28512
rect 33643 28509 33655 28543
rect 33597 28503 33655 28509
rect 33778 28500 33784 28552
rect 33836 28540 33842 28552
rect 33836 28512 34100 28540
rect 33836 28500 33842 28512
rect 17957 28475 18015 28481
rect 17957 28472 17969 28475
rect 14476 28444 17969 28472
rect 17957 28441 17969 28444
rect 18003 28441 18015 28475
rect 17957 28435 18015 28441
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19521 28475 19579 28481
rect 19521 28472 19533 28475
rect 19484 28444 19533 28472
rect 19484 28432 19490 28444
rect 19521 28441 19533 28444
rect 19567 28441 19579 28475
rect 21821 28475 21879 28481
rect 19521 28435 19579 28441
rect 19628 28444 20010 28472
rect 6420 28376 7880 28404
rect 6420 28364 6426 28376
rect 8294 28364 8300 28416
rect 8352 28364 8358 28416
rect 8465 28407 8523 28413
rect 8465 28373 8477 28407
rect 8511 28404 8523 28407
rect 9030 28404 9036 28416
rect 8511 28376 9036 28404
rect 8511 28373 8523 28376
rect 8465 28367 8523 28373
rect 9030 28364 9036 28376
rect 9088 28364 9094 28416
rect 9309 28407 9367 28413
rect 9309 28373 9321 28407
rect 9355 28404 9367 28407
rect 9674 28404 9680 28416
rect 9355 28376 9680 28404
rect 9355 28373 9367 28376
rect 9309 28367 9367 28373
rect 9674 28364 9680 28376
rect 9732 28364 9738 28416
rect 13814 28364 13820 28416
rect 13872 28364 13878 28416
rect 14366 28364 14372 28416
rect 14424 28404 14430 28416
rect 14826 28404 14832 28416
rect 14424 28376 14832 28404
rect 14424 28364 14430 28376
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 17586 28364 17592 28416
rect 17644 28364 17650 28416
rect 17865 28407 17923 28413
rect 17865 28373 17877 28407
rect 17911 28404 17923 28407
rect 18157 28407 18215 28413
rect 18157 28404 18169 28407
rect 17911 28376 18169 28404
rect 17911 28373 17923 28376
rect 17865 28367 17923 28373
rect 18157 28373 18169 28376
rect 18203 28373 18215 28407
rect 18157 28367 18215 28373
rect 19242 28364 19248 28416
rect 19300 28404 19306 28416
rect 19628 28404 19656 28444
rect 21821 28441 21833 28475
rect 21867 28472 21879 28475
rect 22925 28475 22983 28481
rect 21867 28444 22094 28472
rect 21867 28441 21879 28444
rect 21821 28435 21879 28441
rect 19300 28376 19656 28404
rect 22066 28404 22094 28444
rect 22925 28441 22937 28475
rect 22971 28472 22983 28475
rect 23845 28475 23903 28481
rect 23845 28472 23857 28475
rect 22971 28444 23857 28472
rect 22971 28441 22983 28444
rect 22925 28435 22983 28441
rect 23845 28441 23857 28444
rect 23891 28472 23903 28475
rect 24412 28472 24440 28500
rect 23891 28444 24440 28472
rect 25216 28475 25274 28481
rect 23891 28441 23903 28444
rect 23845 28435 23903 28441
rect 25216 28441 25228 28475
rect 25262 28472 25274 28475
rect 25406 28472 25412 28484
rect 25262 28444 25412 28472
rect 25262 28441 25274 28444
rect 25216 28435 25274 28441
rect 25406 28432 25412 28444
rect 25464 28432 25470 28484
rect 27157 28475 27215 28481
rect 27157 28441 27169 28475
rect 27203 28441 27215 28475
rect 27157 28435 27215 28441
rect 23014 28404 23020 28416
rect 22066 28376 23020 28404
rect 19300 28364 19306 28376
rect 23014 28364 23020 28376
rect 23072 28404 23078 28416
rect 27172 28404 27200 28435
rect 31846 28432 31852 28484
rect 31904 28432 31910 28484
rect 32309 28475 32367 28481
rect 32309 28441 32321 28475
rect 32355 28472 32367 28475
rect 33413 28475 33471 28481
rect 33413 28472 33425 28475
rect 32355 28444 33425 28472
rect 32355 28441 32367 28444
rect 32309 28435 32367 28441
rect 33413 28441 33425 28444
rect 33459 28441 33471 28475
rect 33413 28435 33471 28441
rect 33689 28475 33747 28481
rect 33689 28441 33701 28475
rect 33735 28441 33747 28475
rect 33689 28435 33747 28441
rect 23072 28376 27200 28404
rect 30837 28407 30895 28413
rect 23072 28364 23078 28376
rect 30837 28373 30849 28407
rect 30883 28404 30895 28407
rect 32674 28404 32680 28416
rect 30883 28376 32680 28404
rect 30883 28373 30895 28376
rect 30837 28367 30895 28373
rect 32674 28364 32680 28376
rect 32732 28364 32738 28416
rect 33704 28404 33732 28435
rect 33870 28432 33876 28484
rect 33928 28481 33934 28484
rect 33928 28475 33957 28481
rect 33945 28441 33957 28475
rect 34072 28472 34100 28512
rect 34146 28500 34152 28552
rect 34204 28500 34210 28552
rect 34330 28500 34336 28552
rect 34388 28540 34394 28552
rect 35345 28543 35403 28549
rect 34388 28512 34652 28540
rect 34388 28500 34394 28512
rect 34624 28484 34652 28512
rect 35345 28509 35357 28543
rect 35391 28509 35403 28543
rect 35345 28503 35403 28509
rect 34072 28444 34284 28472
rect 33928 28435 33957 28441
rect 33928 28432 33934 28435
rect 34149 28407 34207 28413
rect 34149 28404 34161 28407
rect 33704 28376 34161 28404
rect 34149 28373 34161 28376
rect 34195 28373 34207 28407
rect 34256 28404 34284 28444
rect 34606 28432 34612 28484
rect 34664 28432 34670 28484
rect 35360 28472 35388 28503
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 35989 28543 36047 28549
rect 35989 28540 36001 28543
rect 35952 28512 36001 28540
rect 35952 28500 35958 28512
rect 35989 28509 36001 28512
rect 36035 28509 36047 28543
rect 36096 28540 36124 28568
rect 36173 28543 36231 28549
rect 36173 28540 36185 28543
rect 36096 28512 36185 28540
rect 35989 28503 36047 28509
rect 36173 28509 36185 28512
rect 36219 28509 36231 28543
rect 36173 28503 36231 28509
rect 38930 28500 38936 28552
rect 38988 28500 38994 28552
rect 39390 28500 39396 28552
rect 39448 28500 39454 28552
rect 36081 28475 36139 28481
rect 36081 28472 36093 28475
rect 35360 28444 36093 28472
rect 36081 28441 36093 28444
rect 36127 28441 36139 28475
rect 36081 28435 36139 28441
rect 35986 28404 35992 28416
rect 34256 28376 35992 28404
rect 34149 28367 34207 28373
rect 35986 28364 35992 28376
rect 36044 28364 36050 28416
rect 39684 28404 39712 28580
rect 39758 28568 39764 28620
rect 39816 28568 39822 28620
rect 40497 28611 40555 28617
rect 40497 28608 40509 28611
rect 40328 28580 40509 28608
rect 39776 28540 39804 28568
rect 40328 28552 40356 28580
rect 40497 28577 40509 28580
rect 40543 28577 40555 28611
rect 41386 28608 41414 28716
rect 42794 28704 42800 28756
rect 42852 28744 42858 28756
rect 43349 28747 43407 28753
rect 43349 28744 43361 28747
rect 42852 28716 43361 28744
rect 42852 28704 42858 28716
rect 43349 28713 43361 28716
rect 43395 28713 43407 28747
rect 43349 28707 43407 28713
rect 44082 28636 44088 28688
rect 44140 28676 44146 28688
rect 44177 28679 44235 28685
rect 44177 28676 44189 28679
rect 44140 28648 44189 28676
rect 44140 28636 44146 28648
rect 44177 28645 44189 28648
rect 44223 28645 44235 28679
rect 44177 28639 44235 28645
rect 42242 28608 42248 28620
rect 41386 28580 42248 28608
rect 40497 28571 40555 28577
rect 42242 28568 42248 28580
rect 42300 28608 42306 28620
rect 43438 28608 43444 28620
rect 42300 28580 43444 28608
rect 42300 28568 42306 28580
rect 43438 28568 43444 28580
rect 43496 28568 43502 28620
rect 39853 28543 39911 28549
rect 39853 28540 39865 28543
rect 39776 28512 39865 28540
rect 39853 28509 39865 28512
rect 39899 28509 39911 28543
rect 39853 28503 39911 28509
rect 40034 28500 40040 28552
rect 40092 28500 40098 28552
rect 40310 28500 40316 28552
rect 40368 28500 40374 28552
rect 40405 28543 40463 28549
rect 40405 28509 40417 28543
rect 40451 28540 40463 28543
rect 40586 28540 40592 28552
rect 40451 28512 40592 28540
rect 40451 28509 40463 28512
rect 40405 28503 40463 28509
rect 40586 28500 40592 28512
rect 40644 28500 40650 28552
rect 40862 28500 40868 28552
rect 40920 28500 40926 28552
rect 41690 28500 41696 28552
rect 41748 28540 41754 28552
rect 42061 28543 42119 28549
rect 42061 28540 42073 28543
rect 41748 28512 42073 28540
rect 41748 28500 41754 28512
rect 42061 28509 42073 28512
rect 42107 28509 42119 28543
rect 42061 28503 42119 28509
rect 43530 28500 43536 28552
rect 43588 28540 43594 28552
rect 43901 28543 43959 28549
rect 43901 28540 43913 28543
rect 43588 28512 43913 28540
rect 43588 28500 43594 28512
rect 43901 28509 43913 28512
rect 43947 28509 43959 28543
rect 43901 28503 43959 28509
rect 43990 28500 43996 28552
rect 44048 28540 44054 28552
rect 44177 28543 44235 28549
rect 44177 28540 44189 28543
rect 44048 28512 44189 28540
rect 44048 28500 44054 28512
rect 44177 28509 44189 28512
rect 44223 28509 44235 28543
rect 44177 28503 44235 28509
rect 39942 28432 39948 28484
rect 40000 28472 40006 28484
rect 40681 28475 40739 28481
rect 40681 28472 40693 28475
rect 40000 28444 40693 28472
rect 40000 28432 40006 28444
rect 40681 28441 40693 28444
rect 40727 28441 40739 28475
rect 40681 28435 40739 28441
rect 40880 28404 40908 28500
rect 43254 28432 43260 28484
rect 43312 28472 43318 28484
rect 44008 28472 44036 28500
rect 43312 28444 44036 28472
rect 43312 28432 43318 28444
rect 39684 28376 40908 28404
rect 42886 28364 42892 28416
rect 42944 28404 42950 28416
rect 43806 28404 43812 28416
rect 42944 28376 43812 28404
rect 42944 28364 42950 28376
rect 43806 28364 43812 28376
rect 43864 28404 43870 28416
rect 43993 28407 44051 28413
rect 43993 28404 44005 28407
rect 43864 28376 44005 28404
rect 43864 28364 43870 28376
rect 43993 28373 44005 28376
rect 44039 28404 44051 28407
rect 44174 28404 44180 28416
rect 44039 28376 44180 28404
rect 44039 28373 44051 28376
rect 43993 28367 44051 28373
rect 44174 28364 44180 28376
rect 44232 28364 44238 28416
rect 1104 28314 45172 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 45172 28314
rect 1104 28240 45172 28262
rect 3789 28203 3847 28209
rect 3789 28169 3801 28203
rect 3835 28200 3847 28203
rect 5258 28200 5264 28212
rect 3835 28172 5264 28200
rect 3835 28169 3847 28172
rect 3789 28163 3847 28169
rect 5258 28160 5264 28172
rect 5316 28160 5322 28212
rect 6178 28200 6184 28212
rect 5552 28172 6184 28200
rect 4798 28092 4804 28144
rect 4856 28092 4862 28144
rect 5552 28076 5580 28172
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 6546 28160 6552 28212
rect 6604 28200 6610 28212
rect 7653 28203 7711 28209
rect 6604 28172 6684 28200
rect 6604 28160 6610 28172
rect 5626 28092 5632 28144
rect 5684 28092 5690 28144
rect 5997 28135 6055 28141
rect 5997 28101 6009 28135
rect 6043 28132 6055 28135
rect 6043 28104 6592 28132
rect 6043 28101 6055 28104
rect 5997 28095 6055 28101
rect 934 28024 940 28076
rect 992 28064 998 28076
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 992 28036 1409 28064
rect 992 28024 998 28036
rect 1397 28033 1409 28036
rect 1443 28033 1455 28067
rect 1397 28027 1455 28033
rect 5534 28024 5540 28076
rect 5592 28024 5598 28076
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 5813 28067 5871 28073
rect 5813 28064 5825 28067
rect 5776 28036 5825 28064
rect 5776 28024 5782 28036
rect 5813 28033 5825 28036
rect 5859 28033 5871 28067
rect 5813 28027 5871 28033
rect 4798 27956 4804 28008
rect 4856 27996 4862 28008
rect 5261 27999 5319 28005
rect 5261 27996 5273 27999
rect 4856 27968 5273 27996
rect 4856 27956 4862 27968
rect 5261 27965 5273 27968
rect 5307 27965 5319 27999
rect 5828 27996 5856 28027
rect 6362 28024 6368 28076
rect 6420 28024 6426 28076
rect 6564 28073 6592 28104
rect 6656 28073 6684 28172
rect 7653 28169 7665 28203
rect 7699 28200 7711 28203
rect 7834 28200 7840 28212
rect 7699 28172 7840 28200
rect 7699 28169 7711 28172
rect 7653 28163 7711 28169
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 9030 28160 9036 28212
rect 9088 28200 9094 28212
rect 9398 28200 9404 28212
rect 9088 28172 9404 28200
rect 9088 28160 9094 28172
rect 9398 28160 9404 28172
rect 9456 28200 9462 28212
rect 14461 28203 14519 28209
rect 14461 28200 14473 28203
rect 9456 28172 14473 28200
rect 9456 28160 9462 28172
rect 7098 28092 7104 28144
rect 7156 28132 7162 28144
rect 7156 28104 7958 28132
rect 7156 28092 7162 28104
rect 9214 28092 9220 28144
rect 9272 28132 9278 28144
rect 9272 28104 9628 28132
rect 9272 28092 9278 28104
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28033 6699 28067
rect 6641 28027 6699 28033
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28064 6791 28067
rect 6822 28064 6828 28076
rect 6779 28036 6828 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 8110 28024 8116 28076
rect 8168 28024 8174 28076
rect 8128 27996 8156 28024
rect 5828 27968 8156 27996
rect 5261 27959 5319 27965
rect 9030 27956 9036 28008
rect 9088 27996 9094 28008
rect 9600 28005 9628 28104
rect 12434 28092 12440 28144
rect 12492 28092 12498 28144
rect 9950 28024 9956 28076
rect 10008 28024 10014 28076
rect 12452 28064 12480 28092
rect 12636 28073 12664 28172
rect 14461 28169 14473 28172
rect 14507 28169 14519 28203
rect 14624 28203 14682 28209
rect 14624 28200 14636 28203
rect 14461 28163 14519 28169
rect 14568 28172 14636 28200
rect 12710 28092 12716 28144
rect 12768 28092 12774 28144
rect 12897 28135 12955 28141
rect 12897 28132 12909 28135
rect 12820 28104 12909 28132
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 12452 28036 12541 28064
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 12621 28067 12679 28073
rect 12621 28033 12633 28067
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 9125 27999 9183 28005
rect 9125 27996 9137 27999
rect 9088 27968 9137 27996
rect 9088 27956 9094 27968
rect 9125 27965 9137 27968
rect 9171 27965 9183 27999
rect 9125 27959 9183 27965
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27965 9459 27999
rect 9401 27959 9459 27965
rect 9585 27999 9643 28005
rect 9585 27965 9597 27999
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 1762 27860 1768 27872
rect 1627 27832 1768 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 1762 27820 1768 27832
rect 1820 27820 1826 27872
rect 6914 27820 6920 27872
rect 6972 27860 6978 27872
rect 7009 27863 7067 27869
rect 7009 27860 7021 27863
rect 6972 27832 7021 27860
rect 6972 27820 6978 27832
rect 7009 27829 7021 27832
rect 7055 27829 7067 27863
rect 7009 27823 7067 27829
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 9416 27860 9444 27959
rect 11054 27956 11060 28008
rect 11112 27956 11118 28008
rect 11330 27956 11336 28008
rect 11388 27956 11394 28008
rect 12728 27996 12756 28092
rect 12820 28073 12848 28104
rect 12897 28101 12909 28104
rect 12943 28101 12955 28135
rect 12897 28095 12955 28101
rect 13446 28092 13452 28144
rect 13504 28092 13510 28144
rect 13538 28092 13544 28144
rect 13596 28132 13602 28144
rect 14274 28132 14280 28144
rect 13596 28104 14280 28132
rect 13596 28092 13602 28104
rect 14274 28092 14280 28104
rect 14332 28092 14338 28144
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28033 12863 28067
rect 12805 28027 12863 28033
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28064 13231 28067
rect 13464 28064 13492 28092
rect 13219 28036 13492 28064
rect 13219 28033 13231 28036
rect 13173 28027 13231 28033
rect 13630 28024 13636 28076
rect 13688 28024 13694 28076
rect 14185 28067 14243 28073
rect 14185 28033 14197 28067
rect 14231 28064 14243 28067
rect 14568 28064 14596 28172
rect 14624 28169 14636 28172
rect 14670 28169 14682 28203
rect 14624 28163 14682 28169
rect 17586 28160 17592 28212
rect 17644 28160 17650 28212
rect 21726 28160 21732 28212
rect 21784 28200 21790 28212
rect 21821 28203 21879 28209
rect 21821 28200 21833 28203
rect 21784 28172 21833 28200
rect 21784 28160 21790 28172
rect 21821 28169 21833 28172
rect 21867 28169 21879 28203
rect 21821 28163 21879 28169
rect 23661 28203 23719 28209
rect 23661 28169 23673 28203
rect 23707 28200 23719 28203
rect 23750 28200 23756 28212
rect 23707 28172 23756 28200
rect 23707 28169 23719 28172
rect 23661 28163 23719 28169
rect 23750 28160 23756 28172
rect 23808 28160 23814 28212
rect 24210 28160 24216 28212
rect 24268 28160 24274 28212
rect 25406 28160 25412 28212
rect 25464 28160 25470 28212
rect 25685 28203 25743 28209
rect 25685 28169 25697 28203
rect 25731 28200 25743 28203
rect 27430 28200 27436 28212
rect 25731 28172 27436 28200
rect 25731 28169 25743 28172
rect 25685 28163 25743 28169
rect 14826 28141 14832 28144
rect 14803 28135 14832 28141
rect 14803 28101 14815 28135
rect 14884 28132 14890 28144
rect 16022 28132 16028 28144
rect 14884 28104 16028 28132
rect 14803 28095 14832 28101
rect 14826 28092 14832 28095
rect 14884 28092 14890 28104
rect 16022 28092 16028 28104
rect 16080 28092 16086 28144
rect 15197 28067 15255 28073
rect 14231 28054 14596 28064
rect 14844 28054 15148 28064
rect 14231 28036 15148 28054
rect 14231 28033 14243 28036
rect 14185 28027 14243 28033
rect 14568 28026 14872 28036
rect 12897 27999 12955 28005
rect 12897 27996 12909 27999
rect 12728 27968 12909 27996
rect 12897 27965 12909 27968
rect 12943 27965 12955 27999
rect 12897 27959 12955 27965
rect 13004 27968 14136 27996
rect 12437 27931 12495 27937
rect 12437 27897 12449 27931
rect 12483 27928 12495 27931
rect 12526 27928 12532 27940
rect 12483 27900 12532 27928
rect 12483 27897 12495 27900
rect 12437 27891 12495 27897
rect 12526 27888 12532 27900
rect 12584 27928 12590 27940
rect 13004 27928 13032 27968
rect 12584 27900 13032 27928
rect 13081 27931 13139 27937
rect 12584 27888 12590 27900
rect 13081 27897 13093 27931
rect 13127 27928 13139 27931
rect 14108 27928 14136 27968
rect 14366 27956 14372 28008
rect 14424 27956 14430 28008
rect 14458 27956 14464 28008
rect 14516 27996 14522 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14516 27968 14933 27996
rect 14516 27956 14522 27968
rect 14921 27965 14933 27968
rect 14967 27965 14979 27999
rect 14921 27959 14979 27965
rect 15010 27956 15016 28008
rect 15068 27956 15074 28008
rect 15120 28005 15148 28036
rect 15197 28033 15209 28067
rect 15243 28064 15255 28067
rect 15746 28064 15752 28076
rect 15243 28036 15752 28064
rect 15243 28033 15255 28036
rect 15197 28027 15255 28033
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 17604 28064 17632 28160
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19996 28104 21588 28132
rect 18233 28067 18291 28073
rect 18233 28064 18245 28067
rect 17604 28036 18245 28064
rect 18233 28033 18245 28036
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 19150 28024 19156 28076
rect 19208 28054 19214 28076
rect 19996 28073 20024 28104
rect 21560 28076 21588 28104
rect 20254 28073 20260 28076
rect 19981 28067 20039 28073
rect 19981 28064 19993 28067
rect 19352 28054 19993 28064
rect 19208 28036 19993 28054
rect 19208 28026 19380 28036
rect 19981 28033 19993 28036
rect 20027 28033 20039 28067
rect 20248 28064 20260 28073
rect 20215 28036 20260 28064
rect 19981 28027 20039 28033
rect 20248 28027 20260 28036
rect 19208 28024 19214 28026
rect 20254 28024 20260 28027
rect 20312 28024 20318 28076
rect 21542 28024 21548 28076
rect 21600 28024 21606 28076
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28064 23903 28067
rect 24228 28064 24256 28160
rect 24949 28135 25007 28141
rect 24949 28101 24961 28135
rect 24995 28132 25007 28135
rect 25700 28132 25728 28163
rect 27430 28160 27436 28172
rect 27488 28160 27494 28212
rect 38930 28160 38936 28212
rect 38988 28160 38994 28212
rect 39758 28160 39764 28212
rect 39816 28160 39822 28212
rect 42886 28160 42892 28212
rect 42944 28160 42950 28212
rect 42978 28160 42984 28212
rect 43036 28160 43042 28212
rect 43346 28160 43352 28212
rect 43404 28160 43410 28212
rect 44082 28160 44088 28212
rect 44140 28160 44146 28212
rect 44174 28160 44180 28212
rect 44232 28200 44238 28212
rect 44269 28203 44327 28209
rect 44269 28200 44281 28203
rect 44232 28172 44281 28200
rect 44232 28160 44238 28172
rect 44269 28169 44281 28172
rect 44315 28169 44327 28203
rect 44269 28163 44327 28169
rect 24995 28104 25728 28132
rect 34793 28135 34851 28141
rect 24995 28101 25007 28104
rect 24949 28095 25007 28101
rect 34793 28101 34805 28135
rect 34839 28132 34851 28135
rect 35713 28135 35771 28141
rect 35713 28132 35725 28135
rect 34839 28104 35725 28132
rect 34839 28101 34851 28104
rect 34793 28095 34851 28101
rect 35713 28101 35725 28104
rect 35759 28132 35771 28135
rect 35759 28104 35940 28132
rect 35759 28101 35771 28104
rect 35713 28095 35771 28101
rect 25593 28067 25651 28073
rect 25593 28064 25605 28067
rect 23891 28036 24256 28064
rect 25332 28036 25605 28064
rect 23891 28033 23903 28036
rect 23845 28027 23903 28033
rect 15105 27999 15163 28005
rect 15105 27965 15117 27999
rect 15151 27996 15163 27999
rect 15378 27996 15384 28008
rect 15151 27968 15384 27996
rect 15151 27965 15163 27968
rect 15105 27959 15163 27965
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 17126 27956 17132 28008
rect 17184 27996 17190 28008
rect 17865 27999 17923 28005
rect 17865 27996 17877 27999
rect 17184 27968 17877 27996
rect 17184 27956 17190 27968
rect 17865 27965 17877 27968
rect 17911 27965 17923 27999
rect 17865 27959 17923 27965
rect 19058 27956 19064 28008
rect 19116 27996 19122 28008
rect 19705 27999 19763 28005
rect 19705 27996 19717 27999
rect 19116 27968 19717 27996
rect 19116 27956 19122 27968
rect 19705 27965 19717 27968
rect 19751 27965 19763 27999
rect 22373 27999 22431 28005
rect 22373 27996 22385 27999
rect 19705 27959 19763 27965
rect 22066 27968 22385 27996
rect 15028 27928 15056 27956
rect 13127 27900 14044 27928
rect 14108 27900 15056 27928
rect 21361 27931 21419 27937
rect 13127 27897 13139 27900
rect 13081 27891 13139 27897
rect 8444 27832 9444 27860
rect 8444 27820 8450 27832
rect 12802 27820 12808 27872
rect 12860 27820 12866 27872
rect 13541 27863 13599 27869
rect 13541 27829 13553 27863
rect 13587 27860 13599 27863
rect 13630 27860 13636 27872
rect 13587 27832 13636 27860
rect 13587 27829 13599 27832
rect 13541 27823 13599 27829
rect 13630 27820 13636 27832
rect 13688 27820 13694 27872
rect 14016 27869 14044 27900
rect 21361 27897 21373 27931
rect 21407 27928 21419 27931
rect 22066 27928 22094 27968
rect 22373 27965 22385 27968
rect 22419 27965 22431 27999
rect 22373 27959 22431 27965
rect 23474 27956 23480 28008
rect 23532 27996 23538 28008
rect 24670 27996 24676 28008
rect 23532 27968 24676 27996
rect 23532 27956 23538 27968
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 24854 27956 24860 28008
rect 24912 27956 24918 28008
rect 25332 27937 25360 28036
rect 25593 28033 25605 28036
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 26329 28067 26387 28073
rect 26329 28033 26341 28067
rect 26375 28064 26387 28067
rect 26418 28064 26424 28076
rect 26375 28036 26424 28064
rect 26375 28033 26387 28036
rect 26329 28027 26387 28033
rect 26418 28024 26424 28036
rect 26476 28024 26482 28076
rect 34698 28024 34704 28076
rect 34756 28064 34762 28076
rect 34977 28067 35035 28073
rect 34977 28064 34989 28067
rect 34756 28036 34989 28064
rect 34756 28024 34762 28036
rect 34977 28033 34989 28036
rect 35023 28033 35035 28067
rect 34977 28027 35035 28033
rect 35069 28067 35127 28073
rect 35069 28033 35081 28067
rect 35115 28033 35127 28067
rect 35069 28027 35127 28033
rect 35084 27996 35112 28027
rect 35250 28024 35256 28076
rect 35308 28024 35314 28076
rect 35345 28067 35403 28073
rect 35345 28033 35357 28067
rect 35391 28033 35403 28067
rect 35345 28027 35403 28033
rect 35360 27996 35388 28027
rect 35434 28024 35440 28076
rect 35492 28062 35498 28076
rect 35912 28073 35940 28104
rect 35621 28067 35679 28073
rect 35621 28064 35633 28067
rect 35544 28062 35633 28064
rect 35492 28036 35633 28062
rect 35492 28034 35572 28036
rect 35492 28024 35498 28034
rect 35621 28033 35633 28036
rect 35667 28033 35679 28067
rect 35621 28027 35679 28033
rect 35805 28067 35863 28073
rect 35805 28033 35817 28067
rect 35851 28033 35863 28067
rect 35805 28027 35863 28033
rect 35897 28067 35955 28073
rect 35897 28033 35909 28067
rect 35943 28033 35955 28067
rect 35897 28027 35955 28033
rect 35820 27996 35848 28027
rect 38838 28024 38844 28076
rect 38896 28024 38902 28076
rect 39025 28067 39083 28073
rect 39025 28033 39037 28067
rect 39071 28064 39083 28067
rect 39298 28064 39304 28076
rect 39071 28036 39304 28064
rect 39071 28033 39083 28036
rect 39025 28027 39083 28033
rect 39298 28024 39304 28036
rect 39356 28024 39362 28076
rect 39482 28024 39488 28076
rect 39540 28024 39546 28076
rect 40310 28024 40316 28076
rect 40368 28064 40374 28076
rect 41322 28064 41328 28076
rect 40368 28036 41328 28064
rect 40368 28024 40374 28036
rect 41322 28024 41328 28036
rect 41380 28064 41386 28076
rect 42429 28067 42487 28073
rect 42429 28064 42441 28067
rect 41380 28036 42441 28064
rect 41380 28024 41386 28036
rect 42429 28033 42441 28036
rect 42475 28033 42487 28067
rect 42429 28027 42487 28033
rect 42613 28067 42671 28073
rect 42613 28033 42625 28067
rect 42659 28064 42671 28067
rect 42904 28064 42932 28160
rect 42996 28132 43024 28160
rect 43364 28132 43392 28160
rect 44100 28132 44128 28160
rect 42996 28104 43300 28132
rect 43364 28104 43760 28132
rect 42659 28036 42932 28064
rect 42659 28033 42671 28036
rect 42613 28027 42671 28033
rect 42978 28024 42984 28076
rect 43036 28024 43042 28076
rect 43272 28064 43300 28104
rect 43732 28073 43760 28104
rect 44008 28104 44128 28132
rect 43441 28067 43499 28073
rect 43441 28064 43453 28067
rect 43272 28036 43453 28064
rect 43441 28033 43453 28036
rect 43487 28033 43499 28067
rect 43441 28027 43499 28033
rect 43717 28067 43775 28073
rect 43717 28033 43729 28067
rect 43763 28033 43775 28067
rect 43717 28027 43775 28033
rect 36722 27996 36728 28008
rect 35084 27968 35296 27996
rect 35360 27968 36728 27996
rect 21407 27900 22094 27928
rect 25317 27931 25375 27937
rect 21407 27897 21419 27900
rect 21361 27891 21419 27897
rect 25317 27897 25329 27931
rect 25363 27897 25375 27931
rect 25317 27891 25375 27897
rect 14001 27863 14059 27869
rect 14001 27829 14013 27863
rect 14047 27860 14059 27863
rect 14090 27860 14096 27872
rect 14047 27832 14096 27860
rect 14047 27829 14059 27832
rect 14001 27823 14059 27829
rect 14090 27820 14096 27832
rect 14148 27820 14154 27872
rect 14274 27820 14280 27872
rect 14332 27860 14338 27872
rect 14645 27863 14703 27869
rect 14645 27860 14657 27863
rect 14332 27832 14657 27860
rect 14332 27820 14338 27832
rect 14645 27829 14657 27832
rect 14691 27829 14703 27863
rect 14645 27823 14703 27829
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 15013 27863 15071 27869
rect 15013 27860 15025 27863
rect 14976 27832 15025 27860
rect 14976 27820 14982 27832
rect 15013 27829 15025 27832
rect 15059 27829 15071 27863
rect 15013 27823 15071 27829
rect 34790 27820 34796 27872
rect 34848 27820 34854 27872
rect 35268 27869 35296 27968
rect 36722 27956 36728 27968
rect 36780 27956 36786 28008
rect 42889 27999 42947 28005
rect 42889 27965 42901 27999
rect 42935 27996 42947 27999
rect 43254 27996 43260 28008
rect 42935 27968 43260 27996
rect 42935 27965 42947 27968
rect 42889 27959 42947 27965
rect 43254 27956 43260 27968
rect 43312 27956 43318 28008
rect 43456 27996 43484 28027
rect 43898 28024 43904 28076
rect 43956 28024 43962 28076
rect 44008 28073 44036 28104
rect 43993 28067 44051 28073
rect 43993 28033 44005 28067
rect 44039 28033 44051 28067
rect 43993 28027 44051 28033
rect 44085 28067 44143 28073
rect 44085 28033 44097 28067
rect 44131 28033 44143 28067
rect 44085 28027 44143 28033
rect 44361 28067 44419 28073
rect 44361 28033 44373 28067
rect 44407 28033 44419 28067
rect 44361 28027 44419 28033
rect 44100 27996 44128 28027
rect 43456 27968 44128 27996
rect 43162 27888 43168 27940
rect 43220 27928 43226 27940
rect 43349 27931 43407 27937
rect 43349 27928 43361 27931
rect 43220 27900 43361 27928
rect 43220 27888 43226 27900
rect 43349 27897 43361 27900
rect 43395 27897 43407 27931
rect 43349 27891 43407 27897
rect 43438 27888 43444 27940
rect 43496 27928 43502 27940
rect 44376 27928 44404 28027
rect 43496 27900 44404 27928
rect 43496 27888 43502 27900
rect 35253 27863 35311 27869
rect 35253 27829 35265 27863
rect 35299 27860 35311 27863
rect 35894 27860 35900 27872
rect 35299 27832 35900 27860
rect 35299 27829 35311 27832
rect 35253 27823 35311 27829
rect 35894 27820 35900 27832
rect 35952 27820 35958 27872
rect 35989 27863 36047 27869
rect 35989 27829 36001 27863
rect 36035 27860 36047 27863
rect 36078 27860 36084 27872
rect 36035 27832 36084 27860
rect 36035 27829 36047 27832
rect 35989 27823 36047 27829
rect 36078 27820 36084 27832
rect 36136 27820 36142 27872
rect 36170 27820 36176 27872
rect 36228 27820 36234 27872
rect 42978 27820 42984 27872
rect 43036 27860 43042 27872
rect 43533 27863 43591 27869
rect 43533 27860 43545 27863
rect 43036 27832 43545 27860
rect 43036 27820 43042 27832
rect 43533 27829 43545 27832
rect 43579 27829 43591 27863
rect 43533 27823 43591 27829
rect 44085 27863 44143 27869
rect 44085 27829 44097 27863
rect 44131 27860 44143 27863
rect 44174 27860 44180 27872
rect 44131 27832 44180 27860
rect 44131 27829 44143 27832
rect 44085 27823 44143 27829
rect 44174 27820 44180 27832
rect 44232 27820 44238 27872
rect 1104 27770 45172 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 45172 27770
rect 1104 27696 45172 27718
rect 4798 27616 4804 27668
rect 4856 27616 4862 27668
rect 5442 27616 5448 27668
rect 5500 27616 5506 27668
rect 5626 27616 5632 27668
rect 5684 27616 5690 27668
rect 5813 27659 5871 27665
rect 5813 27625 5825 27659
rect 5859 27656 5871 27659
rect 6546 27656 6552 27668
rect 5859 27628 6552 27656
rect 5859 27625 5871 27628
rect 5813 27619 5871 27625
rect 5261 27591 5319 27597
rect 5261 27557 5273 27591
rect 5307 27557 5319 27591
rect 5261 27551 5319 27557
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27452 4675 27455
rect 5276 27452 5304 27551
rect 4663 27424 5304 27452
rect 5644 27452 5672 27616
rect 5721 27455 5779 27461
rect 5721 27452 5733 27455
rect 5644 27424 5733 27452
rect 4663 27421 4675 27424
rect 4617 27415 4675 27421
rect 5721 27421 5733 27424
rect 5767 27421 5779 27455
rect 5721 27415 5779 27421
rect 5626 27344 5632 27396
rect 5684 27344 5690 27396
rect 5429 27319 5487 27325
rect 5429 27285 5441 27319
rect 5475 27316 5487 27319
rect 5828 27316 5856 27619
rect 6546 27616 6552 27628
rect 6604 27616 6610 27668
rect 8294 27616 8300 27668
rect 8352 27656 8358 27668
rect 8846 27656 8852 27668
rect 8352 27628 8852 27656
rect 8352 27616 8358 27628
rect 8846 27616 8852 27628
rect 8904 27616 8910 27668
rect 9033 27659 9091 27665
rect 9033 27625 9045 27659
rect 9079 27656 9091 27659
rect 9122 27656 9128 27668
rect 9079 27628 9128 27656
rect 9079 27625 9091 27628
rect 9033 27619 9091 27625
rect 9122 27616 9128 27628
rect 9180 27616 9186 27668
rect 11054 27616 11060 27668
rect 11112 27616 11118 27668
rect 12332 27659 12390 27665
rect 12332 27625 12344 27659
rect 12378 27656 12390 27659
rect 12802 27656 12808 27668
rect 12378 27628 12808 27656
rect 12378 27625 12390 27628
rect 12332 27619 12390 27625
rect 12802 27616 12808 27628
rect 12860 27616 12866 27668
rect 13446 27616 13452 27668
rect 13504 27656 13510 27668
rect 13817 27659 13875 27665
rect 13817 27656 13829 27659
rect 13504 27628 13829 27656
rect 13504 27616 13510 27628
rect 13817 27625 13829 27628
rect 13863 27656 13875 27659
rect 14274 27656 14280 27668
rect 13863 27628 14280 27656
rect 13863 27625 13875 27628
rect 13817 27619 13875 27625
rect 14274 27616 14280 27628
rect 14332 27616 14338 27668
rect 16022 27616 16028 27668
rect 16080 27616 16086 27668
rect 21542 27616 21548 27668
rect 21600 27656 21606 27668
rect 26605 27659 26663 27665
rect 21600 27628 22140 27656
rect 21600 27616 21606 27628
rect 10229 27591 10287 27597
rect 10229 27557 10241 27591
rect 10275 27588 10287 27591
rect 11072 27588 11100 27616
rect 22005 27591 22063 27597
rect 22005 27588 22017 27591
rect 10275 27560 11100 27588
rect 21744 27560 22017 27588
rect 10275 27557 10287 27560
rect 10229 27551 10287 27557
rect 11330 27480 11336 27532
rect 11388 27520 11394 27532
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 11388 27492 12081 27520
rect 11388 27480 11394 27492
rect 12069 27489 12081 27492
rect 12115 27520 12127 27523
rect 13722 27520 13728 27532
rect 12115 27492 13728 27520
rect 12115 27489 12127 27492
rect 12069 27483 12127 27489
rect 13722 27480 13728 27492
rect 13780 27520 13786 27532
rect 14277 27523 14335 27529
rect 14277 27520 14289 27523
rect 13780 27492 14289 27520
rect 13780 27480 13786 27492
rect 14277 27489 14289 27492
rect 14323 27520 14335 27523
rect 16666 27520 16672 27532
rect 14323 27492 16672 27520
rect 14323 27489 14335 27492
rect 14277 27483 14335 27489
rect 16666 27480 16672 27492
rect 16724 27480 16730 27532
rect 7006 27412 7012 27464
rect 7064 27412 7070 27464
rect 9214 27412 9220 27464
rect 9272 27412 9278 27464
rect 9398 27412 9404 27464
rect 9456 27412 9462 27464
rect 9674 27412 9680 27464
rect 9732 27452 9738 27464
rect 10045 27455 10103 27461
rect 10045 27452 10057 27455
rect 9732 27424 10057 27452
rect 9732 27412 9738 27424
rect 10045 27421 10057 27424
rect 10091 27421 10103 27455
rect 19889 27455 19947 27461
rect 19889 27452 19901 27455
rect 10045 27415 10103 27421
rect 19260 27424 19901 27452
rect 13630 27384 13636 27396
rect 13570 27356 13636 27384
rect 13630 27344 13636 27356
rect 13688 27344 13694 27396
rect 14550 27344 14556 27396
rect 14608 27344 14614 27396
rect 18138 27384 18144 27396
rect 15778 27356 18144 27384
rect 5475 27288 5856 27316
rect 5475 27285 5487 27288
rect 5429 27279 5487 27285
rect 8202 27276 8208 27328
rect 8260 27316 8266 27328
rect 8297 27319 8355 27325
rect 8297 27316 8309 27319
rect 8260 27288 8309 27316
rect 8260 27276 8266 27288
rect 8297 27285 8309 27288
rect 8343 27316 8355 27319
rect 8386 27316 8392 27328
rect 8343 27288 8392 27316
rect 8343 27285 8355 27288
rect 8297 27279 8355 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 13648 27316 13676 27344
rect 15856 27316 15884 27356
rect 18138 27344 18144 27356
rect 18196 27344 18202 27396
rect 13648 27288 15884 27316
rect 16298 27276 16304 27328
rect 16356 27316 16362 27328
rect 19260 27316 19288 27424
rect 19889 27421 19901 27424
rect 19935 27452 19947 27455
rect 20806 27452 20812 27464
rect 19935 27424 20812 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 20806 27412 20812 27424
rect 20864 27412 20870 27464
rect 20165 27387 20223 27393
rect 20165 27353 20177 27387
rect 20211 27353 20223 27387
rect 21744 27384 21772 27560
rect 22005 27557 22017 27560
rect 22051 27557 22063 27591
rect 22005 27551 22063 27557
rect 22112 27529 22140 27628
rect 26605 27625 26617 27659
rect 26651 27656 26663 27659
rect 26954 27659 27012 27665
rect 26954 27656 26966 27659
rect 26651 27628 26966 27656
rect 26651 27625 26663 27628
rect 26605 27619 26663 27625
rect 26954 27625 26966 27628
rect 27000 27625 27012 27659
rect 26954 27619 27012 27625
rect 27706 27616 27712 27668
rect 27764 27656 27770 27668
rect 31846 27656 31852 27668
rect 27764 27628 31852 27656
rect 27764 27616 27770 27628
rect 31846 27616 31852 27628
rect 31904 27616 31910 27668
rect 34514 27616 34520 27668
rect 34572 27616 34578 27668
rect 36722 27616 36728 27668
rect 36780 27616 36786 27668
rect 36814 27616 36820 27668
rect 36872 27656 36878 27668
rect 38209 27659 38267 27665
rect 38209 27656 38221 27659
rect 36872 27628 38221 27656
rect 36872 27616 36878 27628
rect 38209 27625 38221 27628
rect 38255 27625 38267 27659
rect 38209 27619 38267 27625
rect 39393 27659 39451 27665
rect 39393 27625 39405 27659
rect 39439 27656 39451 27659
rect 39482 27656 39488 27668
rect 39439 27628 39488 27656
rect 39439 27625 39451 27628
rect 39393 27619 39451 27625
rect 39482 27616 39488 27628
rect 39540 27616 39546 27668
rect 43070 27616 43076 27668
rect 43128 27656 43134 27668
rect 43438 27656 43444 27668
rect 43128 27628 43444 27656
rect 43128 27616 43134 27628
rect 43438 27616 43444 27628
rect 43496 27616 43502 27668
rect 23106 27548 23112 27600
rect 23164 27588 23170 27600
rect 23477 27591 23535 27597
rect 23477 27588 23489 27591
rect 23164 27560 23489 27588
rect 23164 27548 23170 27560
rect 23477 27557 23489 27560
rect 23523 27557 23535 27591
rect 23477 27551 23535 27557
rect 34425 27591 34483 27597
rect 34425 27557 34437 27591
rect 34471 27588 34483 27591
rect 34532 27588 34560 27616
rect 34471 27560 34560 27588
rect 34701 27591 34759 27597
rect 34471 27557 34483 27560
rect 34425 27551 34483 27557
rect 34701 27557 34713 27591
rect 34747 27588 34759 27591
rect 34790 27588 34796 27600
rect 34747 27560 34796 27588
rect 34747 27557 34759 27560
rect 34701 27551 34759 27557
rect 34790 27548 34796 27560
rect 34848 27548 34854 27600
rect 39298 27548 39304 27600
rect 39356 27588 39362 27600
rect 39758 27588 39764 27600
rect 39356 27560 39764 27588
rect 39356 27548 39362 27560
rect 39758 27548 39764 27560
rect 39816 27548 39822 27600
rect 22097 27523 22155 27529
rect 22097 27489 22109 27523
rect 22143 27489 22155 27523
rect 22097 27483 22155 27489
rect 24670 27480 24676 27532
rect 24728 27520 24734 27532
rect 24949 27523 25007 27529
rect 24949 27520 24961 27523
rect 24728 27492 24961 27520
rect 24728 27480 24734 27492
rect 24949 27489 24961 27492
rect 24995 27489 25007 27523
rect 24949 27483 25007 27489
rect 26697 27523 26755 27529
rect 26697 27489 26709 27523
rect 26743 27520 26755 27523
rect 26970 27520 26976 27532
rect 26743 27492 26976 27520
rect 26743 27489 26755 27492
rect 26697 27483 26755 27489
rect 26970 27480 26976 27492
rect 27028 27480 27034 27532
rect 34606 27480 34612 27532
rect 34664 27520 34670 27532
rect 35069 27523 35127 27529
rect 35069 27520 35081 27523
rect 34664 27492 35081 27520
rect 34664 27480 34670 27492
rect 35069 27489 35081 27492
rect 35115 27489 35127 27523
rect 35069 27483 35127 27489
rect 38473 27523 38531 27529
rect 38473 27489 38485 27523
rect 38519 27520 38531 27523
rect 42794 27520 42800 27532
rect 38519 27492 42800 27520
rect 38519 27489 38531 27492
rect 38473 27483 38531 27489
rect 42794 27480 42800 27492
rect 42852 27480 42858 27532
rect 21821 27455 21879 27461
rect 21821 27421 21833 27455
rect 21867 27452 21879 27455
rect 22186 27452 22192 27464
rect 21867 27424 22192 27452
rect 21867 27421 21879 27424
rect 21821 27415 21879 27421
rect 22186 27412 22192 27424
rect 22244 27412 22250 27464
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 24029 27455 24087 27461
rect 22704 27424 23704 27452
rect 22704 27412 22710 27424
rect 23676 27393 23704 27424
rect 24029 27421 24041 27455
rect 24075 27452 24087 27455
rect 24578 27452 24584 27464
rect 24075 27424 24584 27452
rect 24075 27421 24087 27424
rect 24029 27415 24087 27421
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27452 24823 27455
rect 25498 27452 25504 27464
rect 24811 27424 25504 27452
rect 24811 27421 24823 27424
rect 24765 27415 24823 27421
rect 25498 27412 25504 27424
rect 25556 27412 25562 27464
rect 26418 27412 26424 27464
rect 26476 27412 26482 27464
rect 34330 27412 34336 27464
rect 34388 27412 34394 27464
rect 34517 27455 34575 27461
rect 34517 27421 34529 27455
rect 34563 27452 34575 27455
rect 34563 27424 34744 27452
rect 34563 27421 34575 27424
rect 34517 27415 34575 27421
rect 22342 27387 22400 27393
rect 22342 27384 22354 27387
rect 21744 27356 22354 27384
rect 20165 27347 20223 27353
rect 22342 27353 22354 27356
rect 22388 27353 22400 27387
rect 22342 27347 22400 27353
rect 23661 27387 23719 27393
rect 23661 27353 23673 27387
rect 23707 27353 23719 27387
rect 23661 27347 23719 27353
rect 24320 27356 27108 27384
rect 16356 27288 19288 27316
rect 16356 27276 16362 27288
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 20180 27316 20208 27347
rect 24320 27316 24348 27356
rect 19392 27288 24348 27316
rect 19392 27276 19398 27288
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 24857 27319 24915 27325
rect 24857 27285 24869 27319
rect 24903 27316 24915 27319
rect 25038 27316 25044 27328
rect 24903 27288 25044 27316
rect 24903 27285 24915 27288
rect 24857 27279 24915 27285
rect 25038 27276 25044 27288
rect 25096 27276 25102 27328
rect 27080 27316 27108 27356
rect 27706 27344 27712 27396
rect 27764 27344 27770 27396
rect 28276 27356 30696 27384
rect 28276 27316 28304 27356
rect 30668 27328 30696 27356
rect 34716 27328 34744 27424
rect 35250 27412 35256 27464
rect 35308 27412 35314 27464
rect 35434 27412 35440 27464
rect 35492 27452 35498 27464
rect 35621 27455 35679 27461
rect 35621 27452 35633 27455
rect 35492 27424 35633 27452
rect 35492 27412 35498 27424
rect 35621 27421 35633 27424
rect 35667 27421 35679 27455
rect 35621 27415 35679 27421
rect 35894 27412 35900 27464
rect 35952 27452 35958 27464
rect 35989 27455 36047 27461
rect 35989 27452 36001 27455
rect 35952 27424 36001 27452
rect 35952 27412 35958 27424
rect 35989 27421 36001 27424
rect 36035 27421 36047 27455
rect 35989 27415 36047 27421
rect 36078 27412 36084 27464
rect 36136 27452 36142 27464
rect 36357 27455 36415 27461
rect 36357 27452 36369 27455
rect 36136 27424 36369 27452
rect 36136 27412 36142 27424
rect 36357 27421 36369 27424
rect 36403 27421 36415 27455
rect 36357 27415 36415 27421
rect 36906 27412 36912 27464
rect 36964 27452 36970 27464
rect 39853 27455 39911 27461
rect 39853 27452 39865 27455
rect 36964 27424 37122 27452
rect 38948 27424 39865 27452
rect 36964 27412 36970 27424
rect 35268 27384 35296 27412
rect 35268 27356 36400 27384
rect 36372 27328 36400 27356
rect 38838 27344 38844 27396
rect 38896 27384 38902 27396
rect 38948 27393 38976 27424
rect 39853 27421 39865 27424
rect 39899 27421 39911 27455
rect 39853 27415 39911 27421
rect 40310 27412 40316 27464
rect 40368 27412 40374 27464
rect 40497 27455 40555 27461
rect 40497 27421 40509 27455
rect 40543 27421 40555 27455
rect 40497 27415 40555 27421
rect 38933 27387 38991 27393
rect 38933 27384 38945 27387
rect 38896 27356 38945 27384
rect 38896 27344 38902 27356
rect 38933 27353 38945 27356
rect 38979 27353 38991 27387
rect 38933 27347 38991 27353
rect 39758 27344 39764 27396
rect 39816 27384 39822 27396
rect 40512 27384 40540 27415
rect 39816 27356 40540 27384
rect 39816 27344 39822 27356
rect 27080 27288 28304 27316
rect 28442 27276 28448 27328
rect 28500 27276 28506 27328
rect 30650 27276 30656 27328
rect 30708 27276 30714 27328
rect 34698 27276 34704 27328
rect 34756 27276 34762 27328
rect 36354 27276 36360 27328
rect 36412 27276 36418 27328
rect 1104 27226 45172 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 45172 27226
rect 1104 27152 45172 27174
rect 8389 27115 8447 27121
rect 8389 27081 8401 27115
rect 8435 27112 8447 27115
rect 8478 27112 8484 27124
rect 8435 27084 8484 27112
rect 8435 27081 8447 27084
rect 8389 27075 8447 27081
rect 8478 27072 8484 27084
rect 8536 27072 8542 27124
rect 8570 27072 8576 27124
rect 8628 27072 8634 27124
rect 8941 27115 8999 27121
rect 8941 27081 8953 27115
rect 8987 27112 8999 27115
rect 9030 27112 9036 27124
rect 8987 27084 9036 27112
rect 8987 27081 8999 27084
rect 8941 27075 8999 27081
rect 9030 27072 9036 27084
rect 9088 27072 9094 27124
rect 13446 27072 13452 27124
rect 13504 27112 13510 27124
rect 13722 27112 13728 27124
rect 13504 27084 13728 27112
rect 13504 27072 13510 27084
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 14550 27072 14556 27124
rect 14608 27112 14614 27124
rect 14921 27115 14979 27121
rect 14921 27112 14933 27115
rect 14608 27084 14933 27112
rect 14608 27072 14614 27084
rect 14921 27081 14933 27084
rect 14967 27081 14979 27115
rect 14921 27075 14979 27081
rect 22186 27072 22192 27124
rect 22244 27112 22250 27124
rect 22373 27115 22431 27121
rect 22373 27112 22385 27115
rect 22244 27084 22385 27112
rect 22244 27072 22250 27084
rect 22373 27081 22385 27084
rect 22419 27081 22431 27115
rect 22373 27075 22431 27081
rect 22741 27115 22799 27121
rect 22741 27081 22753 27115
rect 22787 27112 22799 27115
rect 23106 27112 23112 27124
rect 22787 27084 23112 27112
rect 22787 27081 22799 27084
rect 22741 27075 22799 27081
rect 23106 27072 23112 27084
rect 23164 27072 23170 27124
rect 24394 27112 24400 27124
rect 24136 27084 24400 27112
rect 6641 27047 6699 27053
rect 6641 27013 6653 27047
rect 6687 27044 6699 27047
rect 6914 27044 6920 27056
rect 6687 27016 6920 27044
rect 6687 27013 6699 27016
rect 6641 27007 6699 27013
rect 6914 27004 6920 27016
rect 6972 27004 6978 27056
rect 7098 27004 7104 27056
rect 7156 27004 7162 27056
rect 8588 27044 8616 27072
rect 8588 27016 9076 27044
rect 5534 26936 5540 26988
rect 5592 26976 5598 26988
rect 6365 26979 6423 26985
rect 6365 26976 6377 26979
rect 5592 26948 6377 26976
rect 5592 26936 5598 26948
rect 6365 26945 6377 26948
rect 6411 26945 6423 26979
rect 6365 26939 6423 26945
rect 6380 26908 6408 26939
rect 8202 26936 8208 26988
rect 8260 26936 8266 26988
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 8220 26908 8248 26936
rect 6380 26880 8248 26908
rect 8110 26800 8116 26852
rect 8168 26800 8174 26852
rect 8588 26840 8616 26939
rect 8846 26936 8852 26988
rect 8904 26936 8910 26988
rect 9048 26985 9076 27016
rect 14734 27004 14740 27056
rect 14792 27004 14798 27056
rect 20622 27044 20628 27056
rect 20548 27016 20628 27044
rect 9033 26979 9091 26985
rect 9033 26945 9045 26979
rect 9079 26945 9091 26979
rect 9033 26939 9091 26945
rect 9214 26936 9220 26988
rect 9272 26936 9278 26988
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 14829 26979 14887 26985
rect 14829 26976 14841 26979
rect 14148 26948 14841 26976
rect 14148 26936 14154 26948
rect 14829 26945 14841 26948
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 14918 26936 14924 26988
rect 14976 26976 14982 26988
rect 20548 26985 20576 27016
rect 20622 27004 20628 27016
rect 20680 27004 20686 27056
rect 22462 27044 22468 27056
rect 20732 27016 22468 27044
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14976 26948 15025 26976
rect 14976 26936 14982 26948
rect 15013 26945 15025 26948
rect 15059 26945 15071 26979
rect 15013 26939 15071 26945
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 8757 26911 8815 26917
rect 8757 26877 8769 26911
rect 8803 26908 8815 26911
rect 9232 26908 9260 26936
rect 8803 26880 9260 26908
rect 8803 26877 8815 26880
rect 8757 26871 8815 26877
rect 9398 26868 9404 26920
rect 9456 26868 9462 26920
rect 12066 26868 12072 26920
rect 12124 26868 12130 26920
rect 9416 26840 9444 26868
rect 8588 26812 9444 26840
rect 18156 26840 18184 26939
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 20732 26917 20760 27016
rect 22462 27004 22468 27016
rect 22520 27044 22526 27056
rect 22520 27016 23060 27044
rect 22520 27004 22526 27016
rect 20806 26936 20812 26988
rect 20864 26976 20870 26988
rect 22646 26976 22652 26988
rect 20864 26948 22652 26976
rect 20864 26936 20870 26948
rect 22646 26936 22652 26948
rect 22704 26936 22710 26988
rect 20717 26911 20775 26917
rect 20717 26908 20729 26911
rect 20680 26880 20729 26908
rect 20680 26868 20686 26880
rect 20717 26877 20729 26880
rect 20763 26877 20775 26911
rect 20717 26871 20775 26877
rect 22830 26868 22836 26920
rect 22888 26868 22894 26920
rect 23032 26917 23060 27016
rect 24136 26985 24164 27084
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 25774 27072 25780 27124
rect 25832 27072 25838 27124
rect 26418 27072 26424 27124
rect 26476 27112 26482 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26476 27084 26985 27112
rect 26476 27072 26482 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 27341 27115 27399 27121
rect 27341 27081 27353 27115
rect 27387 27112 27399 27115
rect 28442 27112 28448 27124
rect 27387 27084 28448 27112
rect 27387 27081 27399 27084
rect 27341 27075 27399 27081
rect 28442 27072 28448 27084
rect 28500 27072 28506 27124
rect 28997 27115 29055 27121
rect 28997 27081 29009 27115
rect 29043 27081 29055 27115
rect 28997 27075 29055 27081
rect 24762 27044 24768 27056
rect 24412 27016 24768 27044
rect 24412 26985 24440 27016
rect 24762 27004 24768 27016
rect 24820 27004 24826 27056
rect 29012 27044 29040 27075
rect 29270 27072 29276 27124
rect 29328 27112 29334 27124
rect 30098 27112 30104 27124
rect 29328 27084 30104 27112
rect 29328 27072 29334 27084
rect 30098 27072 30104 27084
rect 30156 27072 30162 27124
rect 34330 27072 34336 27124
rect 34388 27072 34394 27124
rect 35250 27072 35256 27124
rect 35308 27072 35314 27124
rect 35529 27115 35587 27121
rect 35529 27081 35541 27115
rect 35575 27112 35587 27115
rect 36814 27112 36820 27124
rect 35575 27084 36820 27112
rect 35575 27081 35587 27084
rect 35529 27075 35587 27081
rect 36814 27072 36820 27084
rect 36872 27072 36878 27124
rect 43162 27072 43168 27124
rect 43220 27112 43226 27124
rect 43220 27084 43760 27112
rect 43220 27072 43226 27084
rect 34348 27044 34376 27072
rect 29012 27016 30512 27044
rect 34348 27016 35204 27044
rect 24121 26979 24179 26985
rect 24121 26945 24133 26979
rect 24167 26945 24179 26979
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24121 26939 24179 26945
rect 24320 26948 24409 26976
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26908 23075 26911
rect 23474 26908 23480 26920
rect 23063 26880 23480 26908
rect 23063 26877 23075 26880
rect 23017 26871 23075 26877
rect 23474 26868 23480 26880
rect 23532 26868 23538 26920
rect 24320 26908 24348 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24653 26979 24711 26985
rect 24653 26976 24665 26979
rect 24397 26939 24455 26945
rect 24504 26948 24665 26976
rect 24504 26908 24532 26948
rect 24653 26945 24665 26948
rect 24699 26945 24711 26979
rect 24653 26939 24711 26945
rect 28629 26979 28687 26985
rect 28629 26945 28641 26979
rect 28675 26945 28687 26979
rect 28629 26939 28687 26945
rect 24136 26880 24348 26908
rect 24412 26880 24532 26908
rect 24136 26852 24164 26880
rect 21358 26840 21364 26852
rect 18156 26812 21364 26840
rect 21358 26800 21364 26812
rect 21416 26800 21422 26852
rect 24118 26800 24124 26852
rect 24176 26800 24182 26852
rect 24305 26843 24363 26849
rect 24305 26809 24317 26843
rect 24351 26840 24363 26843
rect 24412 26840 24440 26880
rect 27430 26868 27436 26920
rect 27488 26868 27494 26920
rect 27522 26868 27528 26920
rect 27580 26868 27586 26920
rect 28644 26852 28672 26939
rect 28994 26936 29000 26988
rect 29052 26976 29058 26988
rect 29365 26979 29423 26985
rect 29365 26976 29377 26979
rect 29052 26948 29377 26976
rect 29052 26936 29058 26948
rect 29365 26945 29377 26948
rect 29411 26945 29423 26979
rect 30484 26974 30512 27016
rect 30561 26979 30619 26985
rect 30561 26974 30573 26979
rect 30484 26946 30573 26974
rect 29365 26939 29423 26945
rect 30561 26945 30573 26946
rect 30607 26945 30619 26979
rect 30561 26939 30619 26945
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 34609 26979 34667 26985
rect 30708 26948 34560 26976
rect 30708 26936 30714 26948
rect 28721 26911 28779 26917
rect 28721 26877 28733 26911
rect 28767 26908 28779 26911
rect 28810 26908 28816 26920
rect 28767 26880 28816 26908
rect 28767 26877 28779 26880
rect 28721 26871 28779 26877
rect 28810 26868 28816 26880
rect 28868 26868 28874 26920
rect 29638 26868 29644 26920
rect 29696 26868 29702 26920
rect 30193 26911 30251 26917
rect 30193 26877 30205 26911
rect 30239 26908 30251 26911
rect 34333 26911 34391 26917
rect 34333 26908 34345 26911
rect 30239 26880 34345 26908
rect 30239 26877 30251 26880
rect 30193 26871 30251 26877
rect 34333 26877 34345 26880
rect 34379 26908 34391 26911
rect 34422 26908 34428 26920
rect 34379 26880 34428 26908
rect 34379 26877 34391 26880
rect 34333 26871 34391 26877
rect 34422 26868 34428 26880
rect 34480 26868 34486 26920
rect 34532 26908 34560 26948
rect 34609 26945 34621 26979
rect 34655 26976 34667 26979
rect 34790 26976 34796 26988
rect 34655 26948 34796 26976
rect 34655 26945 34667 26948
rect 34609 26939 34667 26945
rect 34790 26936 34796 26948
rect 34848 26936 34854 26988
rect 35176 26976 35204 27016
rect 35618 27004 35624 27056
rect 35676 27044 35682 27056
rect 36015 27047 36073 27053
rect 36015 27044 36027 27047
rect 35676 27016 36027 27044
rect 35676 27004 35682 27016
rect 36015 27013 36027 27016
rect 36061 27013 36073 27047
rect 36015 27007 36073 27013
rect 36354 27004 36360 27056
rect 36412 27004 36418 27056
rect 43732 27053 43760 27084
rect 42613 27047 42671 27053
rect 42613 27013 42625 27047
rect 42659 27013 42671 27047
rect 42613 27007 42671 27013
rect 43717 27047 43775 27053
rect 43717 27013 43729 27047
rect 43763 27013 43775 27047
rect 43717 27007 43775 27013
rect 35713 26979 35771 26985
rect 35713 26976 35725 26979
rect 35176 26948 35725 26976
rect 35713 26945 35725 26948
rect 35759 26945 35771 26979
rect 35713 26939 35771 26945
rect 34532 26880 35296 26908
rect 28626 26840 28632 26852
rect 24351 26812 24440 26840
rect 26160 26812 28632 26840
rect 24351 26809 24363 26812
rect 24305 26803 24363 26809
rect 26160 26784 26188 26812
rect 28626 26800 28632 26812
rect 28684 26800 28690 26852
rect 30653 26843 30711 26849
rect 30653 26809 30665 26843
rect 30699 26840 30711 26843
rect 35158 26840 35164 26852
rect 30699 26812 35164 26840
rect 30699 26809 30711 26812
rect 30653 26803 30711 26809
rect 35158 26800 35164 26812
rect 35216 26800 35222 26852
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 17954 26732 17960 26784
rect 18012 26732 18018 26784
rect 26142 26732 26148 26784
rect 26200 26732 26206 26784
rect 35268 26772 35296 26880
rect 35434 26868 35440 26920
rect 35492 26868 35498 26920
rect 35728 26908 35756 26939
rect 35802 26936 35808 26988
rect 35860 26936 35866 26988
rect 35894 26936 35900 26988
rect 35952 26936 35958 26988
rect 36170 26936 36176 26988
rect 36228 26936 36234 26988
rect 36265 26979 36323 26985
rect 36265 26945 36277 26979
rect 36311 26976 36323 26979
rect 36372 26976 36400 27004
rect 36311 26948 36400 26976
rect 36449 26979 36507 26985
rect 36311 26945 36323 26948
rect 36265 26939 36323 26945
rect 36449 26945 36461 26979
rect 36495 26945 36507 26979
rect 36449 26939 36507 26945
rect 36357 26911 36415 26917
rect 36357 26908 36369 26911
rect 35728 26880 36369 26908
rect 36357 26877 36369 26880
rect 36403 26877 36415 26911
rect 36357 26871 36415 26877
rect 35452 26840 35480 26868
rect 36464 26840 36492 26939
rect 42426 26936 42432 26988
rect 42484 26936 42490 26988
rect 35452 26812 36492 26840
rect 42628 26840 42656 27007
rect 42702 26936 42708 26988
rect 42760 26936 42766 26988
rect 42797 26979 42855 26985
rect 42797 26945 42809 26979
rect 42843 26976 42855 26979
rect 42978 26976 42984 26988
rect 42843 26948 42984 26976
rect 42843 26945 42855 26948
rect 42797 26939 42855 26945
rect 42978 26936 42984 26948
rect 43036 26936 43042 26988
rect 43441 26979 43499 26985
rect 43441 26945 43453 26979
rect 43487 26976 43499 26979
rect 43901 26979 43959 26985
rect 43901 26976 43913 26979
rect 43487 26948 43913 26976
rect 43487 26945 43499 26948
rect 43441 26939 43499 26945
rect 43901 26945 43913 26948
rect 43947 26976 43959 26979
rect 43990 26976 43996 26988
rect 43947 26948 43996 26976
rect 43947 26945 43959 26948
rect 43901 26939 43959 26945
rect 43990 26936 43996 26948
rect 44048 26936 44054 26988
rect 43530 26868 43536 26920
rect 43588 26868 43594 26920
rect 44085 26843 44143 26849
rect 44085 26840 44097 26843
rect 42628 26812 44097 26840
rect 44085 26809 44097 26812
rect 44131 26809 44143 26843
rect 44085 26803 44143 26809
rect 38102 26772 38108 26784
rect 35268 26744 38108 26772
rect 38102 26732 38108 26744
rect 38160 26732 38166 26784
rect 42886 26732 42892 26784
rect 42944 26772 42950 26784
rect 42981 26775 43039 26781
rect 42981 26772 42993 26775
rect 42944 26744 42993 26772
rect 42944 26732 42950 26744
rect 42981 26741 42993 26744
rect 43027 26741 43039 26775
rect 42981 26735 43039 26741
rect 43070 26732 43076 26784
rect 43128 26732 43134 26784
rect 1104 26682 45172 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 45172 26682
rect 1104 26608 45172 26630
rect 11517 26571 11575 26577
rect 11517 26537 11529 26571
rect 11563 26568 11575 26571
rect 12066 26568 12072 26580
rect 11563 26540 12072 26568
rect 11563 26537 11575 26540
rect 11517 26531 11575 26537
rect 12066 26528 12072 26540
rect 12124 26528 12130 26580
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 16301 26571 16359 26577
rect 16301 26568 16313 26571
rect 13136 26540 16313 26568
rect 13136 26528 13142 26540
rect 16301 26537 16313 26540
rect 16347 26537 16359 26571
rect 16301 26531 16359 26537
rect 18046 26528 18052 26580
rect 18104 26528 18110 26580
rect 18414 26528 18420 26580
rect 18472 26568 18478 26580
rect 18509 26571 18567 26577
rect 18509 26568 18521 26571
rect 18472 26540 18521 26568
rect 18472 26528 18478 26540
rect 18509 26537 18521 26540
rect 18555 26537 18567 26571
rect 27430 26568 27436 26580
rect 18509 26531 18567 26537
rect 18616 26540 27436 26568
rect 18064 26500 18092 26528
rect 18616 26500 18644 26540
rect 27430 26528 27436 26540
rect 27488 26528 27494 26580
rect 28810 26528 28816 26580
rect 28868 26528 28874 26580
rect 28994 26528 29000 26580
rect 29052 26568 29058 26580
rect 29549 26571 29607 26577
rect 29549 26568 29561 26571
rect 29052 26540 29561 26568
rect 29052 26528 29058 26540
rect 29549 26537 29561 26540
rect 29595 26537 29607 26571
rect 29549 26531 29607 26537
rect 30006 26528 30012 26580
rect 30064 26528 30070 26580
rect 34698 26528 34704 26580
rect 34756 26568 34762 26580
rect 35069 26571 35127 26577
rect 35069 26568 35081 26571
rect 34756 26540 35081 26568
rect 34756 26528 34762 26540
rect 35069 26537 35081 26540
rect 35115 26537 35127 26571
rect 35069 26531 35127 26537
rect 35342 26528 35348 26580
rect 35400 26528 35406 26580
rect 35713 26571 35771 26577
rect 35713 26537 35725 26571
rect 35759 26568 35771 26571
rect 35802 26568 35808 26580
rect 35759 26540 35808 26568
rect 35759 26537 35771 26540
rect 35713 26531 35771 26537
rect 35802 26528 35808 26540
rect 35860 26528 35866 26580
rect 41509 26571 41567 26577
rect 41509 26568 41521 26571
rect 41156 26540 41521 26568
rect 18064 26472 18644 26500
rect 22925 26503 22983 26509
rect 22925 26469 22937 26503
rect 22971 26500 22983 26503
rect 23014 26500 23020 26512
rect 22971 26472 23020 26500
rect 22971 26469 22983 26472
rect 22925 26463 22983 26469
rect 23014 26460 23020 26472
rect 23072 26460 23078 26512
rect 24213 26503 24271 26509
rect 24213 26469 24225 26503
rect 24259 26469 24271 26503
rect 24213 26463 24271 26469
rect 10965 26435 11023 26441
rect 10965 26401 10977 26435
rect 11011 26432 11023 26435
rect 11238 26432 11244 26444
rect 11011 26404 11244 26432
rect 11011 26401 11023 26404
rect 10965 26395 11023 26401
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 12161 26435 12219 26441
rect 12161 26401 12173 26435
rect 12207 26432 12219 26435
rect 12434 26432 12440 26444
rect 12207 26404 12440 26432
rect 12207 26401 12219 26404
rect 12161 26395 12219 26401
rect 12434 26392 12440 26404
rect 12492 26392 12498 26444
rect 16761 26435 16819 26441
rect 16761 26401 16773 26435
rect 16807 26432 16819 26435
rect 17126 26432 17132 26444
rect 16807 26404 17132 26432
rect 16807 26401 16819 26404
rect 16761 26395 16819 26401
rect 17126 26392 17132 26404
rect 17184 26392 17190 26444
rect 20530 26392 20536 26444
rect 20588 26392 20594 26444
rect 21358 26392 21364 26444
rect 21416 26392 21422 26444
rect 21542 26392 21548 26444
rect 21600 26392 21606 26444
rect 23032 26432 23060 26460
rect 23569 26435 23627 26441
rect 23569 26432 23581 26435
rect 23032 26404 23581 26432
rect 23569 26401 23581 26404
rect 23615 26401 23627 26435
rect 24228 26432 24256 26463
rect 26970 26460 26976 26512
rect 27028 26500 27034 26512
rect 27028 26472 30604 26500
rect 27028 26460 27034 26472
rect 24673 26435 24731 26441
rect 24673 26432 24685 26435
rect 24228 26404 24685 26432
rect 23569 26395 23627 26401
rect 24673 26401 24685 26404
rect 24719 26401 24731 26435
rect 24673 26395 24731 26401
rect 28626 26392 28632 26444
rect 28684 26432 28690 26444
rect 28684 26404 29408 26432
rect 28684 26392 28690 26404
rect 10689 26367 10747 26373
rect 10689 26333 10701 26367
rect 10735 26364 10747 26367
rect 10870 26364 10876 26376
rect 10735 26336 10876 26364
rect 10735 26333 10747 26336
rect 10689 26327 10747 26333
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 11977 26367 12035 26373
rect 11977 26333 11989 26367
rect 12023 26364 12035 26367
rect 15749 26367 15807 26373
rect 12023 26336 15700 26364
rect 12023 26333 12035 26336
rect 11977 26327 12035 26333
rect 10781 26299 10839 26305
rect 10781 26265 10793 26299
rect 10827 26296 10839 26299
rect 11790 26296 11796 26308
rect 10827 26268 11796 26296
rect 10827 26265 10839 26268
rect 10781 26259 10839 26265
rect 11790 26256 11796 26268
rect 11848 26296 11854 26308
rect 11885 26299 11943 26305
rect 11885 26296 11897 26299
rect 11848 26268 11897 26296
rect 11848 26256 11854 26268
rect 11885 26265 11897 26268
rect 11931 26265 11943 26299
rect 11885 26259 11943 26265
rect 15286 26256 15292 26308
rect 15344 26296 15350 26308
rect 15473 26299 15531 26305
rect 15473 26296 15485 26299
rect 15344 26268 15485 26296
rect 15344 26256 15350 26268
rect 15473 26265 15485 26268
rect 15519 26265 15531 26299
rect 15672 26296 15700 26336
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 16298 26364 16304 26376
rect 15795 26336 16304 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 16393 26367 16451 26373
rect 16393 26333 16405 26367
rect 16439 26364 16451 26367
rect 16666 26364 16672 26376
rect 16439 26336 16672 26364
rect 16439 26333 16451 26336
rect 16393 26327 16451 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 18138 26324 18144 26376
rect 18196 26364 18202 26376
rect 19242 26364 19248 26376
rect 18196 26336 19248 26364
rect 18196 26324 18202 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 20438 26324 20444 26376
rect 20496 26324 20502 26376
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 24118 26324 24124 26376
rect 24176 26364 24182 26376
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 24176 26336 24409 26364
rect 24176 26324 24182 26336
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 28994 26324 29000 26376
rect 29052 26324 29058 26376
rect 29089 26367 29147 26373
rect 29089 26333 29101 26367
rect 29135 26333 29147 26367
rect 29089 26327 29147 26333
rect 29181 26367 29239 26373
rect 29181 26333 29193 26367
rect 29227 26333 29239 26367
rect 29181 26327 29239 26333
rect 15672 26268 16988 26296
rect 15473 26259 15531 26265
rect 10226 26188 10232 26240
rect 10284 26228 10290 26240
rect 10321 26231 10379 26237
rect 10321 26228 10333 26231
rect 10284 26200 10333 26228
rect 10284 26188 10290 26200
rect 10321 26197 10333 26200
rect 10367 26197 10379 26231
rect 16960 26228 16988 26268
rect 17034 26256 17040 26308
rect 17092 26256 17098 26308
rect 20254 26296 20260 26308
rect 18340 26268 20260 26296
rect 18340 26228 18368 26268
rect 20254 26256 20260 26268
rect 20312 26256 20318 26308
rect 20349 26299 20407 26305
rect 20349 26265 20361 26299
rect 20395 26296 20407 26299
rect 20809 26299 20867 26305
rect 20809 26296 20821 26299
rect 20395 26268 20821 26296
rect 20395 26265 20407 26268
rect 20349 26259 20407 26265
rect 20809 26265 20821 26268
rect 20855 26265 20867 26299
rect 20809 26259 20867 26265
rect 21634 26256 21640 26308
rect 21692 26296 21698 26308
rect 21790 26299 21848 26305
rect 21790 26296 21802 26299
rect 21692 26268 21802 26296
rect 21692 26256 21698 26268
rect 21790 26265 21802 26268
rect 21836 26265 21848 26299
rect 21790 26259 21848 26265
rect 24670 26256 24676 26308
rect 24728 26296 24734 26308
rect 27706 26296 27712 26308
rect 24728 26268 25162 26296
rect 25976 26268 27712 26296
rect 24728 26256 24734 26268
rect 16960 26200 18368 26228
rect 10321 26191 10379 26197
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 19981 26231 20039 26237
rect 19981 26228 19993 26231
rect 19484 26200 19993 26228
rect 19484 26188 19490 26200
rect 19981 26197 19993 26200
rect 20027 26197 20039 26231
rect 19981 26191 20039 26197
rect 23014 26188 23020 26240
rect 23072 26188 23078 26240
rect 25056 26228 25084 26268
rect 25976 26228 26004 26268
rect 27706 26256 27712 26268
rect 27764 26256 27770 26308
rect 25056 26200 26004 26228
rect 26142 26188 26148 26240
rect 26200 26188 26206 26240
rect 29104 26228 29132 26327
rect 29196 26296 29224 26327
rect 29270 26324 29276 26376
rect 29328 26324 29334 26376
rect 29380 26364 29408 26404
rect 29454 26392 29460 26444
rect 29512 26432 29518 26444
rect 30576 26441 30604 26472
rect 33410 26460 33416 26512
rect 33468 26500 33474 26512
rect 33468 26472 34008 26500
rect 33468 26460 33474 26472
rect 29641 26435 29699 26441
rect 29641 26432 29653 26435
rect 29512 26404 29653 26432
rect 29512 26392 29518 26404
rect 29641 26401 29653 26404
rect 29687 26401 29699 26435
rect 29641 26395 29699 26401
rect 30561 26435 30619 26441
rect 30561 26401 30573 26435
rect 30607 26401 30619 26435
rect 30561 26395 30619 26401
rect 32214 26392 32220 26444
rect 32272 26432 32278 26444
rect 32309 26435 32367 26441
rect 32309 26432 32321 26435
rect 32272 26404 32321 26432
rect 32272 26392 32278 26404
rect 32309 26401 32321 26404
rect 32355 26432 32367 26435
rect 32953 26435 33011 26441
rect 32953 26432 32965 26435
rect 32355 26404 32965 26432
rect 32355 26401 32367 26404
rect 32309 26395 32367 26401
rect 32953 26401 32965 26404
rect 32999 26401 33011 26435
rect 32953 26395 33011 26401
rect 33134 26392 33140 26444
rect 33192 26432 33198 26444
rect 33980 26441 34008 26472
rect 33781 26435 33839 26441
rect 33781 26432 33793 26435
rect 33192 26404 33793 26432
rect 33192 26392 33198 26404
rect 33781 26401 33793 26404
rect 33827 26401 33839 26435
rect 33781 26395 33839 26401
rect 33965 26435 34023 26441
rect 33965 26401 33977 26435
rect 34011 26401 34023 26435
rect 33965 26395 34023 26401
rect 34425 26435 34483 26441
rect 34425 26401 34437 26435
rect 34471 26432 34483 26435
rect 34471 26404 34928 26432
rect 34471 26401 34483 26404
rect 34425 26395 34483 26401
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29380 26336 29837 26364
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 33318 26324 33324 26376
rect 33376 26364 33382 26376
rect 33689 26367 33747 26373
rect 33689 26364 33701 26367
rect 33376 26336 33701 26364
rect 33376 26324 33382 26336
rect 33689 26333 33701 26336
rect 33735 26333 33747 26367
rect 33689 26327 33747 26333
rect 34057 26367 34115 26373
rect 34057 26333 34069 26367
rect 34103 26333 34115 26367
rect 34517 26367 34575 26373
rect 34517 26366 34529 26367
rect 34057 26327 34115 26333
rect 34440 26338 34529 26366
rect 29546 26296 29552 26308
rect 29196 26268 29552 26296
rect 29546 26256 29552 26268
rect 29604 26256 29610 26308
rect 30834 26256 30840 26308
rect 30892 26256 30898 26308
rect 31846 26256 31852 26308
rect 31904 26256 31910 26308
rect 34072 26296 34100 26327
rect 33612 26268 34100 26296
rect 34440 26296 34468 26338
rect 34517 26333 34529 26338
rect 34563 26333 34575 26367
rect 34517 26327 34575 26333
rect 34606 26324 34612 26376
rect 34664 26364 34670 26376
rect 34900 26373 34928 26404
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34664 26336 34713 26364
rect 34664 26324 34670 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26333 34943 26367
rect 35360 26364 35388 26528
rect 39209 26435 39267 26441
rect 39209 26401 39221 26435
rect 39255 26432 39267 26435
rect 39390 26432 39396 26444
rect 39255 26404 39396 26432
rect 39255 26401 39267 26404
rect 39209 26395 39267 26401
rect 39390 26392 39396 26404
rect 39448 26432 39454 26444
rect 40129 26435 40187 26441
rect 40129 26432 40141 26435
rect 39448 26404 40141 26432
rect 39448 26392 39454 26404
rect 40129 26401 40141 26404
rect 40175 26401 40187 26435
rect 40129 26395 40187 26401
rect 40494 26392 40500 26444
rect 40552 26432 40558 26444
rect 40954 26432 40960 26444
rect 40552 26404 40960 26432
rect 40552 26392 40558 26404
rect 40954 26392 40960 26404
rect 41012 26432 41018 26444
rect 41156 26441 41184 26540
rect 41509 26537 41521 26540
rect 41555 26537 41567 26571
rect 41509 26531 41567 26537
rect 42610 26528 42616 26580
rect 42668 26528 42674 26580
rect 42978 26528 42984 26580
rect 43036 26528 43042 26580
rect 43990 26528 43996 26580
rect 44048 26568 44054 26580
rect 44729 26571 44787 26577
rect 44729 26568 44741 26571
rect 44048 26540 44741 26568
rect 44048 26528 44054 26540
rect 44729 26537 44741 26540
rect 44775 26537 44787 26571
rect 44729 26531 44787 26537
rect 42153 26503 42211 26509
rect 42153 26500 42165 26503
rect 41616 26472 42165 26500
rect 41049 26435 41107 26441
rect 41049 26432 41061 26435
rect 41012 26404 41061 26432
rect 41012 26392 41018 26404
rect 41049 26401 41061 26404
rect 41095 26401 41107 26435
rect 41049 26395 41107 26401
rect 41141 26435 41199 26441
rect 41141 26401 41153 26435
rect 41187 26401 41199 26435
rect 41616 26432 41644 26472
rect 42153 26469 42165 26472
rect 42199 26469 42211 26503
rect 42153 26463 42211 26469
rect 42521 26435 42579 26441
rect 42521 26432 42533 26435
rect 41141 26395 41199 26401
rect 41248 26404 41644 26432
rect 41892 26404 42533 26432
rect 35529 26367 35587 26373
rect 35529 26364 35541 26367
rect 35360 26336 35541 26364
rect 34885 26327 34943 26333
rect 35529 26333 35541 26336
rect 35575 26333 35587 26367
rect 35529 26327 35587 26333
rect 36906 26324 36912 26376
rect 36964 26324 36970 26376
rect 37274 26324 37280 26376
rect 37332 26364 37338 26376
rect 37461 26367 37519 26373
rect 37461 26364 37473 26367
rect 37332 26336 37473 26364
rect 37332 26324 37338 26336
rect 37461 26333 37473 26336
rect 37507 26333 37519 26367
rect 37461 26327 37519 26333
rect 39301 26367 39359 26373
rect 39301 26333 39313 26367
rect 39347 26364 39359 26367
rect 39853 26367 39911 26373
rect 39853 26364 39865 26367
rect 39347 26336 39865 26364
rect 39347 26333 39359 26336
rect 39301 26327 39359 26333
rect 39853 26333 39865 26336
rect 39899 26333 39911 26367
rect 39853 26327 39911 26333
rect 39942 26324 39948 26376
rect 40000 26324 40006 26376
rect 40037 26367 40095 26373
rect 40037 26333 40049 26367
rect 40083 26333 40095 26367
rect 40037 26327 40095 26333
rect 34440 26268 34836 26296
rect 33612 26240 33640 26268
rect 34808 26240 34836 26268
rect 35342 26256 35348 26308
rect 35400 26256 35406 26308
rect 36924 26296 36952 26324
rect 36924 26268 37688 26296
rect 29454 26228 29460 26240
rect 29104 26200 29460 26228
rect 29454 26188 29460 26200
rect 29512 26188 29518 26240
rect 32122 26188 32128 26240
rect 32180 26228 32186 26240
rect 32401 26231 32459 26237
rect 32401 26228 32413 26231
rect 32180 26200 32413 26228
rect 32180 26188 32186 26200
rect 32401 26197 32413 26200
rect 32447 26197 32459 26231
rect 32401 26191 32459 26197
rect 33594 26188 33600 26240
rect 33652 26188 33658 26240
rect 33962 26188 33968 26240
rect 34020 26188 34026 26240
rect 34146 26188 34152 26240
rect 34204 26188 34210 26240
rect 34790 26188 34796 26240
rect 34848 26188 34854 26240
rect 37660 26228 37688 26268
rect 37734 26256 37740 26308
rect 37792 26256 37798 26308
rect 37844 26268 38226 26296
rect 37844 26228 37872 26268
rect 37660 26200 37872 26228
rect 38120 26228 38148 26268
rect 39482 26256 39488 26308
rect 39540 26256 39546 26308
rect 39574 26256 39580 26308
rect 39632 26256 39638 26308
rect 39669 26299 39727 26305
rect 39669 26265 39681 26299
rect 39715 26296 39727 26299
rect 39960 26296 39988 26324
rect 39715 26268 39988 26296
rect 39715 26265 39727 26268
rect 39669 26259 39727 26265
rect 38746 26228 38752 26240
rect 38120 26200 38752 26228
rect 38746 26188 38752 26200
rect 38804 26188 38810 26240
rect 39592 26228 39620 26256
rect 40052 26228 40080 26327
rect 40218 26324 40224 26376
rect 40276 26324 40282 26376
rect 40405 26367 40463 26373
rect 40405 26333 40417 26367
rect 40451 26364 40463 26367
rect 40681 26367 40739 26373
rect 40681 26364 40693 26367
rect 40451 26336 40693 26364
rect 40451 26333 40463 26336
rect 40405 26327 40463 26333
rect 40681 26333 40693 26336
rect 40727 26333 40739 26367
rect 40681 26327 40739 26333
rect 40862 26324 40868 26376
rect 40920 26324 40926 26376
rect 41248 26373 41276 26404
rect 41233 26367 41291 26373
rect 41233 26333 41245 26367
rect 41279 26333 41291 26367
rect 41233 26327 41291 26333
rect 41414 26324 41420 26376
rect 41472 26324 41478 26376
rect 41506 26324 41512 26376
rect 41564 26364 41570 26376
rect 41892 26373 41920 26404
rect 42521 26401 42533 26404
rect 42567 26432 42579 26435
rect 42628 26432 42656 26528
rect 42996 26500 43024 26528
rect 42567 26404 42656 26432
rect 42720 26472 43024 26500
rect 42567 26401 42579 26404
rect 42521 26395 42579 26401
rect 42720 26373 42748 26472
rect 42794 26392 42800 26444
rect 42852 26432 42858 26444
rect 42981 26435 43039 26441
rect 42981 26432 42993 26435
rect 42852 26404 42993 26432
rect 42852 26392 42858 26404
rect 42981 26401 42993 26404
rect 43027 26401 43039 26435
rect 42981 26395 43039 26401
rect 41693 26367 41751 26373
rect 41693 26364 41705 26367
rect 41564 26336 41705 26364
rect 41564 26324 41570 26336
rect 41693 26333 41705 26336
rect 41739 26333 41751 26367
rect 41693 26327 41751 26333
rect 41877 26367 41935 26373
rect 41877 26333 41889 26367
rect 41923 26333 41935 26367
rect 41877 26327 41935 26333
rect 42061 26367 42119 26373
rect 42061 26333 42073 26367
rect 42107 26364 42119 26367
rect 42337 26367 42395 26373
rect 42337 26364 42349 26367
rect 42107 26336 42349 26364
rect 42107 26333 42119 26336
rect 42061 26327 42119 26333
rect 42337 26333 42349 26336
rect 42383 26364 42395 26367
rect 42613 26367 42671 26373
rect 42383 26336 42564 26364
rect 42383 26333 42395 26336
rect 42337 26327 42395 26333
rect 42536 26308 42564 26336
rect 42613 26333 42625 26367
rect 42659 26333 42671 26367
rect 42613 26327 42671 26333
rect 42705 26367 42763 26373
rect 42705 26333 42717 26367
rect 42751 26333 42763 26367
rect 42705 26327 42763 26333
rect 40586 26256 40592 26308
rect 40644 26256 40650 26308
rect 41782 26296 41788 26308
rect 41386 26268 41788 26296
rect 39592 26200 40080 26228
rect 41138 26188 41144 26240
rect 41196 26228 41202 26240
rect 41386 26228 41414 26268
rect 41782 26256 41788 26268
rect 41840 26256 41846 26308
rect 42518 26256 42524 26308
rect 42576 26256 42582 26308
rect 41196 26200 41414 26228
rect 42628 26228 42656 26327
rect 42886 26324 42892 26376
rect 42944 26324 42950 26376
rect 43254 26256 43260 26308
rect 43312 26256 43318 26308
rect 43714 26256 43720 26308
rect 43772 26256 43778 26308
rect 42702 26228 42708 26240
rect 42628 26200 42708 26228
rect 41196 26188 41202 26200
rect 42702 26188 42708 26200
rect 42760 26228 42766 26240
rect 43346 26228 43352 26240
rect 42760 26200 43352 26228
rect 42760 26188 42766 26200
rect 43346 26188 43352 26200
rect 43404 26188 43410 26240
rect 1104 26138 45172 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 45172 26138
rect 1104 26064 45172 26086
rect 7098 25984 7104 26036
rect 7156 25984 7162 26036
rect 8128 25996 9812 26024
rect 7116 25956 7144 25984
rect 8128 25956 8156 25996
rect 9784 25956 9812 25996
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12492 25996 13768 26024
rect 12492 25984 12498 25996
rect 9950 25956 9956 25968
rect 7116 25928 8234 25956
rect 9784 25928 9956 25956
rect 9950 25916 9956 25928
rect 10008 25956 10014 25968
rect 10008 25928 10166 25956
rect 10008 25916 10014 25928
rect 11606 25916 11612 25968
rect 11664 25956 11670 25968
rect 13740 25956 13768 25996
rect 17034 25984 17040 26036
rect 17092 26024 17098 26036
rect 17221 26027 17279 26033
rect 17221 26024 17233 26027
rect 17092 25996 17233 26024
rect 17092 25984 17098 25996
rect 17221 25993 17233 25996
rect 17267 25993 17279 26027
rect 17221 25987 17279 25993
rect 17589 26027 17647 26033
rect 17589 25993 17601 26027
rect 17635 25993 17647 26027
rect 17589 25987 17647 25993
rect 17957 26027 18015 26033
rect 17957 25993 17969 26027
rect 18003 26024 18015 26027
rect 18414 26024 18420 26036
rect 18003 25996 18420 26024
rect 18003 25993 18015 25996
rect 17957 25987 18015 25993
rect 11664 25928 13216 25956
rect 13740 25928 13952 25956
rect 11664 25916 11670 25928
rect 12986 25848 12992 25900
rect 13044 25897 13050 25900
rect 13044 25851 13056 25897
rect 13044 25848 13050 25851
rect 7469 25823 7527 25829
rect 7469 25789 7481 25823
rect 7515 25789 7527 25823
rect 7469 25783 7527 25789
rect 7484 25684 7512 25783
rect 7742 25780 7748 25832
rect 7800 25780 7806 25832
rect 9401 25823 9459 25829
rect 9401 25789 9413 25823
rect 9447 25789 9459 25823
rect 9401 25783 9459 25789
rect 9416 25752 9444 25783
rect 9674 25780 9680 25832
rect 9732 25780 9738 25832
rect 10870 25780 10876 25832
rect 10928 25820 10934 25832
rect 11149 25823 11207 25829
rect 11149 25820 11161 25823
rect 10928 25792 11161 25820
rect 10928 25780 10934 25792
rect 11149 25789 11161 25792
rect 11195 25789 11207 25823
rect 13188 25820 13216 25928
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25888 13323 25891
rect 13446 25888 13452 25900
rect 13311 25860 13452 25888
rect 13311 25857 13323 25860
rect 13265 25851 13323 25857
rect 13446 25848 13452 25860
rect 13504 25848 13510 25900
rect 13725 25891 13783 25897
rect 13725 25857 13737 25891
rect 13771 25857 13783 25891
rect 13725 25851 13783 25857
rect 13740 25820 13768 25851
rect 13924 25829 13952 25928
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 16758 25888 16764 25900
rect 16347 25860 16764 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 16758 25848 16764 25860
rect 16816 25848 16822 25900
rect 17405 25891 17463 25897
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 17604 25888 17632 25987
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 19334 25984 19340 26036
rect 19392 25984 19398 26036
rect 19426 25984 19432 26036
rect 19484 25984 19490 26036
rect 19705 26027 19763 26033
rect 19705 25993 19717 26027
rect 19751 25993 19763 26027
rect 19705 25987 19763 25993
rect 21177 26027 21235 26033
rect 21177 25993 21189 26027
rect 21223 26024 21235 26027
rect 21358 26024 21364 26036
rect 21223 25996 21364 26024
rect 21223 25993 21235 25996
rect 21177 25987 21235 25993
rect 19352 25956 19380 25984
rect 19168 25928 19380 25956
rect 17451 25860 17632 25888
rect 18049 25891 18107 25897
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 18049 25857 18061 25891
rect 18095 25888 18107 25891
rect 18690 25888 18696 25900
rect 18095 25860 18696 25888
rect 18095 25857 18107 25860
rect 18049 25851 18107 25857
rect 18690 25848 18696 25860
rect 18748 25848 18754 25900
rect 13188 25792 13768 25820
rect 13817 25823 13875 25829
rect 11149 25783 11207 25789
rect 13817 25789 13829 25823
rect 13863 25789 13875 25823
rect 13817 25783 13875 25789
rect 13909 25823 13967 25829
rect 13909 25789 13921 25823
rect 13955 25789 13967 25823
rect 13909 25783 13967 25789
rect 16025 25823 16083 25829
rect 16025 25789 16037 25823
rect 16071 25820 16083 25823
rect 16206 25820 16212 25832
rect 16071 25792 16212 25820
rect 16071 25789 16083 25792
rect 16025 25783 16083 25789
rect 8772 25724 9444 25752
rect 13832 25752 13860 25783
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 18233 25823 18291 25829
rect 18233 25789 18245 25823
rect 18279 25820 18291 25823
rect 18598 25820 18604 25832
rect 18279 25792 18604 25820
rect 18279 25789 18291 25792
rect 18233 25783 18291 25789
rect 18598 25780 18604 25792
rect 18656 25820 18662 25832
rect 19168 25820 19196 25928
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25888 19303 25891
rect 19334 25888 19340 25900
rect 19291 25860 19340 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 19444 25888 19472 25984
rect 19720 25956 19748 25987
rect 21358 25984 21364 25996
rect 21416 25984 21422 26036
rect 21634 25984 21640 26036
rect 21692 25984 21698 26036
rect 21821 26027 21879 26033
rect 21821 25993 21833 26027
rect 21867 25993 21879 26027
rect 21821 25987 21879 25993
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 23014 26024 23020 26036
rect 22235 25996 23020 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 20064 25959 20122 25965
rect 20064 25956 20076 25959
rect 19720 25928 20076 25956
rect 20064 25925 20076 25928
rect 20110 25925 20122 25959
rect 20064 25919 20122 25925
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19444 25860 19533 25888
rect 19521 25857 19533 25860
rect 19567 25857 19579 25891
rect 19521 25851 19579 25857
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 21836 25888 21864 25987
rect 23014 25984 23020 25996
rect 23072 25984 23078 26036
rect 24026 25984 24032 26036
rect 24084 26024 24090 26036
rect 24213 26027 24271 26033
rect 24213 26024 24225 26027
rect 24084 25996 24225 26024
rect 24084 25984 24090 25996
rect 24213 25993 24225 25996
rect 24259 25993 24271 26027
rect 24213 25987 24271 25993
rect 24581 26027 24639 26033
rect 24581 25993 24593 26027
rect 24627 26024 24639 26027
rect 26142 26024 26148 26036
rect 24627 25996 26148 26024
rect 24627 25993 24639 25996
rect 24581 25987 24639 25993
rect 26142 25984 26148 25996
rect 26200 25984 26206 26036
rect 26789 26027 26847 26033
rect 26789 25993 26801 26027
rect 26835 25993 26847 26027
rect 26789 25987 26847 25993
rect 26804 25956 26832 25987
rect 29638 25984 29644 26036
rect 29696 25984 29702 26036
rect 30834 25984 30840 26036
rect 30892 26024 30898 26036
rect 31297 26027 31355 26033
rect 31297 26024 31309 26027
rect 30892 25996 31309 26024
rect 30892 25984 30898 25996
rect 31297 25993 31309 25996
rect 31343 25993 31355 26027
rect 32493 26027 32551 26033
rect 31297 25987 31355 25993
rect 31864 25996 32444 26024
rect 27249 25959 27307 25965
rect 27249 25956 27261 25959
rect 26804 25928 27261 25956
rect 27249 25925 27261 25928
rect 27295 25925 27307 25959
rect 27249 25919 27307 25925
rect 27706 25916 27712 25968
rect 27764 25916 27770 25968
rect 31864 25965 31892 25996
rect 31849 25959 31907 25965
rect 31849 25925 31861 25959
rect 31895 25925 31907 25959
rect 31849 25919 31907 25925
rect 31941 25959 31999 25965
rect 31941 25925 31953 25959
rect 31987 25956 31999 25959
rect 32122 25956 32128 25968
rect 31987 25928 32128 25956
rect 31987 25925 31999 25928
rect 31941 25919 31999 25925
rect 32122 25916 32128 25928
rect 32180 25916 32186 25968
rect 32416 25956 32444 25996
rect 32493 25993 32505 26027
rect 32539 26024 32551 26027
rect 33134 26024 33140 26036
rect 32539 25996 33140 26024
rect 32539 25993 32551 25996
rect 32493 25987 32551 25993
rect 33134 25984 33140 25996
rect 33192 25984 33198 26036
rect 37734 25984 37740 26036
rect 37792 26024 37798 26036
rect 37829 26027 37887 26033
rect 37829 26024 37841 26027
rect 37792 25996 37841 26024
rect 37792 25984 37798 25996
rect 37829 25993 37841 25996
rect 37875 25993 37887 26027
rect 37829 25987 37887 25993
rect 39390 25984 39396 26036
rect 39448 25984 39454 26036
rect 39574 25984 39580 26036
rect 39632 25984 39638 26036
rect 39942 25984 39948 26036
rect 40000 25984 40006 26036
rect 40218 25984 40224 26036
rect 40276 25984 40282 26036
rect 40957 26027 41015 26033
rect 40957 25993 40969 26027
rect 41003 26024 41015 26027
rect 41414 26024 41420 26036
rect 41003 25996 41420 26024
rect 41003 25993 41015 25996
rect 40957 25987 41015 25993
rect 41414 25984 41420 25996
rect 41472 25984 41478 26036
rect 42426 25984 42432 26036
rect 42484 25984 42490 26036
rect 43162 26024 43168 26036
rect 42628 25996 43168 26024
rect 32416 25928 33088 25956
rect 21499 25860 21864 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 23566 25848 23572 25900
rect 23624 25848 23630 25900
rect 26602 25848 26608 25900
rect 26660 25848 26666 25900
rect 29270 25848 29276 25900
rect 29328 25888 29334 25900
rect 29457 25891 29515 25897
rect 29457 25888 29469 25891
rect 29328 25860 29469 25888
rect 29328 25848 29334 25860
rect 29457 25857 29469 25860
rect 29503 25857 29515 25891
rect 29457 25851 29515 25857
rect 31570 25848 31576 25900
rect 31628 25848 31634 25900
rect 32214 25848 32220 25900
rect 32272 25848 32278 25900
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 18656 25792 19196 25820
rect 18656 25780 18662 25792
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19797 25823 19855 25829
rect 19797 25820 19809 25823
rect 19484 25792 19809 25820
rect 19484 25780 19490 25792
rect 19797 25789 19809 25792
rect 19843 25789 19855 25823
rect 19797 25783 19855 25789
rect 22278 25780 22284 25832
rect 22336 25780 22342 25832
rect 22462 25780 22468 25832
rect 22520 25780 22526 25832
rect 22830 25780 22836 25832
rect 22888 25780 22894 25832
rect 23477 25823 23535 25829
rect 23477 25789 23489 25823
rect 23523 25820 23535 25823
rect 24673 25823 24731 25829
rect 24673 25820 24685 25823
rect 23523 25792 24685 25820
rect 23523 25789 23535 25792
rect 23477 25783 23535 25789
rect 24673 25789 24685 25792
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 24762 25780 24768 25832
rect 24820 25780 24826 25832
rect 26970 25780 26976 25832
rect 27028 25780 27034 25832
rect 29181 25823 29239 25829
rect 29181 25789 29193 25823
rect 29227 25820 29239 25823
rect 29227 25792 29500 25820
rect 29227 25789 29239 25792
rect 29181 25783 29239 25789
rect 29472 25764 29500 25792
rect 31478 25780 31484 25832
rect 31536 25780 31542 25832
rect 32324 25820 32352 25851
rect 32490 25848 32496 25900
rect 32548 25888 32554 25900
rect 32585 25891 32643 25897
rect 32585 25888 32597 25891
rect 32548 25860 32597 25888
rect 32548 25848 32554 25860
rect 32585 25857 32597 25860
rect 32631 25857 32643 25891
rect 32585 25851 32643 25857
rect 32674 25848 32680 25900
rect 32732 25888 32738 25900
rect 32953 25891 33011 25897
rect 32953 25888 32965 25891
rect 32732 25860 32965 25888
rect 32732 25848 32738 25860
rect 32953 25857 32965 25860
rect 32999 25857 33011 25891
rect 32953 25851 33011 25857
rect 33060 25832 33088 25928
rect 33704 25928 34192 25956
rect 33704 25897 33732 25928
rect 34164 25900 34192 25928
rect 33689 25891 33747 25897
rect 33689 25857 33701 25891
rect 33735 25857 33747 25891
rect 33689 25851 33747 25857
rect 33962 25848 33968 25900
rect 34020 25848 34026 25900
rect 34146 25848 34152 25900
rect 34204 25848 34210 25900
rect 39408 25897 39436 25984
rect 39301 25891 39359 25897
rect 39301 25857 39313 25891
rect 39347 25888 39359 25891
rect 39393 25891 39451 25897
rect 39393 25888 39405 25891
rect 39347 25860 39405 25888
rect 39347 25857 39359 25860
rect 39301 25851 39359 25857
rect 39393 25857 39405 25860
rect 39439 25857 39451 25891
rect 39393 25851 39451 25857
rect 39482 25848 39488 25900
rect 39540 25848 39546 25900
rect 39592 25897 39620 25984
rect 39853 25959 39911 25965
rect 39853 25925 39865 25959
rect 39899 25956 39911 25959
rect 39960 25956 39988 25984
rect 39899 25928 39988 25956
rect 39899 25925 39911 25928
rect 39853 25919 39911 25925
rect 40862 25916 40868 25968
rect 40920 25916 40926 25968
rect 41138 25916 41144 25968
rect 41196 25916 41202 25968
rect 41325 25959 41383 25965
rect 41325 25925 41337 25959
rect 41371 25956 41383 25959
rect 41506 25956 41512 25968
rect 41371 25928 41512 25956
rect 41371 25925 41383 25928
rect 41325 25919 41383 25925
rect 41506 25916 41512 25928
rect 41564 25916 41570 25968
rect 39577 25891 39635 25897
rect 39577 25857 39589 25891
rect 39623 25857 39635 25891
rect 39577 25851 39635 25857
rect 39669 25891 39727 25897
rect 39669 25857 39681 25891
rect 39715 25857 39727 25891
rect 39669 25851 39727 25857
rect 39945 25891 40003 25897
rect 39945 25857 39957 25891
rect 39991 25857 40003 25891
rect 39945 25851 40003 25857
rect 40037 25891 40095 25897
rect 40037 25857 40049 25891
rect 40083 25888 40095 25891
rect 40494 25888 40500 25900
rect 40083 25860 40500 25888
rect 40083 25857 40095 25860
rect 40037 25851 40095 25857
rect 32140 25792 32352 25820
rect 32140 25764 32168 25792
rect 33042 25780 33048 25832
rect 33100 25780 33106 25832
rect 34057 25823 34115 25829
rect 34057 25789 34069 25823
rect 34103 25820 34115 25823
rect 35342 25820 35348 25832
rect 34103 25792 35348 25820
rect 34103 25789 34115 25792
rect 34057 25783 34115 25789
rect 35342 25780 35348 25792
rect 35400 25780 35406 25832
rect 38378 25780 38384 25832
rect 38436 25780 38442 25832
rect 39500 25820 39528 25848
rect 39684 25820 39712 25851
rect 39500 25792 39712 25820
rect 39960 25820 39988 25851
rect 40494 25848 40500 25860
rect 40552 25848 40558 25900
rect 40402 25820 40408 25832
rect 39960 25792 40408 25820
rect 40402 25780 40408 25792
rect 40460 25820 40466 25832
rect 40880 25820 40908 25916
rect 42628 25897 42656 25996
rect 43162 25984 43168 25996
rect 43220 25984 43226 26036
rect 43254 25984 43260 26036
rect 43312 25984 43318 26036
rect 42904 25928 44220 25956
rect 42904 25897 42932 25928
rect 44192 25900 44220 25928
rect 42613 25891 42671 25897
rect 42613 25857 42625 25891
rect 42659 25857 42671 25891
rect 42613 25851 42671 25857
rect 42705 25891 42763 25897
rect 42705 25857 42717 25891
rect 42751 25857 42763 25891
rect 42705 25851 42763 25857
rect 42889 25891 42947 25897
rect 42889 25857 42901 25891
rect 42935 25857 42947 25891
rect 42889 25851 42947 25857
rect 40460 25792 40908 25820
rect 40460 25780 40466 25792
rect 42058 25780 42064 25832
rect 42116 25820 42122 25832
rect 42720 25820 42748 25851
rect 42978 25848 42984 25900
rect 43036 25848 43042 25900
rect 43070 25848 43076 25900
rect 43128 25888 43134 25900
rect 43809 25891 43867 25897
rect 43809 25888 43821 25891
rect 43128 25860 43821 25888
rect 43128 25848 43134 25860
rect 43809 25857 43821 25860
rect 43855 25857 43867 25891
rect 43809 25851 43867 25857
rect 44174 25848 44180 25900
rect 44232 25848 44238 25900
rect 42116 25792 43116 25820
rect 42116 25780 42122 25792
rect 17954 25752 17960 25764
rect 13832 25724 17960 25752
rect 8202 25684 8208 25696
rect 7484 25656 8208 25684
rect 8202 25644 8208 25656
rect 8260 25684 8266 25696
rect 8772 25684 8800 25724
rect 8260 25656 8800 25684
rect 9217 25687 9275 25693
rect 8260 25644 8266 25656
rect 9217 25653 9229 25687
rect 9263 25684 9275 25687
rect 9306 25684 9312 25696
rect 9263 25656 9312 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 9306 25644 9312 25656
rect 9364 25644 9370 25696
rect 9416 25684 9444 25724
rect 17954 25712 17960 25724
rect 18012 25712 18018 25764
rect 29454 25712 29460 25764
rect 29512 25712 29518 25764
rect 32122 25712 32128 25764
rect 32180 25712 32186 25764
rect 42518 25712 42524 25764
rect 42576 25752 42582 25764
rect 42886 25752 42892 25764
rect 42576 25724 42892 25752
rect 42576 25712 42582 25724
rect 42886 25712 42892 25724
rect 42944 25712 42950 25764
rect 43088 25752 43116 25792
rect 43346 25780 43352 25832
rect 43404 25820 43410 25832
rect 44545 25823 44603 25829
rect 44545 25820 44557 25823
rect 43404 25792 44557 25820
rect 43404 25780 43410 25792
rect 44545 25789 44557 25792
rect 44591 25789 44603 25823
rect 44545 25783 44603 25789
rect 43162 25752 43168 25764
rect 43088 25724 43168 25752
rect 43162 25712 43168 25724
rect 43220 25752 43226 25764
rect 43898 25752 43904 25764
rect 43220 25724 43904 25752
rect 43220 25712 43226 25724
rect 43898 25712 43904 25724
rect 43956 25712 43962 25764
rect 10318 25684 10324 25696
rect 9416 25656 10324 25684
rect 10318 25644 10324 25656
rect 10376 25644 10382 25696
rect 11882 25644 11888 25696
rect 11940 25644 11946 25696
rect 13354 25644 13360 25696
rect 13412 25644 13418 25696
rect 15194 25644 15200 25696
rect 15252 25684 15258 25696
rect 15381 25687 15439 25693
rect 15381 25684 15393 25687
rect 15252 25656 15393 25684
rect 15252 25644 15258 25656
rect 15381 25653 15393 25656
rect 15427 25653 15439 25687
rect 15381 25647 15439 25653
rect 16114 25644 16120 25696
rect 16172 25644 16178 25696
rect 19429 25687 19487 25693
rect 19429 25653 19441 25687
rect 19475 25684 19487 25687
rect 19518 25684 19524 25696
rect 19475 25656 19524 25684
rect 19475 25653 19487 25656
rect 19429 25647 19487 25653
rect 19518 25644 19524 25656
rect 19576 25644 19582 25696
rect 23750 25644 23756 25696
rect 23808 25644 23814 25696
rect 28721 25687 28779 25693
rect 28721 25653 28733 25687
rect 28767 25684 28779 25687
rect 28994 25684 29000 25696
rect 28767 25656 29000 25684
rect 28767 25653 28779 25656
rect 28721 25647 28779 25653
rect 28994 25644 29000 25656
rect 29052 25644 29058 25696
rect 29273 25687 29331 25693
rect 29273 25653 29285 25687
rect 29319 25684 29331 25687
rect 29546 25684 29552 25696
rect 29319 25656 29552 25684
rect 29319 25653 29331 25656
rect 29273 25647 29331 25653
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 29730 25644 29736 25696
rect 29788 25684 29794 25696
rect 32398 25684 32404 25696
rect 29788 25656 32404 25684
rect 29788 25644 29794 25656
rect 32398 25644 32404 25656
rect 32456 25644 32462 25696
rect 38654 25644 38660 25696
rect 38712 25644 38718 25696
rect 39022 25644 39028 25696
rect 39080 25684 39086 25696
rect 39485 25687 39543 25693
rect 39485 25684 39497 25687
rect 39080 25656 39497 25684
rect 39080 25644 39086 25656
rect 39485 25653 39497 25656
rect 39531 25653 39543 25687
rect 39485 25647 39543 25653
rect 42794 25644 42800 25696
rect 42852 25684 42858 25696
rect 43993 25687 44051 25693
rect 43993 25684 44005 25687
rect 42852 25656 44005 25684
rect 42852 25644 42858 25656
rect 43993 25653 44005 25656
rect 44039 25653 44051 25687
rect 43993 25647 44051 25653
rect 1104 25594 45172 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 45172 25594
rect 1104 25520 45172 25542
rect 7742 25440 7748 25492
rect 7800 25480 7806 25492
rect 8205 25483 8263 25489
rect 8205 25480 8217 25483
rect 7800 25452 8217 25480
rect 7800 25440 7806 25452
rect 8205 25449 8217 25452
rect 8251 25449 8263 25483
rect 8205 25443 8263 25449
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 9861 25483 9919 25489
rect 9861 25480 9873 25483
rect 9732 25452 9873 25480
rect 9732 25440 9738 25452
rect 9861 25449 9873 25452
rect 9907 25449 9919 25483
rect 11238 25480 11244 25492
rect 9861 25443 9919 25449
rect 10152 25452 11244 25480
rect 9585 25347 9643 25353
rect 9585 25313 9597 25347
rect 9631 25344 9643 25347
rect 10152 25344 10180 25452
rect 11238 25440 11244 25452
rect 11296 25440 11302 25492
rect 11790 25440 11796 25492
rect 11848 25480 11854 25492
rect 11885 25483 11943 25489
rect 11885 25480 11897 25483
rect 11848 25452 11897 25480
rect 11848 25440 11854 25452
rect 11885 25449 11897 25452
rect 11931 25449 11943 25483
rect 11885 25443 11943 25449
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 12986 25480 12992 25492
rect 12851 25452 12992 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 12986 25440 12992 25452
rect 13044 25440 13050 25492
rect 13354 25440 13360 25492
rect 13412 25440 13418 25492
rect 15286 25440 15292 25492
rect 15344 25440 15350 25492
rect 15552 25483 15610 25489
rect 15552 25449 15564 25483
rect 15598 25480 15610 25483
rect 16114 25480 16120 25492
rect 15598 25452 16120 25480
rect 15598 25449 15610 25452
rect 15552 25443 15610 25449
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 16666 25440 16672 25492
rect 16724 25480 16730 25492
rect 17034 25480 17040 25492
rect 16724 25452 17040 25480
rect 16724 25440 16730 25452
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 18322 25440 18328 25492
rect 18380 25480 18386 25492
rect 19061 25483 19119 25489
rect 19061 25480 19073 25483
rect 18380 25452 19073 25480
rect 18380 25440 18386 25452
rect 19061 25449 19073 25452
rect 19107 25449 19119 25483
rect 19061 25443 19119 25449
rect 19518 25440 19524 25492
rect 19576 25440 19582 25492
rect 20254 25440 20260 25492
rect 20312 25480 20318 25492
rect 20901 25483 20959 25489
rect 20901 25480 20913 25483
rect 20312 25452 20913 25480
rect 20312 25440 20318 25452
rect 20901 25449 20913 25452
rect 20947 25480 20959 25483
rect 22830 25480 22836 25492
rect 20947 25452 22836 25480
rect 20947 25449 20959 25452
rect 20901 25443 20959 25449
rect 22830 25440 22836 25452
rect 22888 25440 22894 25492
rect 26602 25440 26608 25492
rect 26660 25480 26666 25492
rect 26697 25483 26755 25489
rect 26697 25480 26709 25483
rect 26660 25452 26709 25480
rect 26660 25440 26666 25452
rect 26697 25449 26709 25452
rect 26743 25449 26755 25483
rect 26697 25443 26755 25449
rect 29546 25440 29552 25492
rect 29604 25440 29610 25492
rect 31478 25440 31484 25492
rect 31536 25440 31542 25492
rect 31570 25440 31576 25492
rect 31628 25480 31634 25492
rect 31757 25483 31815 25489
rect 31757 25480 31769 25483
rect 31628 25452 31769 25480
rect 31628 25440 31634 25452
rect 31757 25449 31769 25452
rect 31803 25449 31815 25483
rect 31757 25443 31815 25449
rect 31938 25440 31944 25492
rect 31996 25480 32002 25492
rect 32674 25480 32680 25492
rect 31996 25452 32680 25480
rect 31996 25440 32002 25452
rect 32674 25440 32680 25452
rect 32732 25440 32738 25492
rect 32861 25483 32919 25489
rect 32861 25449 32873 25483
rect 32907 25480 32919 25483
rect 33410 25480 33416 25492
rect 32907 25452 33416 25480
rect 32907 25449 32919 25452
rect 32861 25443 32919 25449
rect 33410 25440 33416 25452
rect 33468 25440 33474 25492
rect 36262 25480 36268 25492
rect 33796 25452 36268 25480
rect 10226 25372 10232 25424
rect 10284 25372 10290 25424
rect 11701 25415 11759 25421
rect 11701 25381 11713 25415
rect 11747 25381 11759 25415
rect 11701 25375 11759 25381
rect 9631 25316 10180 25344
rect 9631 25313 9643 25316
rect 9585 25307 9643 25313
rect 8389 25279 8447 25285
rect 8389 25245 8401 25279
rect 8435 25276 8447 25279
rect 8435 25248 8984 25276
rect 8435 25245 8447 25248
rect 8389 25239 8447 25245
rect 8956 25149 8984 25248
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 10244 25276 10272 25372
rect 10318 25304 10324 25356
rect 10376 25304 10382 25356
rect 11716 25344 11744 25375
rect 12437 25347 12495 25353
rect 12437 25344 12449 25347
rect 11716 25316 12449 25344
rect 12437 25313 12449 25316
rect 12483 25313 12495 25347
rect 12437 25307 12495 25313
rect 10091 25248 10272 25276
rect 12621 25279 12679 25285
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 13372 25276 13400 25440
rect 15304 25412 15332 25440
rect 14752 25384 15332 25412
rect 14752 25353 14780 25384
rect 14737 25347 14795 25353
rect 14737 25313 14749 25347
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 14918 25304 14924 25356
rect 14976 25344 14982 25356
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 14976 25316 15301 25344
rect 14976 25304 14982 25316
rect 15289 25313 15301 25316
rect 15335 25344 15347 25347
rect 17126 25344 17132 25356
rect 15335 25316 17132 25344
rect 15335 25313 15347 25316
rect 15289 25307 15347 25313
rect 17126 25304 17132 25316
rect 17184 25344 17190 25356
rect 17313 25347 17371 25353
rect 17313 25344 17325 25347
rect 17184 25316 17325 25344
rect 17184 25304 17190 25316
rect 17313 25313 17325 25316
rect 17359 25344 17371 25347
rect 19536 25344 19564 25440
rect 31496 25412 31524 25440
rect 31665 25415 31723 25421
rect 31665 25412 31677 25415
rect 31496 25384 31677 25412
rect 31665 25381 31677 25384
rect 31711 25412 31723 25415
rect 33137 25415 33195 25421
rect 31711 25384 32812 25412
rect 31711 25381 31723 25384
rect 31665 25375 31723 25381
rect 17359 25316 19334 25344
rect 19536 25316 19656 25344
rect 17359 25313 17371 25316
rect 17313 25307 17371 25313
rect 12667 25248 13400 25276
rect 13817 25279 13875 25285
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 13817 25245 13829 25279
rect 13863 25276 13875 25279
rect 14553 25279 14611 25285
rect 13863 25248 14136 25276
rect 13863 25245 13875 25248
rect 13817 25239 13875 25245
rect 10588 25211 10646 25217
rect 10588 25177 10600 25211
rect 10634 25208 10646 25211
rect 10870 25208 10876 25220
rect 10634 25180 10876 25208
rect 10634 25177 10646 25180
rect 10588 25171 10646 25177
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 11606 25168 11612 25220
rect 11664 25168 11670 25220
rect 8941 25143 8999 25149
rect 8941 25109 8953 25143
rect 8987 25109 8999 25143
rect 8941 25103 8999 25109
rect 9401 25143 9459 25149
rect 9401 25109 9413 25143
rect 9447 25140 9459 25143
rect 11624 25140 11652 25168
rect 9447 25112 11652 25140
rect 9447 25109 9459 25112
rect 9401 25103 9459 25109
rect 13630 25100 13636 25152
rect 13688 25100 13694 25152
rect 14108 25149 14136 25248
rect 14553 25245 14565 25279
rect 14599 25276 14611 25279
rect 15194 25276 15200 25288
rect 14599 25248 15200 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 19306 25276 19334 25316
rect 19426 25276 19432 25288
rect 19306 25248 19432 25276
rect 19426 25236 19432 25248
rect 19484 25276 19490 25288
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19484 25248 19533 25276
rect 19484 25236 19490 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 19628 25276 19656 25316
rect 23750 25304 23756 25356
rect 23808 25344 23814 25356
rect 23845 25347 23903 25353
rect 23845 25344 23857 25347
rect 23808 25316 23857 25344
rect 23808 25304 23814 25316
rect 23845 25313 23857 25316
rect 23891 25313 23903 25347
rect 23845 25307 23903 25313
rect 24118 25304 24124 25356
rect 24176 25304 24182 25356
rect 24762 25304 24768 25356
rect 24820 25344 24826 25356
rect 27249 25347 27307 25353
rect 27249 25344 27261 25347
rect 24820 25316 27261 25344
rect 24820 25304 24826 25316
rect 27249 25313 27261 25316
rect 27295 25344 27307 25347
rect 27522 25344 27528 25356
rect 27295 25316 27528 25344
rect 27295 25313 27307 25316
rect 27249 25307 27307 25313
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 29086 25304 29092 25356
rect 29144 25304 29150 25356
rect 29365 25347 29423 25353
rect 29365 25313 29377 25347
rect 29411 25344 29423 25347
rect 32122 25344 32128 25356
rect 29411 25316 32128 25344
rect 29411 25313 29423 25316
rect 29365 25307 29423 25313
rect 32122 25304 32128 25316
rect 32180 25304 32186 25356
rect 32784 25344 32812 25384
rect 33137 25381 33149 25415
rect 33183 25412 33195 25415
rect 33594 25412 33600 25424
rect 33183 25384 33600 25412
rect 33183 25381 33195 25384
rect 33137 25375 33195 25381
rect 33594 25372 33600 25384
rect 33652 25372 33658 25424
rect 33229 25347 33287 25353
rect 33229 25344 33241 25347
rect 32784 25316 33241 25344
rect 33229 25313 33241 25316
rect 33275 25344 33287 25347
rect 33410 25344 33416 25356
rect 33275 25316 33416 25344
rect 33275 25313 33287 25316
rect 33229 25307 33287 25313
rect 33410 25304 33416 25316
rect 33468 25304 33474 25356
rect 19777 25279 19835 25285
rect 19777 25276 19789 25279
rect 19628 25248 19789 25276
rect 19521 25239 19579 25245
rect 19777 25245 19789 25248
rect 19823 25245 19835 25279
rect 28997 25279 29055 25285
rect 28997 25276 29009 25279
rect 19777 25239 19835 25245
rect 25976 25248 29009 25276
rect 14461 25211 14519 25217
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 14826 25208 14832 25220
rect 14507 25180 14832 25208
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 16790 25180 16896 25208
rect 14093 25143 14151 25149
rect 14093 25109 14105 25143
rect 14139 25109 14151 25143
rect 16868 25140 16896 25180
rect 17586 25168 17592 25220
rect 17644 25168 17650 25220
rect 18046 25208 18052 25220
rect 17696 25180 18052 25208
rect 17696 25140 17724 25180
rect 18046 25168 18052 25180
rect 18104 25168 18110 25220
rect 18138 25168 18144 25220
rect 18196 25168 18202 25220
rect 24670 25208 24676 25220
rect 23414 25180 24676 25208
rect 24670 25168 24676 25180
rect 24728 25208 24734 25220
rect 24946 25208 24952 25220
rect 24728 25180 24952 25208
rect 24728 25168 24734 25180
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 16868 25112 17724 25140
rect 14093 25103 14151 25109
rect 22370 25100 22376 25152
rect 22428 25140 22434 25152
rect 25976 25140 26004 25248
rect 28997 25245 29009 25248
rect 29043 25276 29055 25279
rect 29733 25279 29791 25285
rect 29733 25276 29745 25279
rect 29043 25248 29745 25276
rect 29043 25245 29055 25248
rect 28997 25239 29055 25245
rect 29733 25245 29745 25248
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25276 31723 25279
rect 31938 25276 31944 25288
rect 31711 25248 31944 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 27065 25211 27123 25217
rect 27065 25177 27077 25211
rect 27111 25208 27123 25211
rect 27111 25180 29040 25208
rect 27111 25177 27123 25180
rect 27065 25171 27123 25177
rect 29012 25152 29040 25180
rect 29822 25168 29828 25220
rect 29880 25208 29886 25220
rect 29917 25211 29975 25217
rect 29917 25208 29929 25211
rect 29880 25180 29929 25208
rect 29880 25168 29886 25180
rect 29917 25177 29929 25180
rect 29963 25177 29975 25211
rect 31496 25208 31524 25239
rect 31938 25236 31944 25248
rect 31996 25236 32002 25288
rect 32033 25279 32091 25285
rect 32033 25245 32045 25279
rect 32079 25245 32091 25279
rect 32033 25239 32091 25245
rect 32048 25208 32076 25239
rect 31496 25180 31754 25208
rect 29917 25171 29975 25177
rect 22428 25112 26004 25140
rect 22428 25100 22434 25112
rect 27154 25100 27160 25152
rect 27212 25100 27218 25152
rect 28994 25100 29000 25152
rect 29052 25100 29058 25152
rect 31726 25140 31754 25180
rect 31864 25180 32076 25208
rect 32140 25208 32168 25304
rect 32214 25236 32220 25288
rect 32272 25276 32278 25288
rect 32677 25279 32735 25285
rect 32677 25276 32689 25279
rect 32272 25248 32689 25276
rect 32272 25236 32278 25248
rect 32677 25245 32689 25248
rect 32723 25245 32735 25279
rect 32677 25239 32735 25245
rect 33045 25279 33103 25285
rect 33045 25245 33057 25279
rect 33091 25245 33103 25279
rect 33045 25239 33103 25245
rect 32493 25211 32551 25217
rect 32493 25208 32505 25211
rect 32140 25180 32505 25208
rect 31864 25152 31892 25180
rect 32493 25177 32505 25180
rect 32539 25177 32551 25211
rect 32493 25171 32551 25177
rect 33060 25208 33088 25239
rect 33318 25236 33324 25288
rect 33376 25236 33382 25288
rect 33505 25279 33563 25285
rect 33505 25245 33517 25279
rect 33551 25276 33563 25279
rect 33689 25279 33747 25285
rect 33689 25276 33701 25279
rect 33551 25248 33701 25276
rect 33551 25245 33563 25248
rect 33505 25239 33563 25245
rect 33689 25245 33701 25248
rect 33735 25245 33747 25279
rect 33689 25239 33747 25245
rect 33796 25208 33824 25452
rect 36262 25440 36268 25452
rect 36320 25440 36326 25492
rect 37829 25483 37887 25489
rect 37829 25449 37841 25483
rect 37875 25480 37887 25483
rect 38378 25480 38384 25492
rect 37875 25452 38384 25480
rect 37875 25449 37887 25452
rect 37829 25443 37887 25449
rect 38378 25440 38384 25452
rect 38436 25440 38442 25492
rect 38654 25440 38660 25492
rect 38712 25440 38718 25492
rect 43349 25483 43407 25489
rect 43349 25480 43361 25483
rect 41984 25452 43361 25480
rect 34241 25415 34299 25421
rect 34241 25381 34253 25415
rect 34287 25381 34299 25415
rect 34241 25375 34299 25381
rect 34256 25344 34284 25375
rect 36265 25347 36323 25353
rect 36265 25344 36277 25347
rect 34256 25316 36277 25344
rect 36265 25313 36277 25316
rect 36311 25313 36323 25347
rect 36265 25307 36323 25313
rect 36541 25347 36599 25353
rect 36541 25313 36553 25347
rect 36587 25344 36599 25347
rect 37274 25344 37280 25356
rect 36587 25316 37280 25344
rect 36587 25313 36599 25316
rect 36541 25307 36599 25313
rect 37274 25304 37280 25316
rect 37332 25304 37338 25356
rect 38197 25347 38255 25353
rect 38197 25313 38209 25347
rect 38243 25344 38255 25347
rect 38470 25344 38476 25356
rect 38243 25316 38476 25344
rect 38243 25313 38255 25316
rect 38197 25307 38255 25313
rect 38470 25304 38476 25316
rect 38528 25304 38534 25356
rect 34054 25236 34060 25288
rect 34112 25236 34118 25288
rect 36906 25236 36912 25288
rect 36964 25236 36970 25288
rect 38105 25279 38163 25285
rect 38105 25245 38117 25279
rect 38151 25276 38163 25279
rect 38672 25276 38700 25440
rect 41984 25285 42012 25452
rect 43349 25449 43361 25452
rect 43395 25480 43407 25483
rect 43530 25480 43536 25492
rect 43395 25452 43536 25480
rect 43395 25449 43407 25452
rect 43349 25443 43407 25449
rect 43530 25440 43536 25452
rect 43588 25440 43594 25492
rect 42058 25372 42064 25424
rect 42116 25372 42122 25424
rect 42245 25415 42303 25421
rect 42245 25381 42257 25415
rect 42291 25381 42303 25415
rect 42245 25375 42303 25381
rect 42076 25285 42104 25372
rect 42260 25344 42288 25375
rect 43901 25347 43959 25353
rect 43901 25344 43913 25347
rect 42260 25316 43913 25344
rect 43901 25313 43913 25316
rect 43947 25313 43959 25347
rect 43901 25307 43959 25313
rect 38151 25248 38700 25276
rect 41969 25279 42027 25285
rect 38151 25245 38163 25248
rect 38105 25239 38163 25245
rect 41969 25245 41981 25279
rect 42015 25245 42027 25279
rect 41969 25239 42027 25245
rect 42061 25279 42119 25285
rect 42061 25245 42073 25279
rect 42107 25245 42119 25279
rect 42061 25239 42119 25245
rect 42245 25279 42303 25285
rect 42245 25245 42257 25279
rect 42291 25276 42303 25279
rect 42794 25276 42800 25288
rect 42291 25248 42800 25276
rect 42291 25245 42303 25248
rect 42245 25239 42303 25245
rect 42794 25236 42800 25248
rect 42852 25236 42858 25288
rect 42886 25236 42892 25288
rect 42944 25236 42950 25288
rect 43165 25279 43223 25285
rect 43165 25245 43177 25279
rect 43211 25245 43223 25279
rect 43165 25239 43223 25245
rect 44545 25279 44603 25285
rect 44545 25245 44557 25279
rect 44591 25276 44603 25279
rect 44637 25279 44695 25285
rect 44637 25276 44649 25279
rect 44591 25248 44649 25276
rect 44591 25245 44603 25248
rect 44545 25239 44603 25245
rect 44637 25245 44649 25248
rect 44683 25245 44695 25279
rect 44637 25239 44695 25245
rect 44821 25279 44879 25285
rect 44821 25245 44833 25279
rect 44867 25245 44879 25279
rect 44821 25239 44879 25245
rect 33060 25180 33824 25208
rect 31846 25140 31852 25152
rect 31726 25112 31852 25140
rect 31846 25100 31852 25112
rect 31904 25100 31910 25152
rect 32398 25100 32404 25152
rect 32456 25140 32462 25152
rect 33060 25140 33088 25180
rect 33870 25168 33876 25220
rect 33928 25168 33934 25220
rect 33962 25168 33968 25220
rect 34020 25168 34026 25220
rect 32456 25112 33088 25140
rect 32456 25100 32462 25112
rect 33134 25100 33140 25152
rect 33192 25140 33198 25152
rect 34072 25140 34100 25236
rect 36924 25208 36952 25236
rect 42978 25208 42984 25220
rect 35834 25180 36952 25208
rect 42812 25180 42984 25208
rect 42812 25152 42840 25180
rect 42978 25168 42984 25180
rect 43036 25208 43042 25220
rect 43180 25208 43208 25239
rect 43036 25180 43208 25208
rect 43036 25168 43042 25180
rect 43254 25168 43260 25220
rect 43312 25208 43318 25220
rect 44836 25208 44864 25239
rect 43312 25180 44864 25208
rect 43312 25168 43318 25180
rect 33192 25112 34100 25140
rect 33192 25100 33198 25112
rect 34790 25100 34796 25152
rect 34848 25140 34854 25152
rect 34974 25140 34980 25152
rect 34848 25112 34980 25140
rect 34848 25100 34854 25112
rect 34974 25100 34980 25112
rect 35032 25100 35038 25152
rect 42334 25100 42340 25152
rect 42392 25100 42398 25152
rect 42794 25100 42800 25152
rect 42852 25100 42858 25152
rect 44358 25100 44364 25152
rect 44416 25140 44422 25152
rect 44729 25143 44787 25149
rect 44729 25140 44741 25143
rect 44416 25112 44741 25140
rect 44416 25100 44422 25112
rect 44729 25109 44741 25112
rect 44775 25109 44787 25143
rect 44729 25103 44787 25109
rect 1104 25050 45172 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 45172 25050
rect 1104 24976 45172 24998
rect 10870 24896 10876 24948
rect 10928 24896 10934 24948
rect 11517 24939 11575 24945
rect 11517 24905 11529 24939
rect 11563 24936 11575 24939
rect 11606 24936 11612 24948
rect 11563 24908 11612 24936
rect 11563 24905 11575 24908
rect 11517 24899 11575 24905
rect 11606 24896 11612 24908
rect 11664 24896 11670 24948
rect 13446 24896 13452 24948
rect 13504 24896 13510 24948
rect 14737 24939 14795 24945
rect 14737 24905 14749 24939
rect 14783 24936 14795 24939
rect 14826 24936 14832 24948
rect 14783 24908 14832 24936
rect 14783 24905 14795 24908
rect 14737 24899 14795 24905
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 16206 24896 16212 24948
rect 16264 24896 16270 24948
rect 16758 24896 16764 24948
rect 16816 24896 16822 24948
rect 17034 24896 17040 24948
rect 17092 24936 17098 24948
rect 17129 24939 17187 24945
rect 17129 24936 17141 24939
rect 17092 24908 17141 24936
rect 17092 24896 17098 24908
rect 17129 24905 17141 24908
rect 17175 24905 17187 24939
rect 17129 24899 17187 24905
rect 17586 24896 17592 24948
rect 17644 24936 17650 24948
rect 17681 24939 17739 24945
rect 17681 24936 17693 24939
rect 17644 24908 17693 24936
rect 17644 24896 17650 24908
rect 17681 24905 17693 24908
rect 17727 24905 17739 24939
rect 17681 24899 17739 24905
rect 18322 24896 18328 24948
rect 18380 24896 18386 24948
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19889 24939 19947 24945
rect 19889 24936 19901 24939
rect 19392 24908 19901 24936
rect 19392 24896 19398 24908
rect 19889 24905 19901 24908
rect 19935 24905 19947 24939
rect 19889 24899 19947 24905
rect 20254 24896 20260 24948
rect 20312 24896 20318 24948
rect 22370 24896 22376 24948
rect 22428 24936 22434 24948
rect 23017 24939 23075 24945
rect 23017 24936 23029 24939
rect 22428 24908 23029 24936
rect 22428 24896 22434 24908
rect 23017 24905 23029 24908
rect 23063 24905 23075 24939
rect 23017 24899 23075 24905
rect 23385 24939 23443 24945
rect 23385 24905 23397 24939
rect 23431 24936 23443 24939
rect 23566 24936 23572 24948
rect 23431 24908 23572 24936
rect 23431 24905 23443 24908
rect 23385 24899 23443 24905
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 24857 24939 24915 24945
rect 24857 24905 24869 24939
rect 24903 24905 24915 24939
rect 24857 24899 24915 24905
rect 13464 24868 13492 24896
rect 13004 24840 13492 24868
rect 11057 24803 11115 24809
rect 11057 24769 11069 24803
rect 11103 24800 11115 24803
rect 11514 24800 11520 24812
rect 11103 24772 11520 24800
rect 11103 24769 11115 24772
rect 11057 24763 11115 24769
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11882 24760 11888 24812
rect 11940 24800 11946 24812
rect 13004 24809 13032 24840
rect 13722 24828 13728 24880
rect 13780 24828 13786 24880
rect 24872 24868 24900 24899
rect 24946 24896 24952 24948
rect 25004 24936 25010 24948
rect 25004 24908 25636 24936
rect 25004 24896 25010 24908
rect 25225 24871 25283 24877
rect 25225 24868 25237 24871
rect 17788 24840 18092 24868
rect 24872 24840 25237 24868
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11940 24772 12081 24800
rect 11940 24760 11946 24772
rect 12069 24769 12081 24772
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 14829 24803 14887 24809
rect 14829 24769 14841 24803
rect 14875 24800 14887 24803
rect 14918 24800 14924 24812
rect 14875 24772 14924 24800
rect 14875 24769 14887 24772
rect 14829 24763 14887 24769
rect 14918 24760 14924 24772
rect 14976 24760 14982 24812
rect 15102 24809 15108 24812
rect 15096 24763 15108 24809
rect 15102 24760 15108 24763
rect 15160 24760 15166 24812
rect 15838 24760 15844 24812
rect 15896 24800 15902 24812
rect 17788 24800 17816 24840
rect 15896 24772 17816 24800
rect 17865 24803 17923 24809
rect 15896 24760 15902 24772
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 18064 24800 18092 24840
rect 25225 24837 25237 24840
rect 25271 24837 25283 24871
rect 25608 24868 25636 24908
rect 26970 24896 26976 24948
rect 27028 24936 27034 24948
rect 27249 24939 27307 24945
rect 27249 24936 27261 24939
rect 27028 24908 27261 24936
rect 27028 24896 27034 24908
rect 27249 24905 27261 24908
rect 27295 24905 27307 24939
rect 27249 24899 27307 24905
rect 28997 24939 29055 24945
rect 28997 24905 29009 24939
rect 29043 24936 29055 24939
rect 29086 24936 29092 24948
rect 29043 24908 29092 24936
rect 29043 24905 29055 24908
rect 28997 24899 29055 24905
rect 29086 24896 29092 24908
rect 29144 24896 29150 24948
rect 29270 24896 29276 24948
rect 29328 24936 29334 24948
rect 29914 24936 29920 24948
rect 29328 24908 29920 24936
rect 29328 24896 29334 24908
rect 29914 24896 29920 24908
rect 29972 24936 29978 24948
rect 30377 24939 30435 24945
rect 30377 24936 30389 24939
rect 29972 24908 30389 24936
rect 29972 24896 29978 24908
rect 30377 24905 30389 24908
rect 30423 24905 30435 24939
rect 30377 24899 30435 24905
rect 31938 24896 31944 24948
rect 31996 24936 32002 24948
rect 31996 24908 32444 24936
rect 31996 24896 32002 24908
rect 25608 24840 25714 24868
rect 29196 24840 30604 24868
rect 25225 24831 25283 24837
rect 22002 24800 22008 24812
rect 17911 24772 18000 24800
rect 18064 24772 22008 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13630 24732 13636 24744
rect 13311 24704 13636 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13630 24692 13636 24704
rect 13688 24692 13694 24744
rect 17218 24692 17224 24744
rect 17276 24692 17282 24744
rect 17405 24735 17463 24741
rect 17405 24701 17417 24735
rect 17451 24732 17463 24735
rect 17451 24704 17908 24732
rect 17451 24701 17463 24704
rect 17405 24695 17463 24701
rect 17880 24596 17908 24704
rect 17972 24673 18000 24772
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 22925 24803 22983 24809
rect 22925 24800 22937 24803
rect 22603 24772 22937 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 22925 24769 22937 24772
rect 22971 24769 22983 24803
rect 22925 24763 22983 24769
rect 24670 24760 24676 24812
rect 24728 24760 24734 24812
rect 28718 24760 28724 24812
rect 28776 24760 28782 24812
rect 29196 24809 29224 24840
rect 29181 24803 29239 24809
rect 29181 24769 29193 24803
rect 29227 24800 29239 24803
rect 29270 24800 29276 24812
rect 29227 24772 29276 24800
rect 29227 24769 29239 24772
rect 29181 24763 29239 24769
rect 29270 24760 29276 24772
rect 29328 24760 29334 24812
rect 29822 24800 29828 24812
rect 29472 24772 29828 24800
rect 18414 24692 18420 24744
rect 18472 24692 18478 24744
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 20346 24692 20352 24744
rect 20404 24692 20410 24744
rect 20530 24692 20536 24744
rect 20588 24692 20594 24744
rect 21910 24692 21916 24744
rect 21968 24692 21974 24744
rect 22833 24735 22891 24741
rect 22833 24701 22845 24735
rect 22879 24732 22891 24735
rect 24762 24732 24768 24744
rect 22879 24704 24768 24732
rect 22879 24701 22891 24704
rect 22833 24695 22891 24701
rect 24762 24692 24768 24704
rect 24820 24692 24826 24744
rect 29472 24741 29500 24772
rect 29822 24760 29828 24772
rect 29880 24760 29886 24812
rect 30576 24809 30604 24840
rect 31846 24828 31852 24880
rect 31904 24868 31910 24880
rect 32214 24868 32220 24880
rect 31904 24840 32220 24868
rect 31904 24828 31910 24840
rect 32214 24828 32220 24840
rect 32272 24828 32278 24880
rect 32416 24877 32444 24908
rect 33318 24896 33324 24948
rect 33376 24896 33382 24948
rect 33597 24939 33655 24945
rect 33597 24905 33609 24939
rect 33643 24936 33655 24939
rect 33870 24936 33876 24948
rect 33643 24908 33876 24936
rect 33643 24905 33655 24908
rect 33597 24899 33655 24905
rect 33870 24896 33876 24908
rect 33928 24896 33934 24948
rect 33962 24896 33968 24948
rect 34020 24936 34026 24948
rect 34425 24939 34483 24945
rect 34425 24936 34437 24939
rect 34020 24908 34437 24936
rect 34020 24896 34026 24908
rect 34425 24905 34437 24908
rect 34471 24905 34483 24939
rect 34425 24899 34483 24905
rect 39482 24896 39488 24948
rect 39540 24896 39546 24948
rect 42981 24939 43039 24945
rect 42981 24905 42993 24939
rect 43027 24936 43039 24939
rect 43254 24936 43260 24948
rect 43027 24908 43260 24936
rect 43027 24905 43039 24908
rect 42981 24899 43039 24905
rect 32401 24871 32459 24877
rect 32401 24837 32413 24871
rect 32447 24837 32459 24871
rect 32401 24831 32459 24837
rect 32585 24871 32643 24877
rect 32585 24837 32597 24871
rect 32631 24868 32643 24871
rect 33336 24868 33364 24896
rect 32631 24840 33364 24868
rect 32631 24837 32643 24840
rect 32585 24831 32643 24837
rect 30561 24803 30619 24809
rect 30561 24769 30573 24803
rect 30607 24769 30619 24803
rect 32122 24800 32128 24812
rect 30561 24763 30619 24769
rect 31772 24772 32128 24800
rect 24949 24735 25007 24741
rect 24949 24701 24961 24735
rect 24995 24701 25007 24735
rect 29457 24735 29515 24741
rect 29457 24732 29469 24735
rect 24949 24695 25007 24701
rect 28644 24704 29469 24732
rect 17957 24667 18015 24673
rect 17957 24633 17969 24667
rect 18003 24633 18015 24667
rect 17957 24627 18015 24633
rect 18616 24596 18644 24692
rect 24964 24608 24992 24695
rect 26970 24664 26976 24676
rect 26252 24636 26976 24664
rect 17880 24568 18644 24596
rect 24946 24556 24952 24608
rect 25004 24596 25010 24608
rect 26252 24596 26280 24636
rect 26970 24624 26976 24636
rect 27028 24624 27034 24676
rect 25004 24568 26280 24596
rect 25004 24556 25010 24568
rect 26694 24556 26700 24608
rect 26752 24596 26758 24608
rect 28644 24596 28672 24704
rect 29457 24701 29469 24704
rect 29503 24701 29515 24735
rect 29457 24695 29515 24701
rect 29730 24692 29736 24744
rect 29788 24692 29794 24744
rect 30193 24735 30251 24741
rect 30193 24701 30205 24735
rect 30239 24732 30251 24735
rect 31772 24732 31800 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32600 24800 32628 24831
rect 33336 24809 33364 24840
rect 34054 24828 34060 24880
rect 34112 24868 34118 24880
rect 35434 24868 35440 24880
rect 34112 24840 35440 24868
rect 34112 24828 34118 24840
rect 35434 24828 35440 24840
rect 35492 24828 35498 24880
rect 38841 24871 38899 24877
rect 38841 24837 38853 24871
rect 38887 24868 38899 24871
rect 39500 24868 39528 24896
rect 38887 24840 39528 24868
rect 42613 24871 42671 24877
rect 38887 24837 38899 24840
rect 38841 24831 38899 24837
rect 39132 24812 39160 24840
rect 42613 24837 42625 24871
rect 42659 24868 42671 24871
rect 42702 24868 42708 24880
rect 42659 24840 42708 24868
rect 42659 24837 42671 24840
rect 42613 24831 42671 24837
rect 42702 24828 42708 24840
rect 42760 24828 42766 24880
rect 42794 24828 42800 24880
rect 42852 24877 42858 24880
rect 42852 24871 42871 24877
rect 42859 24837 42871 24871
rect 42852 24831 42871 24837
rect 42852 24828 42858 24831
rect 32309 24763 32367 24769
rect 32508 24772 32628 24800
rect 32769 24803 32827 24809
rect 32318 24732 32346 24763
rect 30239 24704 31800 24732
rect 32048 24704 32346 24732
rect 30239 24701 30251 24704
rect 30193 24695 30251 24701
rect 26752 24568 28672 24596
rect 29365 24599 29423 24605
rect 26752 24556 26758 24568
rect 29365 24565 29377 24599
rect 29411 24596 29423 24599
rect 29454 24596 29460 24608
rect 29411 24568 29460 24596
rect 29411 24565 29423 24568
rect 29365 24559 29423 24565
rect 29454 24556 29460 24568
rect 29512 24556 29518 24608
rect 32048 24596 32076 24704
rect 32125 24667 32183 24673
rect 32125 24633 32137 24667
rect 32171 24664 32183 24667
rect 32508 24664 32536 24772
rect 32769 24769 32781 24803
rect 32815 24800 32827 24803
rect 32861 24803 32919 24809
rect 32861 24800 32873 24803
rect 32815 24772 32873 24800
rect 32815 24769 32827 24772
rect 32769 24763 32827 24769
rect 32861 24769 32873 24772
rect 32907 24769 32919 24803
rect 32861 24763 32919 24769
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33321 24803 33379 24809
rect 33321 24769 33333 24803
rect 33367 24769 33379 24803
rect 33321 24763 33379 24769
rect 32171 24636 32536 24664
rect 32171 24633 32183 24636
rect 32125 24627 32183 24633
rect 32674 24624 32680 24676
rect 32732 24664 32738 24676
rect 33060 24664 33088 24763
rect 33410 24760 33416 24812
rect 33468 24760 33474 24812
rect 34974 24760 34980 24812
rect 35032 24760 35038 24812
rect 38105 24803 38163 24809
rect 38105 24769 38117 24803
rect 38151 24800 38163 24803
rect 38197 24803 38255 24809
rect 38197 24800 38209 24803
rect 38151 24772 38209 24800
rect 38151 24769 38163 24772
rect 38105 24763 38163 24769
rect 38197 24769 38209 24772
rect 38243 24769 38255 24803
rect 38197 24763 38255 24769
rect 38381 24803 38439 24809
rect 38381 24769 38393 24803
rect 38427 24800 38439 24803
rect 38657 24803 38715 24809
rect 38657 24800 38669 24803
rect 38427 24772 38669 24800
rect 38427 24769 38439 24772
rect 38381 24763 38439 24769
rect 38657 24769 38669 24772
rect 38703 24769 38715 24803
rect 38657 24763 38715 24769
rect 39025 24803 39083 24809
rect 39025 24769 39037 24803
rect 39071 24769 39083 24803
rect 39025 24763 39083 24769
rect 33226 24692 33232 24744
rect 33284 24692 33290 24744
rect 33594 24692 33600 24744
rect 33652 24692 33658 24744
rect 38470 24692 38476 24744
rect 38528 24732 38534 24744
rect 38565 24735 38623 24741
rect 38565 24732 38577 24735
rect 38528 24704 38577 24732
rect 38528 24692 38534 24704
rect 38565 24701 38577 24704
rect 38611 24701 38623 24735
rect 39040 24732 39068 24763
rect 39114 24760 39120 24812
rect 39172 24760 39178 24812
rect 39301 24803 39359 24809
rect 39301 24769 39313 24803
rect 39347 24800 39359 24803
rect 39347 24772 39436 24800
rect 39347 24769 39359 24772
rect 39301 24763 39359 24769
rect 39408 24744 39436 24772
rect 40034 24760 40040 24812
rect 40092 24800 40098 24812
rect 40497 24803 40555 24809
rect 40497 24800 40509 24803
rect 40092 24772 40509 24800
rect 40092 24760 40098 24772
rect 40497 24769 40509 24772
rect 40543 24769 40555 24803
rect 40497 24763 40555 24769
rect 40589 24803 40647 24809
rect 40589 24769 40601 24803
rect 40635 24800 40647 24803
rect 40678 24800 40684 24812
rect 40635 24772 40684 24800
rect 40635 24769 40647 24772
rect 40589 24763 40647 24769
rect 40678 24760 40684 24772
rect 40736 24760 40742 24812
rect 40770 24760 40776 24812
rect 40828 24760 40834 24812
rect 41693 24803 41751 24809
rect 41693 24769 41705 24803
rect 41739 24769 41751 24803
rect 41693 24763 41751 24769
rect 41877 24803 41935 24809
rect 41877 24769 41889 24803
rect 41923 24800 41935 24803
rect 42334 24800 42340 24812
rect 41923 24772 42340 24800
rect 41923 24769 41935 24772
rect 41877 24763 41935 24769
rect 39390 24732 39396 24744
rect 39040 24704 39396 24732
rect 38565 24695 38623 24701
rect 32732 24636 33088 24664
rect 32732 24624 32738 24636
rect 33244 24596 33272 24692
rect 38580 24664 38608 24695
rect 39390 24692 39396 24704
rect 39448 24692 39454 24744
rect 41598 24692 41604 24744
rect 41656 24732 41662 24744
rect 41708 24732 41736 24763
rect 42334 24760 42340 24772
rect 42392 24760 42398 24812
rect 42996 24732 43024 24899
rect 43254 24896 43260 24908
rect 43312 24896 43318 24948
rect 43070 24760 43076 24812
rect 43128 24760 43134 24812
rect 41656 24704 43024 24732
rect 41656 24692 41662 24704
rect 39209 24667 39267 24673
rect 39209 24664 39221 24667
rect 38580 24636 39221 24664
rect 39209 24633 39221 24636
rect 39255 24633 39267 24667
rect 43714 24664 43720 24676
rect 39209 24627 39267 24633
rect 39316 24636 43720 24664
rect 32048 24568 33272 24596
rect 37734 24556 37740 24608
rect 37792 24596 37798 24608
rect 37921 24599 37979 24605
rect 37921 24596 37933 24599
rect 37792 24568 37933 24596
rect 37792 24556 37798 24568
rect 37921 24565 37933 24568
rect 37967 24565 37979 24599
rect 37921 24559 37979 24565
rect 38746 24556 38752 24608
rect 38804 24596 38810 24608
rect 39316 24596 39344 24636
rect 43714 24624 43720 24636
rect 43772 24624 43778 24676
rect 38804 24568 39344 24596
rect 38804 24556 38810 24568
rect 40126 24556 40132 24608
rect 40184 24596 40190 24608
rect 40773 24599 40831 24605
rect 40773 24596 40785 24599
rect 40184 24568 40785 24596
rect 40184 24556 40190 24568
rect 40773 24565 40785 24568
rect 40819 24565 40831 24599
rect 40773 24559 40831 24565
rect 41690 24556 41696 24608
rect 41748 24556 41754 24608
rect 42797 24599 42855 24605
rect 42797 24565 42809 24599
rect 42843 24596 42855 24599
rect 43162 24596 43168 24608
rect 42843 24568 43168 24596
rect 42843 24565 42855 24568
rect 42797 24559 42855 24565
rect 43162 24556 43168 24568
rect 43220 24556 43226 24608
rect 44542 24556 44548 24608
rect 44600 24556 44606 24608
rect 1104 24506 45172 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 45172 24506
rect 1104 24432 45172 24454
rect 8018 24352 8024 24404
rect 8076 24392 8082 24404
rect 11054 24392 11060 24404
rect 8076 24364 11060 24392
rect 8076 24352 8082 24364
rect 11054 24352 11060 24364
rect 11112 24352 11118 24404
rect 15013 24395 15071 24401
rect 15013 24361 15025 24395
rect 15059 24392 15071 24395
rect 15102 24392 15108 24404
rect 15059 24364 15108 24392
rect 15059 24361 15071 24364
rect 15013 24355 15071 24361
rect 15102 24352 15108 24364
rect 15160 24352 15166 24404
rect 15838 24352 15844 24404
rect 15896 24352 15902 24404
rect 16758 24352 16764 24404
rect 16816 24392 16822 24404
rect 16816 24364 18092 24392
rect 16816 24352 16822 24364
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 11609 24327 11667 24333
rect 11609 24324 11621 24327
rect 11020 24296 11621 24324
rect 11020 24284 11026 24296
rect 11609 24293 11621 24296
rect 11655 24324 11667 24327
rect 14274 24324 14280 24336
rect 11655 24296 14280 24324
rect 11655 24293 11667 24296
rect 11609 24287 11667 24293
rect 14274 24284 14280 24296
rect 14332 24284 14338 24336
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24256 10103 24259
rect 11238 24256 11244 24268
rect 10091 24228 11244 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 12345 24259 12403 24265
rect 12345 24225 12357 24259
rect 12391 24256 12403 24259
rect 12434 24256 12440 24268
rect 12391 24228 12440 24256
rect 12391 24225 12403 24228
rect 12345 24219 12403 24225
rect 12434 24216 12440 24228
rect 12492 24256 12498 24268
rect 12802 24256 12808 24268
rect 12492 24228 12808 24256
rect 12492 24216 12498 24228
rect 12802 24216 12808 24228
rect 12860 24256 12866 24268
rect 14369 24259 14427 24265
rect 14369 24256 14381 24259
rect 12860 24228 14381 24256
rect 12860 24216 12866 24228
rect 14369 24225 14381 24228
rect 14415 24256 14427 24259
rect 15749 24259 15807 24265
rect 15749 24256 15761 24259
rect 14415 24228 15761 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 15749 24225 15761 24228
rect 15795 24256 15807 24259
rect 15856 24256 15884 24352
rect 18064 24324 18092 24364
rect 18690 24352 18696 24404
rect 18748 24392 18754 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 18748 24364 19257 24392
rect 18748 24352 18754 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 24670 24352 24676 24404
rect 24728 24392 24734 24404
rect 24857 24395 24915 24401
rect 24857 24392 24869 24395
rect 24728 24364 24869 24392
rect 24728 24352 24734 24364
rect 24857 24361 24869 24364
rect 24903 24361 24915 24395
rect 24857 24355 24915 24361
rect 29270 24352 29276 24404
rect 29328 24352 29334 24404
rect 29730 24352 29736 24404
rect 29788 24352 29794 24404
rect 32122 24352 32128 24404
rect 32180 24392 32186 24404
rect 32674 24392 32680 24404
rect 32180 24364 32680 24392
rect 32180 24352 32186 24364
rect 32674 24352 32680 24364
rect 32732 24352 32738 24404
rect 37632 24395 37690 24401
rect 37632 24361 37644 24395
rect 37678 24392 37690 24395
rect 37734 24392 37740 24404
rect 37678 24364 37740 24392
rect 37678 24361 37690 24364
rect 37632 24355 37690 24361
rect 37734 24352 37740 24364
rect 37792 24352 37798 24404
rect 39114 24352 39120 24404
rect 39172 24352 39178 24404
rect 40037 24395 40095 24401
rect 40037 24361 40049 24395
rect 40083 24392 40095 24395
rect 41782 24392 41788 24404
rect 40083 24364 41788 24392
rect 40083 24361 40095 24364
rect 40037 24355 40095 24361
rect 41782 24352 41788 24364
rect 41840 24352 41846 24404
rect 42702 24352 42708 24404
rect 42760 24392 42766 24404
rect 42889 24395 42947 24401
rect 42889 24392 42901 24395
rect 42760 24364 42901 24392
rect 42760 24352 42766 24364
rect 42889 24361 42901 24364
rect 42935 24361 42947 24395
rect 42889 24355 42947 24361
rect 44542 24352 44548 24404
rect 44600 24352 44606 24404
rect 22370 24324 22376 24336
rect 18064 24296 22376 24324
rect 22370 24284 22376 24296
rect 22428 24324 22434 24336
rect 27154 24324 27160 24336
rect 22428 24296 27160 24324
rect 22428 24284 22434 24296
rect 27154 24284 27160 24296
rect 27212 24284 27218 24336
rect 31938 24284 31944 24336
rect 31996 24324 32002 24336
rect 32858 24324 32864 24336
rect 31996 24296 32864 24324
rect 31996 24284 32002 24296
rect 32858 24284 32864 24296
rect 32916 24284 32922 24336
rect 40770 24284 40776 24336
rect 40828 24324 40834 24336
rect 40957 24327 41015 24333
rect 40957 24324 40969 24327
rect 40828 24296 40969 24324
rect 40828 24284 40834 24296
rect 40957 24293 40969 24296
rect 41003 24293 41015 24327
rect 40957 24287 41015 24293
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 15795 24228 15884 24256
rect 17972 24228 18429 24256
rect 15795 24225 15807 24228
rect 15749 24219 15807 24225
rect 10410 24148 10416 24200
rect 10468 24148 10474 24200
rect 10873 24191 10931 24197
rect 10873 24157 10885 24191
rect 10919 24188 10931 24191
rect 10962 24188 10968 24200
rect 10919 24160 10968 24188
rect 10919 24157 10931 24160
rect 10873 24151 10931 24157
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11790 24188 11796 24200
rect 11112 24160 11796 24188
rect 11112 24148 11118 24160
rect 11790 24148 11796 24160
rect 11848 24148 11854 24200
rect 12066 24148 12072 24200
rect 12124 24148 12130 24200
rect 14090 24148 14096 24200
rect 14148 24148 14154 24200
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24188 14887 24191
rect 14875 24160 15148 24188
rect 14875 24157 14887 24160
rect 14829 24151 14887 24157
rect 9861 24123 9919 24129
rect 9861 24089 9873 24123
rect 9907 24120 9919 24123
rect 12618 24120 12624 24132
rect 9907 24092 10824 24120
rect 9907 24089 9919 24092
rect 9861 24083 9919 24089
rect 9214 24012 9220 24064
rect 9272 24052 9278 24064
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 9272 24024 9413 24052
rect 9272 24012 9278 24024
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 9766 24012 9772 24064
rect 9824 24012 9830 24064
rect 10226 24012 10232 24064
rect 10284 24012 10290 24064
rect 10594 24012 10600 24064
rect 10652 24012 10658 24064
rect 10796 24052 10824 24092
rect 11164 24092 12624 24120
rect 11164 24052 11192 24092
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 10796 24024 11192 24052
rect 11882 24012 11888 24064
rect 11940 24012 11946 24064
rect 12434 24012 12440 24064
rect 12492 24012 12498 24064
rect 12526 24012 12532 24064
rect 12584 24012 12590 24064
rect 12894 24012 12900 24064
rect 12952 24012 12958 24064
rect 15120 24061 15148 24160
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 15252 24160 15485 24188
rect 15252 24148 15258 24160
rect 15473 24157 15485 24160
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24188 15623 24191
rect 17972 24188 18000 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 19061 24259 19119 24265
rect 19061 24225 19073 24259
rect 19107 24256 19119 24259
rect 19107 24228 21956 24256
rect 19107 24225 19119 24228
rect 19061 24219 19119 24225
rect 15611 24160 18000 24188
rect 18049 24191 18107 24197
rect 15611 24157 15623 24160
rect 15565 24151 15623 24157
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 18095 24160 18184 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 17586 24080 17592 24132
rect 17644 24120 17650 24132
rect 17782 24123 17840 24129
rect 17782 24120 17794 24123
rect 17644 24092 17794 24120
rect 17644 24080 17650 24092
rect 17782 24089 17794 24092
rect 17828 24089 17840 24123
rect 17782 24083 17840 24089
rect 18156 24064 18184 24160
rect 18432 24120 18460 24219
rect 21928 24200 21956 24228
rect 25314 24216 25320 24268
rect 25372 24256 25378 24268
rect 25409 24259 25467 24265
rect 25409 24256 25421 24259
rect 25372 24228 25421 24256
rect 25372 24216 25378 24228
rect 25409 24225 25421 24228
rect 25455 24225 25467 24259
rect 33502 24256 33508 24268
rect 25409 24219 25467 24225
rect 32876 24228 33508 24256
rect 18690 24148 18696 24200
rect 18748 24188 18754 24200
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 18748 24160 19809 24188
rect 18748 24148 18754 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 21910 24148 21916 24200
rect 21968 24148 21974 24200
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 26237 24191 26295 24197
rect 26237 24188 26249 24191
rect 23440 24160 26249 24188
rect 23440 24148 23446 24160
rect 26237 24157 26249 24160
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24188 28135 24191
rect 28166 24188 28172 24200
rect 28123 24160 28172 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 20254 24120 20260 24132
rect 18432 24092 20260 24120
rect 20254 24080 20260 24092
rect 20312 24080 20318 24132
rect 25225 24123 25283 24129
rect 25225 24089 25237 24123
rect 25271 24120 25283 24123
rect 26694 24120 26700 24132
rect 25271 24092 26700 24120
rect 25271 24089 25283 24092
rect 25225 24083 25283 24089
rect 26694 24080 26700 24092
rect 26752 24080 26758 24132
rect 27798 24080 27804 24132
rect 27856 24120 27862 24132
rect 27893 24123 27951 24129
rect 27893 24120 27905 24123
rect 27856 24092 27905 24120
rect 27856 24080 27862 24092
rect 27893 24089 27905 24092
rect 27939 24120 27951 24123
rect 28368 24120 28396 24151
rect 29178 24148 29184 24200
rect 29236 24148 29242 24200
rect 29641 24191 29699 24197
rect 29641 24157 29653 24191
rect 29687 24157 29699 24191
rect 29641 24151 29699 24157
rect 29825 24191 29883 24197
rect 29825 24157 29837 24191
rect 29871 24188 29883 24191
rect 29914 24188 29920 24200
rect 29871 24160 29920 24188
rect 29871 24157 29883 24160
rect 29825 24151 29883 24157
rect 27939 24092 28396 24120
rect 27939 24089 27951 24092
rect 27893 24083 27951 24089
rect 29454 24080 29460 24132
rect 29512 24120 29518 24132
rect 29656 24120 29684 24151
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 32306 24148 32312 24200
rect 32364 24188 32370 24200
rect 32677 24191 32735 24197
rect 32677 24188 32689 24191
rect 32364 24160 32689 24188
rect 32364 24148 32370 24160
rect 32677 24157 32689 24160
rect 32723 24157 32735 24191
rect 32677 24151 32735 24157
rect 32876 24129 32904 24228
rect 33502 24216 33508 24228
rect 33560 24216 33566 24268
rect 35529 24259 35587 24265
rect 35529 24225 35541 24259
rect 35575 24256 35587 24259
rect 37369 24259 37427 24265
rect 37369 24256 37381 24259
rect 35575 24228 37381 24256
rect 35575 24225 35587 24228
rect 35529 24219 35587 24225
rect 37369 24225 37381 24228
rect 37415 24256 37427 24259
rect 38654 24256 38660 24268
rect 37415 24228 38660 24256
rect 37415 24225 37427 24228
rect 37369 24219 37427 24225
rect 38654 24216 38660 24228
rect 38712 24256 38718 24268
rect 41049 24259 41107 24265
rect 41049 24256 41061 24259
rect 38712 24228 41061 24256
rect 38712 24216 38718 24228
rect 41049 24225 41061 24228
rect 41095 24225 41107 24259
rect 41049 24219 41107 24225
rect 41414 24216 41420 24268
rect 41472 24256 41478 24268
rect 42797 24259 42855 24265
rect 42797 24256 42809 24259
rect 41472 24228 42809 24256
rect 41472 24216 41478 24228
rect 42797 24225 42809 24228
rect 42843 24256 42855 24259
rect 42886 24256 42892 24268
rect 42843 24228 42892 24256
rect 42843 24225 42855 24228
rect 42797 24219 42855 24225
rect 42886 24216 42892 24228
rect 42944 24216 42950 24268
rect 44358 24216 44364 24268
rect 44416 24216 44422 24268
rect 44560 24256 44588 24352
rect 44637 24259 44695 24265
rect 44637 24256 44649 24259
rect 44560 24228 44649 24256
rect 44637 24225 44649 24228
rect 44683 24225 44695 24259
rect 44637 24219 44695 24225
rect 33042 24148 33048 24200
rect 33100 24148 33106 24200
rect 38746 24148 38752 24200
rect 38804 24148 38810 24200
rect 39390 24148 39396 24200
rect 39448 24148 39454 24200
rect 39577 24191 39635 24197
rect 39577 24157 39589 24191
rect 39623 24188 39635 24191
rect 40126 24188 40132 24200
rect 39623 24160 40132 24188
rect 39623 24157 39635 24160
rect 39577 24151 39635 24157
rect 40126 24148 40132 24160
rect 40184 24148 40190 24200
rect 40402 24188 40408 24200
rect 40236 24160 40408 24188
rect 32861 24123 32919 24129
rect 32861 24120 32873 24123
rect 29512 24092 29684 24120
rect 32692 24092 32873 24120
rect 29512 24080 29518 24092
rect 32692 24064 32720 24092
rect 32861 24089 32873 24092
rect 32907 24089 32919 24123
rect 32861 24083 32919 24089
rect 32953 24123 33011 24129
rect 32953 24089 32965 24123
rect 32999 24089 33011 24123
rect 32953 24083 33011 24089
rect 15105 24055 15163 24061
rect 15105 24021 15117 24055
rect 15151 24021 15163 24055
rect 15105 24015 15163 24021
rect 16666 24012 16672 24064
rect 16724 24012 16730 24064
rect 18138 24012 18144 24064
rect 18196 24012 18202 24064
rect 25317 24055 25375 24061
rect 25317 24021 25329 24055
rect 25363 24052 25375 24055
rect 25685 24055 25743 24061
rect 25685 24052 25697 24055
rect 25363 24024 25697 24052
rect 25363 24021 25375 24024
rect 25317 24015 25375 24021
rect 25685 24021 25697 24024
rect 25731 24021 25743 24055
rect 25685 24015 25743 24021
rect 27706 24012 27712 24064
rect 27764 24012 27770 24064
rect 28258 24012 28264 24064
rect 28316 24012 28322 24064
rect 32674 24012 32680 24064
rect 32732 24012 32738 24064
rect 32766 24012 32772 24064
rect 32824 24052 32830 24064
rect 32968 24052 32996 24083
rect 35802 24080 35808 24132
rect 35860 24080 35866 24132
rect 37918 24120 37924 24132
rect 37030 24092 37924 24120
rect 37918 24080 37924 24092
rect 37976 24080 37982 24132
rect 39408 24120 39436 24148
rect 40236 24129 40264 24160
rect 40402 24148 40408 24160
rect 40460 24148 40466 24200
rect 40221 24123 40279 24129
rect 39408 24092 39896 24120
rect 32824 24024 32996 24052
rect 33229 24055 33287 24061
rect 32824 24012 32830 24024
rect 33229 24021 33241 24055
rect 33275 24052 33287 24055
rect 33686 24052 33692 24064
rect 33275 24024 33692 24052
rect 33275 24021 33287 24024
rect 33229 24015 33287 24021
rect 33686 24012 33692 24024
rect 33744 24012 33750 24064
rect 35342 24012 35348 24064
rect 35400 24052 35406 24064
rect 36446 24052 36452 24064
rect 35400 24024 36452 24052
rect 35400 24012 35406 24024
rect 36446 24012 36452 24024
rect 36504 24012 36510 24064
rect 37274 24012 37280 24064
rect 37332 24012 37338 24064
rect 39206 24012 39212 24064
rect 39264 24052 39270 24064
rect 39868 24061 39896 24092
rect 40221 24089 40233 24123
rect 40267 24089 40279 24123
rect 40221 24083 40279 24089
rect 41325 24123 41383 24129
rect 41325 24089 41337 24123
rect 41371 24089 41383 24123
rect 42610 24120 42616 24132
rect 42550 24092 42616 24120
rect 41325 24083 41383 24089
rect 40034 24061 40040 24064
rect 39485 24055 39543 24061
rect 39485 24052 39497 24055
rect 39264 24024 39497 24052
rect 39264 24012 39270 24024
rect 39485 24021 39497 24024
rect 39531 24021 39543 24055
rect 39485 24015 39543 24021
rect 39853 24055 39911 24061
rect 39853 24021 39865 24055
rect 39899 24021 39911 24055
rect 39853 24015 39911 24021
rect 40021 24055 40040 24061
rect 40021 24021 40033 24055
rect 40021 24015 40040 24021
rect 40034 24012 40040 24015
rect 40092 24012 40098 24064
rect 41340 24052 41368 24083
rect 42610 24080 42616 24092
rect 42668 24080 42674 24132
rect 43714 24080 43720 24132
rect 43772 24080 43778 24132
rect 42058 24052 42064 24064
rect 41340 24024 42064 24052
rect 42058 24012 42064 24024
rect 42116 24012 42122 24064
rect 1104 23962 45172 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 45172 23962
rect 1104 23888 45172 23910
rect 10410 23808 10416 23860
rect 10468 23848 10474 23860
rect 10597 23851 10655 23857
rect 10597 23848 10609 23851
rect 10468 23820 10609 23848
rect 10468 23808 10474 23820
rect 10597 23817 10609 23820
rect 10643 23817 10655 23851
rect 10597 23811 10655 23817
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 10965 23851 11023 23857
rect 10965 23848 10977 23851
rect 10744 23820 10977 23848
rect 10744 23808 10750 23820
rect 10965 23817 10977 23820
rect 11011 23848 11023 23851
rect 11054 23848 11060 23860
rect 11011 23820 11060 23848
rect 11011 23817 11023 23820
rect 10965 23811 11023 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12253 23851 12311 23857
rect 12253 23848 12265 23851
rect 12124 23820 12265 23848
rect 12124 23808 12130 23820
rect 12253 23817 12265 23820
rect 12299 23817 12311 23851
rect 12526 23848 12532 23860
rect 12253 23811 12311 23817
rect 12406 23820 12532 23848
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23712 11115 23715
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11103 23684 12173 23712
rect 11103 23681 11115 23684
rect 11057 23675 11115 23681
rect 12161 23681 12173 23684
rect 12207 23712 12219 23715
rect 12406 23712 12434 23820
rect 12526 23808 12532 23820
rect 12584 23808 12590 23860
rect 12618 23808 12624 23860
rect 12676 23848 12682 23860
rect 13081 23851 13139 23857
rect 13081 23848 13093 23851
rect 12676 23820 13093 23848
rect 12676 23808 12682 23820
rect 13081 23817 13093 23820
rect 13127 23817 13139 23851
rect 16758 23848 16764 23860
rect 13081 23811 13139 23817
rect 14568 23820 16764 23848
rect 12713 23783 12771 23789
rect 12713 23749 12725 23783
rect 12759 23780 12771 23783
rect 14568 23780 14596 23820
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 16853 23851 16911 23857
rect 16853 23817 16865 23851
rect 16899 23848 16911 23851
rect 17218 23848 17224 23860
rect 16899 23820 17224 23848
rect 16899 23817 16911 23820
rect 16853 23811 16911 23817
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 17586 23808 17592 23860
rect 17644 23808 17650 23860
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 18417 23851 18475 23857
rect 18417 23848 18429 23851
rect 18196 23820 18429 23848
rect 18196 23808 18202 23820
rect 18417 23817 18429 23820
rect 18463 23848 18475 23851
rect 19426 23848 19432 23860
rect 18463 23820 19432 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 19426 23808 19432 23820
rect 19484 23848 19490 23860
rect 34790 23848 34796 23860
rect 19484 23820 19840 23848
rect 19484 23808 19490 23820
rect 12759 23752 14596 23780
rect 12759 23749 12771 23752
rect 12713 23743 12771 23749
rect 19812 23724 19840 23820
rect 25792 23820 34796 23848
rect 25792 23789 25820 23820
rect 34790 23808 34796 23820
rect 34848 23808 34854 23860
rect 35342 23848 35348 23860
rect 35176 23820 35348 23848
rect 24029 23783 24087 23789
rect 24029 23780 24041 23783
rect 19996 23752 24041 23780
rect 12207 23684 12434 23712
rect 12207 23681 12219 23684
rect 12161 23675 12219 23681
rect 10520 23576 10548 23675
rect 16666 23672 16672 23724
rect 16724 23712 16730 23724
rect 17405 23715 17463 23721
rect 17405 23712 17417 23715
rect 16724 23684 17417 23712
rect 16724 23672 16730 23684
rect 17405 23681 17417 23684
rect 17451 23681 17463 23715
rect 17405 23675 17463 23681
rect 17770 23672 17776 23724
rect 17828 23672 17834 23724
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19705 23715 19763 23721
rect 19705 23712 19717 23715
rect 19484 23684 19717 23712
rect 19484 23672 19490 23684
rect 19705 23681 19717 23684
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 19794 23672 19800 23724
rect 19852 23672 19858 23724
rect 19996 23712 20024 23752
rect 24029 23749 24041 23752
rect 24075 23749 24087 23783
rect 24029 23743 24087 23749
rect 25777 23783 25835 23789
rect 25777 23749 25789 23783
rect 25823 23749 25835 23783
rect 25777 23743 25835 23749
rect 20070 23721 20076 23724
rect 19904 23684 20024 23712
rect 11238 23604 11244 23656
rect 11296 23604 11302 23656
rect 11514 23604 11520 23656
rect 11572 23604 11578 23656
rect 12434 23604 12440 23656
rect 12492 23604 12498 23656
rect 12802 23604 12808 23656
rect 12860 23604 12866 23656
rect 13630 23604 13636 23656
rect 13688 23604 13694 23656
rect 14642 23604 14648 23656
rect 14700 23644 14706 23656
rect 19904 23644 19932 23684
rect 20064 23675 20076 23721
rect 20070 23672 20076 23675
rect 20128 23672 20134 23724
rect 22738 23721 22744 23724
rect 22732 23675 22744 23721
rect 22738 23672 22744 23675
rect 22796 23672 22802 23724
rect 14700 23616 19932 23644
rect 14700 23604 14706 23616
rect 21910 23604 21916 23656
rect 21968 23604 21974 23656
rect 22462 23604 22468 23656
rect 22520 23604 22526 23656
rect 12066 23576 12072 23588
rect 10520 23548 12072 23576
rect 12066 23536 12072 23548
rect 12124 23536 12130 23588
rect 8570 23468 8576 23520
rect 8628 23508 8634 23520
rect 9033 23511 9091 23517
rect 9033 23508 9045 23511
rect 8628 23480 9045 23508
rect 8628 23468 8634 23480
rect 9033 23477 9045 23480
rect 9079 23477 9091 23511
rect 12452 23508 12480 23604
rect 21177 23579 21235 23585
rect 21177 23545 21189 23579
rect 21223 23576 21235 23579
rect 21928 23576 21956 23604
rect 21223 23548 21956 23576
rect 24044 23576 24072 23743
rect 26510 23740 26516 23792
rect 26568 23780 26574 23792
rect 27338 23780 27344 23792
rect 26568 23752 27344 23780
rect 26568 23740 26574 23752
rect 27338 23740 27344 23752
rect 27396 23740 27402 23792
rect 28534 23780 28540 23792
rect 28474 23752 28540 23780
rect 28534 23740 28540 23752
rect 28592 23740 28598 23792
rect 32309 23783 32367 23789
rect 32309 23749 32321 23783
rect 32355 23780 32367 23783
rect 32674 23780 32680 23792
rect 32355 23752 32680 23780
rect 32355 23749 32367 23752
rect 32309 23743 32367 23749
rect 32674 23740 32680 23752
rect 32732 23740 32738 23792
rect 32766 23740 32772 23792
rect 32824 23780 32830 23792
rect 32861 23783 32919 23789
rect 32861 23780 32873 23783
rect 32824 23752 32873 23780
rect 32824 23740 32830 23752
rect 32861 23749 32873 23752
rect 32907 23749 32919 23783
rect 32861 23743 32919 23749
rect 33226 23740 33232 23792
rect 33284 23780 33290 23792
rect 33689 23783 33747 23789
rect 33689 23780 33701 23783
rect 33284 23752 33701 23780
rect 33284 23740 33290 23752
rect 33689 23749 33701 23752
rect 33735 23749 33747 23783
rect 33689 23743 33747 23749
rect 26970 23672 26976 23724
rect 27028 23672 27034 23724
rect 28460 23684 32076 23712
rect 27246 23604 27252 23656
rect 27304 23604 27310 23656
rect 27338 23604 27344 23656
rect 27396 23644 27402 23656
rect 28460 23644 28488 23684
rect 27396 23616 28488 23644
rect 28721 23647 28779 23653
rect 27396 23604 27402 23616
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 29362 23644 29368 23656
rect 28767 23616 29368 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 29362 23604 29368 23616
rect 29420 23604 29426 23656
rect 31938 23576 31944 23588
rect 24044 23548 27108 23576
rect 21223 23545 21235 23548
rect 21177 23539 21235 23545
rect 23382 23508 23388 23520
rect 12452 23480 23388 23508
rect 9033 23471 9091 23477
rect 23382 23468 23388 23480
rect 23440 23508 23446 23520
rect 23845 23511 23903 23517
rect 23845 23508 23857 23511
rect 23440 23480 23857 23508
rect 23440 23468 23446 23480
rect 23845 23477 23857 23480
rect 23891 23477 23903 23511
rect 23845 23471 23903 23477
rect 26234 23468 26240 23520
rect 26292 23468 26298 23520
rect 27080 23508 27108 23548
rect 28276 23548 31944 23576
rect 28276 23508 28304 23548
rect 31938 23536 31944 23548
rect 31996 23536 32002 23588
rect 27080 23480 28304 23508
rect 28810 23468 28816 23520
rect 28868 23468 28874 23520
rect 32048 23508 32076 23684
rect 32122 23672 32128 23724
rect 32180 23672 32186 23724
rect 32398 23672 32404 23724
rect 32456 23672 32462 23724
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23712 32551 23715
rect 33042 23712 33048 23724
rect 32539 23684 33048 23712
rect 32539 23681 32551 23684
rect 32493 23675 32551 23681
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 35176 23721 35204 23820
rect 35342 23808 35348 23820
rect 35400 23808 35406 23860
rect 35437 23851 35495 23857
rect 35437 23817 35449 23851
rect 35483 23848 35495 23851
rect 35802 23848 35808 23860
rect 35483 23820 35808 23848
rect 35483 23817 35495 23820
rect 35437 23811 35495 23817
rect 35802 23808 35808 23820
rect 35860 23808 35866 23860
rect 37918 23808 37924 23860
rect 37976 23848 37982 23860
rect 38197 23851 38255 23857
rect 38197 23848 38209 23851
rect 37976 23820 38209 23848
rect 37976 23808 37982 23820
rect 38197 23817 38209 23820
rect 38243 23848 38255 23851
rect 38562 23848 38568 23860
rect 38243 23820 38568 23848
rect 38243 23817 38255 23820
rect 38197 23811 38255 23817
rect 38562 23808 38568 23820
rect 38620 23808 38626 23860
rect 39206 23848 39212 23860
rect 39040 23820 39212 23848
rect 39040 23789 39068 23820
rect 39206 23808 39212 23820
rect 39264 23808 39270 23860
rect 40402 23808 40408 23860
rect 40460 23848 40466 23860
rect 40497 23851 40555 23857
rect 40497 23848 40509 23851
rect 40460 23820 40509 23848
rect 40460 23808 40466 23820
rect 40497 23817 40509 23820
rect 40543 23817 40555 23851
rect 40497 23811 40555 23817
rect 40678 23808 40684 23860
rect 40736 23848 40742 23860
rect 41325 23851 41383 23857
rect 41325 23848 41337 23851
rect 40736 23820 41337 23848
rect 40736 23808 40742 23820
rect 41325 23817 41337 23820
rect 41371 23817 41383 23851
rect 41325 23811 41383 23817
rect 41598 23808 41604 23860
rect 41656 23808 41662 23860
rect 41690 23808 41696 23860
rect 41748 23808 41754 23860
rect 42058 23808 42064 23860
rect 42116 23848 42122 23860
rect 42153 23851 42211 23857
rect 42153 23848 42165 23851
rect 42116 23820 42165 23848
rect 42116 23808 42122 23820
rect 42153 23817 42165 23820
rect 42199 23817 42211 23851
rect 42153 23811 42211 23817
rect 42794 23808 42800 23860
rect 42852 23808 42858 23860
rect 44542 23808 44548 23860
rect 44600 23808 44606 23860
rect 45278 23808 45284 23860
rect 45336 23808 45342 23860
rect 35253 23783 35311 23789
rect 35253 23749 35265 23783
rect 35299 23780 35311 23783
rect 37277 23783 37335 23789
rect 37277 23780 37289 23783
rect 35299 23752 35848 23780
rect 35299 23749 35311 23752
rect 35253 23743 35311 23749
rect 33597 23715 33655 23721
rect 33597 23712 33609 23715
rect 33428 23684 33609 23712
rect 33428 23656 33456 23684
rect 33597 23681 33609 23684
rect 33643 23681 33655 23715
rect 33597 23675 33655 23681
rect 35161 23715 35219 23721
rect 35161 23681 35173 23715
rect 35207 23681 35219 23715
rect 35161 23675 35219 23681
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 32766 23644 32772 23656
rect 32692 23616 32772 23644
rect 32692 23585 32720 23616
rect 32766 23604 32772 23616
rect 32824 23604 32830 23656
rect 33410 23604 33416 23656
rect 33468 23604 33474 23656
rect 32677 23579 32735 23585
rect 32677 23545 32689 23579
rect 32723 23545 32735 23579
rect 35360 23576 35388 23675
rect 35434 23672 35440 23724
rect 35492 23712 35498 23724
rect 35820 23721 35848 23752
rect 35912 23752 37289 23780
rect 35621 23715 35679 23721
rect 35621 23712 35633 23715
rect 35492 23684 35633 23712
rect 35492 23672 35498 23684
rect 35621 23681 35633 23684
rect 35667 23681 35679 23715
rect 35621 23675 35679 23681
rect 35713 23715 35771 23721
rect 35713 23681 35725 23715
rect 35759 23681 35771 23715
rect 35713 23675 35771 23681
rect 35805 23715 35863 23721
rect 35805 23681 35817 23715
rect 35851 23681 35863 23715
rect 35805 23675 35863 23681
rect 35728 23644 35756 23675
rect 35912 23644 35940 23752
rect 37277 23749 37289 23752
rect 37323 23749 37335 23783
rect 37277 23743 37335 23749
rect 39025 23783 39083 23789
rect 39025 23749 39037 23783
rect 39071 23749 39083 23783
rect 41616 23780 41644 23808
rect 39025 23743 39083 23749
rect 41064 23752 41644 23780
rect 35989 23715 36047 23721
rect 35989 23681 36001 23715
rect 36035 23712 36047 23715
rect 36081 23715 36139 23721
rect 36081 23712 36093 23715
rect 36035 23684 36093 23712
rect 36035 23681 36047 23684
rect 35989 23675 36047 23681
rect 36081 23681 36093 23684
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 38105 23715 38163 23721
rect 38105 23681 38117 23715
rect 38151 23681 38163 23715
rect 38105 23675 38163 23681
rect 36538 23644 36544 23656
rect 35728 23616 35940 23644
rect 36096 23616 36544 23644
rect 36096 23576 36124 23616
rect 36538 23604 36544 23616
rect 36596 23604 36602 23656
rect 37274 23604 37280 23656
rect 37332 23644 37338 23656
rect 37829 23647 37887 23653
rect 37829 23644 37841 23647
rect 37332 23616 37841 23644
rect 37332 23604 37338 23616
rect 37829 23613 37841 23616
rect 37875 23613 37887 23647
rect 37829 23607 37887 23613
rect 38120 23644 38148 23675
rect 38654 23672 38660 23724
rect 38712 23712 38718 23724
rect 41064 23721 41092 23752
rect 38749 23715 38807 23721
rect 38749 23712 38761 23715
rect 38712 23684 38761 23712
rect 38712 23672 38718 23684
rect 38749 23681 38761 23684
rect 38795 23681 38807 23715
rect 41049 23715 41107 23721
rect 38749 23675 38807 23681
rect 40144 23644 40172 23698
rect 41049 23681 41061 23715
rect 41095 23681 41107 23715
rect 41049 23675 41107 23681
rect 41233 23715 41291 23721
rect 41233 23681 41245 23715
rect 41279 23712 41291 23715
rect 41414 23712 41420 23724
rect 41279 23684 41420 23712
rect 41279 23681 41291 23684
rect 41233 23675 41291 23681
rect 41414 23672 41420 23684
rect 41472 23672 41478 23724
rect 41708 23712 41736 23808
rect 42610 23740 42616 23792
rect 42668 23780 42674 23792
rect 42668 23752 43102 23780
rect 42668 23740 42674 23752
rect 42061 23715 42119 23721
rect 42061 23712 42073 23715
rect 41708 23684 42073 23712
rect 42061 23681 42073 23684
rect 42107 23681 42119 23715
rect 42061 23675 42119 23681
rect 42245 23715 42303 23721
rect 42245 23681 42257 23715
rect 42291 23681 42303 23715
rect 42245 23675 42303 23681
rect 38120 23616 40172 23644
rect 38120 23576 38148 23616
rect 41782 23604 41788 23656
rect 41840 23644 41846 23656
rect 41877 23647 41935 23653
rect 41877 23644 41889 23647
rect 41840 23616 41889 23644
rect 41840 23604 41846 23616
rect 41877 23613 41889 23616
rect 41923 23613 41935 23647
rect 41877 23607 41935 23613
rect 35360 23548 36124 23576
rect 36372 23548 38148 23576
rect 32677 23539 32735 23545
rect 36372 23508 36400 23548
rect 40034 23536 40040 23588
rect 40092 23576 40098 23588
rect 40865 23579 40923 23585
rect 40865 23576 40877 23579
rect 40092 23548 40877 23576
rect 40092 23536 40098 23548
rect 40865 23545 40877 23548
rect 40911 23576 40923 23579
rect 42260 23576 42288 23675
rect 40911 23548 42288 23576
rect 40911 23545 40923 23548
rect 40865 23539 40923 23545
rect 32048 23480 36400 23508
rect 36446 23468 36452 23520
rect 36504 23468 36510 23520
rect 38562 23468 38568 23520
rect 38620 23508 38626 23520
rect 41598 23508 41604 23520
rect 38620 23480 41604 23508
rect 38620 23468 38626 23480
rect 41598 23468 41604 23480
rect 41656 23508 41662 23520
rect 42628 23508 42656 23740
rect 44560 23721 44588 23808
rect 44545 23715 44603 23721
rect 44545 23681 44557 23715
rect 44591 23681 44603 23715
rect 44545 23675 44603 23681
rect 44821 23715 44879 23721
rect 44821 23681 44833 23715
rect 44867 23712 44879 23715
rect 45296 23712 45324 23808
rect 44867 23684 45324 23712
rect 44867 23681 44879 23684
rect 44821 23675 44879 23681
rect 43254 23604 43260 23656
rect 43312 23644 43318 23656
rect 44269 23647 44327 23653
rect 44269 23644 44281 23647
rect 43312 23616 44281 23644
rect 43312 23604 43318 23616
rect 44269 23613 44281 23616
rect 44315 23613 44327 23647
rect 44269 23607 44327 23613
rect 41656 23480 42656 23508
rect 41656 23468 41662 23480
rect 44634 23468 44640 23520
rect 44692 23468 44698 23520
rect 1104 23418 45172 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 45172 23418
rect 1104 23344 45172 23366
rect 11054 23264 11060 23316
rect 11112 23264 11118 23316
rect 11333 23307 11391 23313
rect 11333 23273 11345 23307
rect 11379 23304 11391 23307
rect 11514 23304 11520 23316
rect 11379 23276 11520 23304
rect 11379 23273 11391 23276
rect 11333 23267 11391 23273
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 14461 23307 14519 23313
rect 14461 23273 14473 23307
rect 14507 23304 14519 23307
rect 17405 23307 17463 23313
rect 14507 23276 16712 23304
rect 14507 23273 14519 23276
rect 14461 23267 14519 23273
rect 16684 23236 16712 23276
rect 17405 23273 17417 23307
rect 17451 23304 17463 23307
rect 17770 23304 17776 23316
rect 17451 23276 17776 23304
rect 17451 23273 17463 23276
rect 17405 23267 17463 23273
rect 17770 23264 17776 23276
rect 17828 23264 17834 23316
rect 19613 23307 19671 23313
rect 19613 23273 19625 23307
rect 19659 23304 19671 23307
rect 20070 23304 20076 23316
rect 19659 23276 20076 23304
rect 19659 23273 19671 23276
rect 19613 23267 19671 23273
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 22370 23264 22376 23316
rect 22428 23264 22434 23316
rect 27246 23264 27252 23316
rect 27304 23304 27310 23316
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 27304 23276 27537 23304
rect 27304 23264 27310 23276
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 27525 23267 27583 23273
rect 28994 23264 29000 23316
rect 29052 23304 29058 23316
rect 29730 23304 29736 23316
rect 29052 23276 29736 23304
rect 29052 23264 29058 23276
rect 29730 23264 29736 23276
rect 29788 23264 29794 23316
rect 31389 23307 31447 23313
rect 29840 23276 30328 23304
rect 16684 23208 16804 23236
rect 16776 23180 16804 23208
rect 19794 23196 19800 23248
rect 19852 23236 19858 23248
rect 29365 23239 29423 23245
rect 19852 23208 21036 23236
rect 19852 23196 19858 23208
rect 9309 23171 9367 23177
rect 9309 23168 9321 23171
rect 8588 23140 9321 23168
rect 8588 23112 8616 23140
rect 9309 23137 9321 23140
rect 9355 23137 9367 23171
rect 9309 23131 9367 23137
rect 9585 23171 9643 23177
rect 9585 23137 9597 23171
rect 9631 23168 9643 23171
rect 10226 23168 10232 23180
rect 9631 23140 10232 23168
rect 9631 23137 9643 23140
rect 9585 23131 9643 23137
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 14645 23171 14703 23177
rect 14645 23137 14657 23171
rect 14691 23168 14703 23171
rect 14691 23140 16712 23168
rect 14691 23137 14703 23140
rect 14645 23131 14703 23137
rect 8570 23060 8576 23112
rect 8628 23060 8634 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9214 23100 9220 23112
rect 9171 23072 9220 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 10652 23072 10718 23100
rect 10652 23060 10658 23072
rect 11606 23060 11612 23112
rect 11664 23100 11670 23112
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 11664 23072 12725 23100
rect 11664 23060 11670 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 12989 23103 13047 23109
rect 12989 23100 13001 23103
rect 12952 23072 13001 23100
rect 12952 23060 12958 23072
rect 12989 23069 13001 23072
rect 13035 23069 13047 23103
rect 12989 23063 13047 23069
rect 16022 23060 16028 23112
rect 16080 23060 16086 23112
rect 16684 23100 16712 23140
rect 16758 23128 16764 23180
rect 16816 23128 16822 23180
rect 19978 23128 19984 23180
rect 20036 23168 20042 23180
rect 20441 23171 20499 23177
rect 20441 23168 20453 23171
rect 20036 23140 20453 23168
rect 20036 23128 20042 23140
rect 20441 23137 20453 23140
rect 20487 23137 20499 23171
rect 20441 23131 20499 23137
rect 16850 23100 16856 23112
rect 16684 23072 16856 23100
rect 16850 23060 16856 23072
rect 16908 23100 16914 23112
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 16908 23072 17509 23100
rect 16908 23060 16914 23072
rect 17497 23069 17509 23072
rect 17543 23100 17555 23103
rect 18138 23100 18144 23112
rect 17543 23072 18144 23100
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23100 19487 23103
rect 19475 23072 19932 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 12468 23035 12526 23041
rect 12468 23001 12480 23035
rect 12514 23032 12526 23035
rect 12514 23004 12848 23032
rect 12514 23001 12526 23004
rect 12468 22995 12526 23001
rect 8938 22924 8944 22976
rect 8996 22924 9002 22976
rect 12820 22973 12848 23004
rect 14090 22992 14096 23044
rect 14148 23032 14154 23044
rect 14185 23035 14243 23041
rect 14185 23032 14197 23035
rect 14148 23004 14197 23032
rect 14148 22992 14154 23004
rect 14185 23001 14197 23004
rect 14231 23032 14243 23035
rect 14826 23032 14832 23044
rect 14231 23004 14832 23032
rect 14231 23001 14243 23004
rect 14185 22995 14243 23001
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 14918 22992 14924 23044
rect 14976 22992 14982 23044
rect 17037 23035 17095 23041
rect 17037 23001 17049 23035
rect 17083 23032 17095 23035
rect 17218 23032 17224 23044
rect 17083 23004 17224 23032
rect 17083 23001 17095 23004
rect 17037 22995 17095 23001
rect 17218 22992 17224 23004
rect 17276 22992 17282 23044
rect 17764 23035 17822 23041
rect 17764 23001 17776 23035
rect 17810 23032 17822 23035
rect 17862 23032 17868 23044
rect 17810 23004 17868 23032
rect 17810 23001 17822 23004
rect 17764 22995 17822 23001
rect 17862 22992 17868 23004
rect 17920 22992 17926 23044
rect 19242 23032 19248 23044
rect 18800 23004 19248 23032
rect 12805 22967 12863 22973
rect 12805 22933 12817 22967
rect 12851 22933 12863 22967
rect 12805 22927 12863 22933
rect 16390 22924 16396 22976
rect 16448 22924 16454 22976
rect 16945 22967 17003 22973
rect 16945 22933 16957 22967
rect 16991 22964 17003 22967
rect 18800 22964 18828 23004
rect 19242 22992 19248 23004
rect 19300 22992 19306 23044
rect 16991 22936 18828 22964
rect 16991 22933 17003 22936
rect 16945 22927 17003 22933
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 19904 22973 19932 23072
rect 20254 23060 20260 23112
rect 20312 23060 20318 23112
rect 20714 23060 20720 23112
rect 20772 23060 20778 23112
rect 21008 23109 21036 23208
rect 28966 23208 29316 23236
rect 22462 23128 22468 23180
rect 22520 23128 22526 23180
rect 23014 23128 23020 23180
rect 23072 23128 23078 23180
rect 24946 23128 24952 23180
rect 25004 23168 25010 23180
rect 25866 23168 25872 23180
rect 25004 23140 25872 23168
rect 25004 23128 25010 23140
rect 25866 23128 25872 23140
rect 25924 23128 25930 23180
rect 28169 23171 28227 23177
rect 28169 23137 28181 23171
rect 28215 23168 28227 23171
rect 28810 23168 28816 23180
rect 28215 23140 28816 23168
rect 28215 23137 28227 23140
rect 28169 23131 28227 23137
rect 28810 23128 28816 23140
rect 28868 23128 28874 23180
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23100 21051 23103
rect 22480 23100 22508 23128
rect 21039 23072 22508 23100
rect 21039 23069 21051 23072
rect 20993 23063 21051 23069
rect 22646 23060 22652 23112
rect 22704 23100 22710 23112
rect 22925 23103 22983 23109
rect 22925 23100 22937 23103
rect 22704 23072 22937 23100
rect 22704 23060 22710 23072
rect 22925 23069 22937 23072
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 24673 23103 24731 23109
rect 24673 23069 24685 23103
rect 24719 23100 24731 23103
rect 24762 23100 24768 23112
rect 24719 23072 24768 23100
rect 24719 23069 24731 23072
rect 24673 23063 24731 23069
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 26234 23060 26240 23112
rect 26292 23100 26298 23112
rect 26292 23072 26358 23100
rect 26292 23060 26298 23072
rect 27706 23060 27712 23112
rect 27764 23060 27770 23112
rect 27801 23103 27859 23109
rect 27801 23069 27813 23103
rect 27847 23100 27859 23103
rect 28258 23100 28264 23112
rect 27847 23072 28264 23100
rect 27847 23069 27859 23072
rect 27801 23063 27859 23069
rect 28258 23060 28264 23072
rect 28316 23100 28322 23112
rect 28966 23100 28994 23208
rect 28316 23072 28994 23100
rect 28316 23060 28322 23072
rect 29086 23060 29092 23112
rect 29144 23060 29150 23112
rect 29288 23100 29316 23208
rect 29365 23205 29377 23239
rect 29411 23205 29423 23239
rect 29365 23199 29423 23205
rect 29380 23168 29408 23199
rect 29840 23168 29868 23276
rect 29917 23239 29975 23245
rect 29917 23205 29929 23239
rect 29963 23205 29975 23239
rect 29917 23199 29975 23205
rect 29380 23140 29868 23168
rect 29932 23168 29960 23199
rect 29932 23140 30236 23168
rect 30101 23103 30159 23109
rect 30101 23100 30113 23103
rect 29288 23072 30113 23100
rect 30101 23069 30113 23072
rect 30147 23069 30159 23103
rect 30101 23063 30159 23069
rect 21238 23035 21296 23041
rect 21238 23032 21250 23035
rect 20916 23004 21250 23032
rect 19889 22967 19947 22973
rect 19889 22933 19901 22967
rect 19935 22933 19947 22967
rect 19889 22927 19947 22933
rect 20349 22967 20407 22973
rect 20349 22933 20361 22967
rect 20395 22964 20407 22967
rect 20806 22964 20812 22976
rect 20395 22936 20812 22964
rect 20395 22933 20407 22936
rect 20349 22927 20407 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 20916 22973 20944 23004
rect 21238 23001 21250 23004
rect 21284 23001 21296 23035
rect 21238 22995 21296 23001
rect 22833 23035 22891 23041
rect 22833 23001 22845 23035
rect 22879 23032 22891 23035
rect 23400 23032 23428 23060
rect 22879 23004 23428 23032
rect 25225 23035 25283 23041
rect 22879 23001 22891 23004
rect 22833 22995 22891 23001
rect 25225 23001 25237 23035
rect 25271 23001 25283 23035
rect 25225 22995 25283 23001
rect 27893 23035 27951 23041
rect 27893 23001 27905 23035
rect 27939 23001 27951 23035
rect 27893 22995 27951 23001
rect 28031 23035 28089 23041
rect 28031 23001 28043 23035
rect 28077 23032 28089 23035
rect 28810 23032 28816 23044
rect 28077 23004 28816 23032
rect 28077 23001 28089 23004
rect 28031 22995 28089 23001
rect 20901 22967 20959 22973
rect 20901 22933 20913 22967
rect 20947 22933 20959 22967
rect 20901 22927 20959 22933
rect 22462 22924 22468 22976
rect 22520 22924 22526 22976
rect 24857 22967 24915 22973
rect 24857 22933 24869 22967
rect 24903 22964 24915 22967
rect 25240 22964 25268 22995
rect 24903 22936 25268 22964
rect 24903 22933 24915 22936
rect 24857 22927 24915 22933
rect 25498 22924 25504 22976
rect 25556 22964 25562 22976
rect 26697 22967 26755 22973
rect 26697 22964 26709 22967
rect 25556 22936 26709 22964
rect 25556 22924 25562 22936
rect 26697 22933 26709 22936
rect 26743 22964 26755 22967
rect 27798 22964 27804 22976
rect 26743 22936 27804 22964
rect 26743 22933 26755 22936
rect 26697 22927 26755 22933
rect 27798 22924 27804 22936
rect 27856 22924 27862 22976
rect 27908 22964 27936 22995
rect 28810 22992 28816 23004
rect 28868 22992 28874 23044
rect 28994 22992 29000 23044
rect 29052 23032 29058 23044
rect 29181 23035 29239 23041
rect 29181 23032 29193 23035
rect 29052 23004 29193 23032
rect 29052 22992 29058 23004
rect 29181 23001 29193 23004
rect 29227 23001 29239 23035
rect 29362 23032 29368 23044
rect 29323 23004 29368 23032
rect 29181 22995 29239 23001
rect 29362 22992 29368 23004
rect 29420 23032 29426 23044
rect 29549 23035 29607 23041
rect 29549 23032 29561 23035
rect 29420 23004 29561 23032
rect 29420 22992 29426 23004
rect 29549 23001 29561 23004
rect 29595 23001 29607 23035
rect 29549 22995 29607 23001
rect 28166 22964 28172 22976
rect 27908 22936 28172 22964
rect 28166 22924 28172 22936
rect 28224 22924 28230 22976
rect 29086 22924 29092 22976
rect 29144 22964 29150 22976
rect 29749 22967 29807 22973
rect 29749 22964 29761 22967
rect 29144 22936 29761 22964
rect 29144 22924 29150 22936
rect 29749 22933 29761 22936
rect 29795 22933 29807 22967
rect 30116 22964 30144 23063
rect 30208 23032 30236 23140
rect 30300 23112 30328 23276
rect 31389 23273 31401 23307
rect 31435 23304 31447 23307
rect 32122 23304 32128 23316
rect 31435 23276 32128 23304
rect 31435 23273 31447 23276
rect 31389 23267 31447 23273
rect 32122 23264 32128 23276
rect 32180 23264 32186 23316
rect 32398 23264 32404 23316
rect 32456 23264 32462 23316
rect 32677 23307 32735 23313
rect 32677 23273 32689 23307
rect 32723 23304 32735 23307
rect 33410 23304 33416 23316
rect 32723 23276 33416 23304
rect 32723 23273 32735 23276
rect 32677 23267 32735 23273
rect 33410 23264 33416 23276
rect 33468 23264 33474 23316
rect 36449 23307 36507 23313
rect 36449 23273 36461 23307
rect 36495 23304 36507 23307
rect 36538 23304 36544 23316
rect 36495 23276 36544 23304
rect 36495 23273 36507 23276
rect 36449 23267 36507 23273
rect 36538 23264 36544 23276
rect 36596 23264 36602 23316
rect 38654 23264 38660 23316
rect 38712 23304 38718 23316
rect 39209 23307 39267 23313
rect 39209 23304 39221 23307
rect 38712 23276 39221 23304
rect 38712 23264 38718 23276
rect 39209 23273 39221 23276
rect 39255 23273 39267 23307
rect 39209 23267 39267 23273
rect 31941 23239 31999 23245
rect 31941 23205 31953 23239
rect 31987 23236 31999 23239
rect 32416 23236 32444 23264
rect 31987 23208 32444 23236
rect 31987 23205 31999 23208
rect 31941 23199 31999 23205
rect 30926 23128 30932 23180
rect 30984 23128 30990 23180
rect 31726 23140 33088 23168
rect 30282 23060 30288 23112
rect 30340 23060 30346 23112
rect 30561 23103 30619 23109
rect 30561 23069 30573 23103
rect 30607 23069 30619 23103
rect 31021 23103 31079 23109
rect 31021 23100 31033 23103
rect 30561 23063 30619 23069
rect 30668 23072 31033 23100
rect 30374 23032 30380 23044
rect 30208 23004 30380 23032
rect 30374 22992 30380 23004
rect 30432 23032 30438 23044
rect 30576 23032 30604 23063
rect 30432 23004 30604 23032
rect 30432 22992 30438 23004
rect 30668 22964 30696 23072
rect 31021 23069 31033 23072
rect 31067 23069 31079 23103
rect 31021 23063 31079 23069
rect 30834 22992 30840 23044
rect 30892 23032 30898 23044
rect 31726 23032 31754 23140
rect 33060 23112 33088 23140
rect 33686 23128 33692 23180
rect 33744 23168 33750 23180
rect 34149 23171 34207 23177
rect 34149 23168 34161 23171
rect 33744 23140 34161 23168
rect 33744 23128 33750 23140
rect 34149 23137 34161 23140
rect 34195 23137 34207 23171
rect 39224 23168 39252 23267
rect 41782 23264 41788 23316
rect 41840 23304 41846 23316
rect 41969 23307 42027 23313
rect 41969 23304 41981 23307
rect 41840 23276 41981 23304
rect 41840 23264 41846 23276
rect 41969 23273 41981 23276
rect 42015 23273 42027 23307
rect 41969 23267 42027 23273
rect 43254 23264 43260 23316
rect 43312 23264 43318 23316
rect 40221 23171 40279 23177
rect 40221 23168 40233 23171
rect 39224 23140 40233 23168
rect 34149 23131 34207 23137
rect 40221 23137 40233 23140
rect 40267 23137 40279 23171
rect 40221 23131 40279 23137
rect 32582 23060 32588 23112
rect 32640 23060 32646 23112
rect 33042 23060 33048 23112
rect 33100 23060 33106 23112
rect 34425 23103 34483 23109
rect 34425 23069 34437 23103
rect 34471 23100 34483 23103
rect 34514 23100 34520 23112
rect 34471 23072 34520 23100
rect 34471 23069 34483 23072
rect 34425 23063 34483 23069
rect 34514 23060 34520 23072
rect 34572 23060 34578 23112
rect 36354 23060 36360 23112
rect 36412 23060 36418 23112
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 30892 23004 31754 23032
rect 30892 22992 30898 23004
rect 35986 22992 35992 23044
rect 36044 23032 36050 23044
rect 36556 23032 36584 23063
rect 41598 23060 41604 23112
rect 41656 23060 41662 23112
rect 43165 23103 43223 23109
rect 43165 23069 43177 23103
rect 43211 23100 43223 23103
rect 43530 23100 43536 23112
rect 43211 23072 43536 23100
rect 43211 23069 43223 23072
rect 43165 23063 43223 23069
rect 43530 23060 43536 23072
rect 43588 23060 43594 23112
rect 36044 23004 36584 23032
rect 36044 22992 36050 23004
rect 36630 22992 36636 23044
rect 36688 23032 36694 23044
rect 37921 23035 37979 23041
rect 37921 23032 37933 23035
rect 36688 23004 37933 23032
rect 36688 22992 36694 23004
rect 37921 23001 37933 23004
rect 37967 23032 37979 23035
rect 37967 23004 39344 23032
rect 37967 23001 37979 23004
rect 37921 22995 37979 23001
rect 30116 22936 30696 22964
rect 30745 22967 30803 22973
rect 29749 22927 29807 22933
rect 30745 22933 30757 22967
rect 30791 22964 30803 22967
rect 34606 22964 34612 22976
rect 30791 22936 34612 22964
rect 30791 22933 30803 22936
rect 30745 22927 30803 22933
rect 34606 22924 34612 22936
rect 34664 22924 34670 22976
rect 35618 22924 35624 22976
rect 35676 22964 35682 22976
rect 36538 22964 36544 22976
rect 35676 22936 36544 22964
rect 35676 22924 35682 22936
rect 36538 22924 36544 22936
rect 36596 22924 36602 22976
rect 39316 22964 39344 23004
rect 40494 22992 40500 23044
rect 40552 22992 40558 23044
rect 41892 23004 43116 23032
rect 41892 22964 41920 23004
rect 43088 22976 43116 23004
rect 39316 22936 41920 22964
rect 43070 22924 43076 22976
rect 43128 22924 43134 22976
rect 1104 22874 45172 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 45172 22874
rect 1104 22800 45172 22822
rect 9766 22720 9772 22772
rect 9824 22720 9830 22772
rect 12897 22763 12955 22769
rect 12897 22729 12909 22763
rect 12943 22760 12955 22763
rect 13630 22760 13636 22772
rect 12943 22732 13636 22760
rect 12943 22729 12955 22732
rect 12897 22723 12955 22729
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 14918 22720 14924 22772
rect 14976 22760 14982 22772
rect 15013 22763 15071 22769
rect 15013 22760 15025 22763
rect 14976 22732 15025 22760
rect 14976 22720 14982 22732
rect 15013 22729 15025 22732
rect 15059 22729 15071 22763
rect 15013 22723 15071 22729
rect 15654 22720 15660 22772
rect 15712 22760 15718 22772
rect 16390 22760 16396 22772
rect 15712 22732 16396 22760
rect 15712 22720 15718 22732
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 17862 22720 17868 22772
rect 17920 22720 17926 22772
rect 18414 22720 18420 22772
rect 18472 22760 18478 22772
rect 18509 22763 18567 22769
rect 18509 22760 18521 22763
rect 18472 22732 18521 22760
rect 18472 22720 18478 22732
rect 18509 22729 18521 22732
rect 18555 22729 18567 22763
rect 18509 22723 18567 22729
rect 18874 22720 18880 22772
rect 18932 22720 18938 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 21821 22763 21879 22769
rect 21821 22760 21833 22763
rect 20772 22732 21833 22760
rect 20772 22720 20778 22732
rect 21821 22729 21833 22732
rect 21867 22729 21879 22763
rect 21821 22723 21879 22729
rect 22189 22763 22247 22769
rect 22189 22729 22201 22763
rect 22235 22760 22247 22763
rect 22370 22760 22376 22772
rect 22235 22732 22376 22760
rect 22235 22729 22247 22732
rect 22189 22723 22247 22729
rect 22370 22720 22376 22732
rect 22428 22720 22434 22772
rect 22462 22720 22468 22772
rect 22520 22720 22526 22772
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 22833 22763 22891 22769
rect 22833 22760 22845 22763
rect 22796 22732 22845 22760
rect 22796 22720 22802 22732
rect 22833 22729 22845 22732
rect 22879 22729 22891 22763
rect 22833 22723 22891 22729
rect 24762 22720 24768 22772
rect 24820 22760 24826 22772
rect 25133 22763 25191 22769
rect 25133 22760 25145 22763
rect 24820 22732 25145 22760
rect 24820 22720 24826 22732
rect 25133 22729 25145 22732
rect 25179 22729 25191 22763
rect 25133 22723 25191 22729
rect 25498 22720 25504 22772
rect 25556 22720 25562 22772
rect 26510 22720 26516 22772
rect 26568 22720 26574 22772
rect 28166 22720 28172 22772
rect 28224 22720 28230 22772
rect 29362 22720 29368 22772
rect 29420 22760 29426 22772
rect 29457 22763 29515 22769
rect 29457 22760 29469 22763
rect 29420 22732 29469 22760
rect 29420 22720 29426 22732
rect 29457 22729 29469 22732
rect 29503 22729 29515 22763
rect 29457 22723 29515 22729
rect 29730 22720 29736 22772
rect 29788 22760 29794 22772
rect 29825 22763 29883 22769
rect 29825 22760 29837 22763
rect 29788 22732 29837 22760
rect 29788 22720 29794 22732
rect 29825 22729 29837 22732
rect 29871 22729 29883 22763
rect 29825 22723 29883 22729
rect 30282 22720 30288 22772
rect 30340 22720 30346 22772
rect 30374 22720 30380 22772
rect 30432 22720 30438 22772
rect 30561 22763 30619 22769
rect 30561 22729 30573 22763
rect 30607 22760 30619 22763
rect 30926 22760 30932 22772
rect 30607 22732 30932 22760
rect 30607 22729 30619 22732
rect 30561 22723 30619 22729
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 32582 22720 32588 22772
rect 32640 22760 32646 22772
rect 33873 22763 33931 22769
rect 33873 22760 33885 22763
rect 32640 22732 33885 22760
rect 32640 22720 32646 22732
rect 33873 22729 33885 22732
rect 33919 22729 33931 22763
rect 33873 22723 33931 22729
rect 34072 22732 35940 22760
rect 8570 22692 8576 22704
rect 8036 22664 8576 22692
rect 8036 22633 8064 22664
rect 8570 22652 8576 22664
rect 8628 22652 8634 22704
rect 10962 22692 10968 22704
rect 9522 22664 10968 22692
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 11784 22695 11842 22701
rect 11784 22661 11796 22695
rect 11830 22692 11842 22695
rect 11882 22692 11888 22704
rect 11830 22664 11888 22692
rect 11830 22661 11842 22664
rect 11784 22655 11842 22661
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 13538 22652 13544 22704
rect 13596 22692 13602 22704
rect 14369 22695 14427 22701
rect 14369 22692 14381 22695
rect 13596 22664 14381 22692
rect 13596 22652 13602 22664
rect 14369 22661 14381 22664
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 15749 22695 15807 22701
rect 15749 22661 15761 22695
rect 15795 22692 15807 22695
rect 16574 22692 16580 22704
rect 15795 22664 16580 22692
rect 15795 22661 15807 22664
rect 15749 22655 15807 22661
rect 16574 22652 16580 22664
rect 16632 22652 16638 22704
rect 18601 22695 18659 22701
rect 18601 22661 18613 22695
rect 18647 22692 18659 22695
rect 18647 22664 18828 22692
rect 18647 22661 18659 22664
rect 18601 22655 18659 22661
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 11606 22624 11612 22636
rect 11563 22596 11612 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 11606 22584 11612 22596
rect 11664 22584 11670 22636
rect 14458 22584 14464 22636
rect 14516 22584 14522 22636
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22624 15255 22627
rect 15243 22596 15332 22624
rect 15243 22593 15255 22596
rect 15197 22587 15255 22593
rect 8297 22559 8355 22565
rect 8297 22525 8309 22559
rect 8343 22556 8355 22559
rect 8938 22556 8944 22568
rect 8343 22528 8944 22556
rect 8343 22525 8355 22528
rect 8297 22519 8355 22525
rect 8938 22516 8944 22528
rect 8996 22516 9002 22568
rect 15304 22497 15332 22596
rect 18046 22584 18052 22636
rect 18104 22584 18110 22636
rect 15378 22516 15384 22568
rect 15436 22556 15442 22568
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 15436 22528 15853 22556
rect 15436 22516 15442 22528
rect 15841 22525 15853 22528
rect 15887 22525 15899 22559
rect 15841 22519 15899 22525
rect 17218 22516 17224 22568
rect 17276 22516 17282 22568
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18693 22559 18751 22565
rect 18693 22556 18705 22559
rect 17920 22528 18705 22556
rect 17920 22516 17926 22528
rect 18693 22525 18705 22528
rect 18739 22525 18751 22559
rect 18800 22556 18828 22664
rect 18892 22624 18920 22720
rect 20533 22695 20591 22701
rect 20533 22661 20545 22695
rect 20579 22692 20591 22695
rect 20622 22692 20628 22704
rect 20579 22664 20628 22692
rect 20579 22661 20591 22664
rect 20533 22655 20591 22661
rect 20622 22652 20628 22664
rect 20680 22652 20686 22704
rect 19521 22627 19579 22633
rect 19521 22624 19533 22627
rect 18892 22596 19533 22624
rect 19521 22593 19533 22596
rect 19567 22593 19579 22627
rect 22480 22624 22508 22720
rect 24673 22695 24731 22701
rect 24673 22692 24685 22695
rect 23400 22664 24685 22692
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 22480 22596 22661 22624
rect 19521 22587 19579 22593
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 18800 22528 22232 22556
rect 18693 22519 18751 22525
rect 15289 22491 15347 22497
rect 14292 22460 14504 22488
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 12158 22420 12164 22432
rect 11848 22392 12164 22420
rect 11848 22380 11854 22392
rect 12158 22380 12164 22392
rect 12216 22420 12222 22432
rect 14292 22420 14320 22460
rect 12216 22392 14320 22420
rect 14476 22420 14504 22460
rect 15289 22457 15301 22491
rect 15335 22457 15347 22491
rect 15289 22451 15347 22457
rect 16592 22460 18276 22488
rect 16592 22420 16620 22460
rect 14476 22392 16620 22420
rect 12216 22380 12222 22392
rect 16666 22380 16672 22432
rect 16724 22380 16730 22432
rect 18138 22380 18144 22432
rect 18196 22380 18202 22432
rect 18248 22420 18276 22460
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 18969 22491 19027 22497
rect 18969 22488 18981 22491
rect 18472 22460 18981 22488
rect 18472 22448 18478 22460
rect 18969 22457 18981 22460
rect 19015 22457 19027 22491
rect 22204 22488 22232 22528
rect 22278 22516 22284 22568
rect 22336 22516 22342 22568
rect 22462 22516 22468 22568
rect 22520 22556 22526 22568
rect 23014 22556 23020 22568
rect 22520 22528 23020 22556
rect 22520 22516 22526 22528
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 23106 22516 23112 22568
rect 23164 22516 23170 22568
rect 22370 22488 22376 22500
rect 18969 22451 19027 22457
rect 19076 22460 22094 22488
rect 22204 22460 22376 22488
rect 19076 22420 19104 22460
rect 18248 22392 19104 22420
rect 19978 22380 19984 22432
rect 20036 22420 20042 22432
rect 20257 22423 20315 22429
rect 20257 22420 20269 22423
rect 20036 22392 20269 22420
rect 20036 22380 20042 22392
rect 20257 22389 20269 22392
rect 20303 22389 20315 22423
rect 22066 22420 22094 22460
rect 22370 22448 22376 22460
rect 22428 22448 22434 22500
rect 23400 22420 23428 22664
rect 24673 22661 24685 22664
rect 24719 22661 24731 22695
rect 24673 22655 24731 22661
rect 25041 22695 25099 22701
rect 25041 22661 25053 22695
rect 25087 22692 25099 22695
rect 26528 22692 26556 22720
rect 25087 22664 26556 22692
rect 28184 22692 28212 22720
rect 28184 22664 30144 22692
rect 25087 22661 25099 22664
rect 25041 22655 25099 22661
rect 24118 22584 24124 22636
rect 24176 22624 24182 22636
rect 24397 22627 24455 22633
rect 24397 22624 24409 22627
rect 24176 22596 24409 22624
rect 24176 22584 24182 22596
rect 24397 22593 24409 22596
rect 24443 22624 24455 22627
rect 25056 22624 25084 22655
rect 24443 22596 25084 22624
rect 24443 22593 24455 22596
rect 24397 22587 24455 22593
rect 25314 22584 25320 22636
rect 25372 22624 25378 22636
rect 25372 22596 25728 22624
rect 25372 22584 25378 22596
rect 25700 22565 25728 22596
rect 27798 22584 27804 22636
rect 27856 22624 27862 22636
rect 28166 22624 28172 22636
rect 27856 22596 28172 22624
rect 27856 22584 27862 22596
rect 28166 22584 28172 22596
rect 28224 22624 28230 22636
rect 28629 22627 28687 22633
rect 28629 22624 28641 22627
rect 28224 22596 28641 22624
rect 28224 22584 28230 22596
rect 28629 22593 28641 22596
rect 28675 22593 28687 22627
rect 28629 22587 28687 22593
rect 28813 22627 28871 22633
rect 28813 22593 28825 22627
rect 28859 22624 28871 22627
rect 28902 22624 28908 22636
rect 28859 22596 28908 22624
rect 28859 22593 28871 22596
rect 28813 22587 28871 22593
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29089 22627 29147 22633
rect 29089 22593 29101 22627
rect 29135 22624 29147 22627
rect 29178 22624 29184 22636
rect 29135 22596 29184 22624
rect 29135 22593 29147 22596
rect 29089 22587 29147 22593
rect 29178 22584 29184 22596
rect 29236 22584 29242 22636
rect 29270 22584 29276 22636
rect 29328 22624 29334 22636
rect 29365 22627 29423 22633
rect 29365 22624 29377 22627
rect 29328 22596 29377 22624
rect 29328 22584 29334 22596
rect 29365 22593 29377 22596
rect 29411 22593 29423 22627
rect 29365 22587 29423 22593
rect 29641 22627 29699 22633
rect 29641 22593 29653 22627
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 23753 22559 23811 22565
rect 23753 22525 23765 22559
rect 23799 22556 23811 22559
rect 25593 22559 25651 22565
rect 25593 22556 25605 22559
rect 23799 22528 25605 22556
rect 23799 22525 23811 22528
rect 23753 22519 23811 22525
rect 25593 22525 25605 22528
rect 25639 22525 25651 22559
rect 25593 22519 25651 22525
rect 25685 22559 25743 22565
rect 25685 22525 25697 22559
rect 25731 22556 25743 22559
rect 27522 22556 27528 22568
rect 25731 22528 27528 22556
rect 25731 22525 25743 22528
rect 25685 22519 25743 22525
rect 27522 22516 27528 22528
rect 27580 22516 27586 22568
rect 28920 22556 28948 22584
rect 29656 22556 29684 22587
rect 28920 22528 29684 22556
rect 30116 22556 30144 22664
rect 30193 22627 30251 22633
rect 30193 22593 30205 22627
rect 30239 22624 30251 22627
rect 30300 22624 30328 22720
rect 30392 22633 30420 22720
rect 33042 22652 33048 22704
rect 33100 22652 33106 22704
rect 30239 22596 30328 22624
rect 30377 22627 30435 22633
rect 30239 22593 30251 22596
rect 30193 22587 30251 22593
rect 30377 22593 30389 22627
rect 30423 22593 30435 22627
rect 33888 22624 33916 22723
rect 33965 22627 34023 22633
rect 33965 22624 33977 22627
rect 33888 22596 33977 22624
rect 30377 22587 30435 22593
rect 33965 22593 33977 22596
rect 34011 22593 34023 22627
rect 33965 22587 34023 22593
rect 30116 22528 32076 22556
rect 28534 22448 28540 22500
rect 28592 22488 28598 22500
rect 30834 22488 30840 22500
rect 28592 22460 30840 22488
rect 28592 22448 28598 22460
rect 30834 22448 30840 22460
rect 30892 22448 30898 22500
rect 22066 22392 23428 22420
rect 20257 22383 20315 22389
rect 24302 22380 24308 22432
rect 24360 22380 24366 22432
rect 29273 22423 29331 22429
rect 29273 22389 29285 22423
rect 29319 22420 29331 22423
rect 29638 22420 29644 22432
rect 29319 22392 29644 22420
rect 29319 22389 29331 22392
rect 29273 22383 29331 22389
rect 29638 22380 29644 22392
rect 29696 22380 29702 22432
rect 32048 22420 32076 22528
rect 32122 22516 32128 22568
rect 32180 22516 32186 22568
rect 32401 22559 32459 22565
rect 32401 22525 32413 22559
rect 32447 22556 32459 22559
rect 32766 22556 32772 22568
rect 32447 22528 32772 22556
rect 32447 22525 32459 22528
rect 32401 22519 32459 22525
rect 32766 22516 32772 22528
rect 32824 22516 32830 22568
rect 34072 22556 34100 22732
rect 34606 22652 34612 22704
rect 34664 22692 34670 22704
rect 35342 22692 35348 22704
rect 34664 22664 35348 22692
rect 34664 22652 34670 22664
rect 35342 22652 35348 22664
rect 35400 22652 35406 22704
rect 35618 22652 35624 22704
rect 35676 22692 35682 22704
rect 35912 22701 35940 22732
rect 36354 22720 36360 22772
rect 36412 22720 36418 22772
rect 40494 22720 40500 22772
rect 40552 22720 40558 22772
rect 35759 22695 35817 22701
rect 35759 22692 35771 22695
rect 35676 22664 35771 22692
rect 35676 22652 35682 22664
rect 35759 22661 35771 22664
rect 35805 22661 35817 22695
rect 35759 22655 35817 22661
rect 35897 22695 35955 22701
rect 35897 22661 35909 22695
rect 35943 22661 35955 22695
rect 35897 22655 35955 22661
rect 35989 22695 36047 22701
rect 35989 22661 36001 22695
rect 36035 22692 36047 22695
rect 36372 22692 36400 22720
rect 36035 22664 36400 22692
rect 36035 22661 36047 22664
rect 35989 22655 36047 22661
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22593 35219 22627
rect 36004 22624 36032 22655
rect 35161 22587 35219 22593
rect 35866 22596 36032 22624
rect 33980 22528 34100 22556
rect 35176 22556 35204 22587
rect 35434 22556 35440 22568
rect 35176 22528 35440 22556
rect 33980 22420 34008 22528
rect 35434 22516 35440 22528
rect 35492 22516 35498 22568
rect 35618 22516 35624 22568
rect 35676 22516 35682 22568
rect 35529 22491 35587 22497
rect 35529 22457 35541 22491
rect 35575 22488 35587 22491
rect 35866 22488 35894 22596
rect 36078 22584 36084 22636
rect 36136 22584 36142 22636
rect 40129 22627 40187 22633
rect 40129 22593 40141 22627
rect 40175 22593 40187 22627
rect 40129 22587 40187 22593
rect 36357 22559 36415 22565
rect 36357 22556 36369 22559
rect 35575 22460 35894 22488
rect 36050 22528 36369 22556
rect 35575 22457 35587 22460
rect 35529 22451 35587 22457
rect 32048 22392 34008 22420
rect 34054 22380 34060 22432
rect 34112 22380 34118 22432
rect 35618 22380 35624 22432
rect 35676 22420 35682 22432
rect 36050 22420 36078 22528
rect 36357 22525 36369 22528
rect 36403 22525 36415 22559
rect 36357 22519 36415 22525
rect 37001 22559 37059 22565
rect 37001 22525 37013 22559
rect 37047 22556 37059 22559
rect 37734 22556 37740 22568
rect 37047 22528 37740 22556
rect 37047 22525 37059 22528
rect 37001 22519 37059 22525
rect 36170 22448 36176 22500
rect 36228 22488 36234 22500
rect 37016 22488 37044 22519
rect 37734 22516 37740 22528
rect 37792 22516 37798 22568
rect 40034 22516 40040 22568
rect 40092 22516 40098 22568
rect 36228 22460 37044 22488
rect 40144 22488 40172 22587
rect 40512 22565 40540 22720
rect 41693 22627 41751 22633
rect 41693 22593 41705 22627
rect 41739 22624 41751 22627
rect 41782 22624 41788 22636
rect 41739 22596 41788 22624
rect 41739 22593 41751 22596
rect 41693 22587 41751 22593
rect 41782 22584 41788 22596
rect 41840 22584 41846 22636
rect 40497 22559 40555 22565
rect 40497 22525 40509 22559
rect 40543 22525 40555 22559
rect 40497 22519 40555 22525
rect 41049 22491 41107 22497
rect 41049 22488 41061 22491
rect 40144 22460 41061 22488
rect 36228 22448 36234 22460
rect 41049 22457 41061 22460
rect 41095 22457 41107 22491
rect 41049 22451 41107 22457
rect 35676 22392 36078 22420
rect 35676 22380 35682 22392
rect 36262 22380 36268 22432
rect 36320 22380 36326 22432
rect 1104 22330 45172 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 45172 22330
rect 1104 22256 45172 22278
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 14884 22188 16252 22216
rect 14884 22176 14890 22188
rect 16224 22148 16252 22188
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17589 22219 17647 22225
rect 17589 22216 17601 22219
rect 16632 22188 17601 22216
rect 16632 22176 16638 22188
rect 17589 22185 17601 22188
rect 17635 22185 17647 22219
rect 17589 22179 17647 22185
rect 18046 22176 18052 22228
rect 18104 22216 18110 22228
rect 18141 22219 18199 22225
rect 18141 22216 18153 22219
rect 18104 22188 18153 22216
rect 18104 22176 18110 22188
rect 18141 22185 18153 22188
rect 18187 22185 18199 22219
rect 20530 22216 20536 22228
rect 18141 22179 18199 22185
rect 18248 22188 20536 22216
rect 18248 22148 18276 22188
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 20625 22219 20683 22225
rect 20625 22185 20637 22219
rect 20671 22216 20683 22219
rect 25314 22216 25320 22228
rect 20671 22188 21404 22216
rect 20671 22185 20683 22188
rect 20625 22179 20683 22185
rect 16224 22120 18276 22148
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17402 22080 17408 22092
rect 16908 22052 17408 22080
rect 16908 22040 16914 22052
rect 17402 22040 17408 22052
rect 17460 22080 17466 22092
rect 21376 22089 21404 22188
rect 25056 22188 25320 22216
rect 23216 22120 24716 22148
rect 19245 22083 19303 22089
rect 19245 22080 19257 22083
rect 17460 22052 19257 22080
rect 17460 22040 17466 22052
rect 19245 22049 19257 22052
rect 19291 22049 19303 22083
rect 19245 22043 19303 22049
rect 21361 22083 21419 22089
rect 21361 22049 21373 22083
rect 21407 22080 21419 22083
rect 23106 22080 23112 22092
rect 21407 22052 23112 22080
rect 21407 22049 21419 22052
rect 21361 22043 21419 22049
rect 23106 22040 23112 22052
rect 23164 22040 23170 22092
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 14642 22012 14648 22024
rect 13587 21984 14648 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 22012 15347 22015
rect 16868 22012 16896 22040
rect 23216 22024 23244 22120
rect 24688 22080 24716 22120
rect 24762 22108 24768 22160
rect 24820 22148 24826 22160
rect 25056 22148 25084 22188
rect 25314 22176 25320 22188
rect 25372 22176 25378 22228
rect 29086 22176 29092 22228
rect 29144 22176 29150 22228
rect 31938 22176 31944 22228
rect 31996 22216 32002 22228
rect 34146 22216 34152 22228
rect 31996 22188 34152 22216
rect 31996 22176 32002 22188
rect 34146 22176 34152 22188
rect 34204 22176 34210 22228
rect 35986 22216 35992 22228
rect 35866 22188 35992 22216
rect 24820 22120 25084 22148
rect 24820 22108 24826 22120
rect 25056 22089 25084 22120
rect 28166 22108 28172 22160
rect 28224 22148 28230 22160
rect 29362 22148 29368 22160
rect 28224 22120 29368 22148
rect 28224 22108 28230 22120
rect 24857 22083 24915 22089
rect 24857 22080 24869 22083
rect 24688 22052 24869 22080
rect 24857 22049 24869 22052
rect 24903 22049 24915 22083
rect 24857 22043 24915 22049
rect 25041 22083 25099 22089
rect 25041 22049 25053 22083
rect 25087 22080 25099 22083
rect 25087 22052 25121 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 25866 22040 25872 22092
rect 25924 22040 25930 22092
rect 15335 21984 16896 22012
rect 16945 22015 17003 22021
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 16945 21981 16957 22015
rect 16991 21981 17003 22015
rect 16945 21975 17003 21981
rect 15556 21947 15614 21953
rect 15556 21913 15568 21947
rect 15602 21944 15614 21947
rect 15746 21944 15752 21956
rect 15602 21916 15752 21944
rect 15602 21913 15614 21916
rect 15556 21907 15614 21913
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 13078 21836 13084 21888
rect 13136 21876 13142 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 13136 21848 13369 21876
rect 13136 21836 13142 21848
rect 13357 21845 13369 21848
rect 13403 21845 13415 21879
rect 13357 21839 13415 21845
rect 16669 21879 16727 21885
rect 16669 21845 16681 21879
rect 16715 21876 16727 21879
rect 16960 21876 16988 21975
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 18196 21984 18705 22012
rect 18196 21972 18202 21984
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 23198 22012 23204 22024
rect 22428 21984 23204 22012
rect 22428 21972 22434 21984
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 21981 23811 22015
rect 29012 22012 29040 22120
rect 29362 22108 29368 22120
rect 29420 22108 29426 22160
rect 30101 22151 30159 22157
rect 30101 22117 30113 22151
rect 30147 22148 30159 22151
rect 34241 22151 34299 22157
rect 30147 22120 31708 22148
rect 30147 22117 30159 22120
rect 30101 22111 30159 22117
rect 29638 22040 29644 22092
rect 29696 22040 29702 22092
rect 29089 22015 29147 22021
rect 29089 22012 29101 22015
rect 29012 21984 29101 22012
rect 23753 21975 23811 21981
rect 29089 21981 29101 21984
rect 29135 21981 29147 22015
rect 29089 21975 29147 21981
rect 19058 21904 19064 21956
rect 19116 21944 19122 21956
rect 19490 21947 19548 21953
rect 19490 21944 19502 21947
rect 19116 21916 19502 21944
rect 19116 21904 19122 21916
rect 19490 21913 19502 21916
rect 19536 21913 19548 21947
rect 19490 21907 19548 21913
rect 16715 21848 16988 21876
rect 16715 21845 16727 21848
rect 16669 21839 16727 21845
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 20717 21879 20775 21885
rect 20717 21876 20729 21879
rect 19300 21848 20729 21876
rect 19300 21836 19306 21848
rect 20717 21845 20729 21848
rect 20763 21845 20775 21879
rect 20717 21839 20775 21845
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 23658 21876 23664 21888
rect 23615 21848 23664 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 23768 21876 23796 21975
rect 29270 21972 29276 22024
rect 29328 21972 29334 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 21981 29791 22015
rect 31680 22012 31708 22120
rect 34241 22117 34253 22151
rect 34287 22148 34299 22151
rect 34287 22120 34652 22148
rect 34287 22117 34299 22120
rect 34241 22111 34299 22117
rect 34624 22080 34652 22120
rect 35866 22080 35894 22188
rect 35986 22176 35992 22188
rect 36044 22176 36050 22228
rect 36262 22225 36268 22228
rect 36252 22219 36268 22225
rect 36252 22185 36264 22219
rect 36252 22179 36268 22185
rect 36262 22176 36268 22179
rect 36320 22176 36326 22228
rect 37734 22176 37740 22228
rect 37792 22176 37798 22228
rect 34624 22052 34928 22080
rect 34900 22021 34928 22052
rect 35176 22052 35894 22080
rect 35989 22083 36047 22089
rect 35176 22021 35204 22052
rect 35989 22049 36001 22083
rect 36035 22080 36047 22083
rect 37829 22083 37887 22089
rect 37829 22080 37841 22083
rect 36035 22052 37841 22080
rect 36035 22049 36047 22052
rect 35989 22043 36047 22049
rect 37829 22049 37841 22052
rect 37875 22080 37887 22083
rect 38194 22080 38200 22092
rect 37875 22052 38200 22080
rect 37875 22049 37887 22052
rect 37829 22043 37887 22049
rect 38194 22040 38200 22052
rect 38252 22080 38258 22092
rect 38746 22080 38752 22092
rect 38252 22052 38752 22080
rect 38252 22040 38258 22052
rect 38746 22040 38752 22052
rect 38804 22040 38810 22092
rect 39577 22083 39635 22089
rect 39577 22049 39589 22083
rect 39623 22080 39635 22083
rect 39758 22080 39764 22092
rect 39623 22052 39764 22080
rect 39623 22049 39635 22052
rect 39577 22043 39635 22049
rect 39758 22040 39764 22052
rect 39816 22080 39822 22092
rect 40405 22083 40463 22089
rect 40405 22080 40417 22083
rect 39816 22052 40417 22080
rect 39816 22040 39822 22052
rect 40405 22049 40417 22052
rect 40451 22049 40463 22083
rect 40405 22043 40463 22049
rect 33873 22015 33931 22021
rect 33873 22012 33885 22015
rect 31680 21984 33885 22012
rect 29733 21975 29791 21981
rect 33873 21981 33885 21984
rect 33919 22012 33931 22015
rect 34333 22015 34391 22021
rect 34333 22012 34345 22015
rect 33919 21984 34345 22012
rect 33919 21981 33931 21984
rect 33873 21975 33931 21981
rect 34333 21981 34345 21984
rect 34379 21981 34391 22015
rect 34517 22015 34575 22021
rect 34517 22012 34529 22015
rect 34333 21975 34391 21981
rect 34440 21984 34529 22012
rect 26142 21904 26148 21956
rect 26200 21904 26206 21956
rect 27706 21944 27712 21956
rect 27370 21916 27712 21944
rect 27706 21904 27712 21916
rect 27764 21944 27770 21956
rect 28534 21944 28540 21956
rect 27764 21916 28540 21944
rect 27764 21904 27770 21916
rect 28534 21904 28540 21916
rect 28592 21904 28598 21956
rect 28813 21947 28871 21953
rect 28813 21913 28825 21947
rect 28859 21913 28871 21947
rect 28813 21907 28871 21913
rect 24397 21879 24455 21885
rect 24397 21876 24409 21879
rect 23768 21848 24409 21876
rect 24397 21845 24409 21848
rect 24443 21845 24455 21879
rect 24397 21839 24455 21845
rect 24765 21879 24823 21885
rect 24765 21845 24777 21879
rect 24811 21876 24823 21879
rect 25130 21876 25136 21888
rect 24811 21848 25136 21876
rect 24811 21845 24823 21848
rect 24765 21839 24823 21845
rect 25130 21836 25136 21848
rect 25188 21836 25194 21888
rect 27614 21836 27620 21888
rect 27672 21836 27678 21888
rect 28828 21876 28856 21907
rect 28902 21904 28908 21956
rect 28960 21944 28966 21956
rect 28997 21947 29055 21953
rect 28997 21944 29009 21947
rect 28960 21916 29009 21944
rect 28960 21904 28966 21916
rect 28997 21913 29009 21916
rect 29043 21913 29055 21947
rect 28997 21907 29055 21913
rect 29288 21876 29316 21972
rect 29748 21888 29776 21975
rect 34054 21904 34060 21956
rect 34112 21944 34118 21956
rect 34440 21944 34468 21984
rect 34517 21981 34529 21984
rect 34563 21981 34575 22015
rect 34517 21975 34575 21981
rect 34701 22015 34759 22021
rect 34701 21981 34713 22015
rect 34747 21981 34759 22015
rect 34701 21975 34759 21981
rect 34885 22015 34943 22021
rect 34885 21981 34897 22015
rect 34931 22012 34943 22015
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 34931 21984 35173 22012
rect 34931 21981 34943 21984
rect 34885 21975 34943 21981
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 34716 21944 34744 21975
rect 35342 21972 35348 22024
rect 35400 21972 35406 22024
rect 35434 21972 35440 22024
rect 35492 21972 35498 22024
rect 35526 21972 35532 22024
rect 35584 21972 35590 22024
rect 34112 21916 34468 21944
rect 34532 21916 34744 21944
rect 34793 21947 34851 21953
rect 34112 21904 34118 21916
rect 28828 21848 29316 21876
rect 29730 21836 29736 21888
rect 29788 21836 29794 21888
rect 34532 21885 34560 21916
rect 34793 21913 34805 21947
rect 34839 21944 34851 21947
rect 35452 21944 35480 21972
rect 34839 21916 35480 21944
rect 37490 21916 38056 21944
rect 34839 21913 34851 21916
rect 34793 21907 34851 21913
rect 34517 21879 34575 21885
rect 34517 21845 34529 21879
rect 34563 21845 34575 21879
rect 34517 21839 34575 21845
rect 35802 21836 35808 21888
rect 35860 21836 35866 21888
rect 38028 21876 38056 21916
rect 38102 21904 38108 21956
rect 38160 21904 38166 21956
rect 38562 21944 38568 21956
rect 38212 21916 38568 21944
rect 38212 21876 38240 21916
rect 38562 21904 38568 21916
rect 38620 21904 38626 21956
rect 38028 21848 38240 21876
rect 39850 21836 39856 21888
rect 39908 21836 39914 21888
rect 1104 21786 45172 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 45172 21786
rect 1104 21712 45172 21734
rect 14458 21632 14464 21684
rect 14516 21672 14522 21684
rect 14553 21675 14611 21681
rect 14553 21672 14565 21675
rect 14516 21644 14565 21672
rect 14516 21632 14522 21644
rect 14553 21641 14565 21644
rect 14599 21641 14611 21675
rect 14553 21635 14611 21641
rect 13078 21564 13084 21616
rect 13136 21564 13142 21616
rect 14568 21604 14596 21635
rect 14642 21632 14648 21684
rect 14700 21632 14706 21684
rect 15746 21632 15752 21684
rect 15804 21632 15810 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16632 21644 17049 21672
rect 16632 21632 16638 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 19058 21632 19064 21684
rect 19116 21632 19122 21684
rect 19242 21632 19248 21684
rect 19300 21672 19306 21684
rect 19521 21675 19579 21681
rect 19521 21672 19533 21675
rect 19300 21644 19533 21672
rect 19300 21632 19306 21644
rect 19521 21641 19533 21644
rect 19567 21641 19579 21675
rect 19521 21635 19579 21641
rect 23198 21632 23204 21684
rect 23256 21632 23262 21684
rect 25130 21632 25136 21684
rect 25188 21632 25194 21684
rect 26142 21632 26148 21684
rect 26200 21632 26206 21684
rect 26973 21675 27031 21681
rect 26973 21641 26985 21675
rect 27019 21641 27031 21675
rect 26973 21635 27031 21641
rect 15013 21607 15071 21613
rect 15013 21604 15025 21607
rect 14568 21576 15025 21604
rect 15013 21573 15025 21576
rect 15059 21573 15071 21607
rect 16022 21604 16028 21616
rect 15013 21567 15071 21573
rect 15111 21576 16028 21604
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 15111 21536 15139 21576
rect 16022 21564 16028 21576
rect 16080 21564 16086 21616
rect 21805 21576 23428 21604
rect 14240 21508 15139 21536
rect 15933 21539 15991 21545
rect 14240 21496 14246 21508
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16666 21536 16672 21548
rect 15979 21508 16672 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 18877 21539 18935 21545
rect 16816 21508 17356 21536
rect 16816 21496 16822 21508
rect 11974 21428 11980 21480
rect 12032 21468 12038 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12032 21440 12817 21468
rect 12032 21428 12038 21440
rect 12805 21437 12817 21440
rect 12851 21437 12863 21471
rect 12805 21431 12863 21437
rect 12820 21332 12848 21431
rect 15102 21428 15108 21480
rect 15160 21428 15166 21480
rect 15194 21428 15200 21480
rect 15252 21428 15258 21480
rect 17328 21477 17356 21508
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 21361 21539 21419 21545
rect 18923 21508 19196 21536
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 17313 21471 17371 21477
rect 17313 21437 17325 21471
rect 17359 21468 17371 21471
rect 17862 21468 17868 21480
rect 17359 21440 17868 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 17144 21400 17172 21431
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18601 21471 18659 21477
rect 18601 21468 18613 21471
rect 18380 21440 18613 21468
rect 18380 21428 18386 21440
rect 18601 21437 18613 21440
rect 18647 21437 18659 21471
rect 18601 21431 18659 21437
rect 19168 21409 19196 21508
rect 21361 21505 21373 21539
rect 21407 21536 21419 21539
rect 21450 21536 21456 21548
rect 21407 21508 21456 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 21805 21545 21833 21576
rect 21805 21539 21879 21545
rect 21805 21512 21833 21539
rect 21821 21505 21833 21512
rect 21867 21505 21879 21539
rect 22077 21539 22135 21545
rect 22077 21536 22089 21539
rect 21821 21499 21879 21505
rect 21928 21508 22089 21536
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 19613 21471 19671 21477
rect 19613 21468 19625 21471
rect 19300 21440 19625 21468
rect 19300 21428 19306 21440
rect 19613 21437 19625 21440
rect 19659 21437 19671 21471
rect 19613 21431 19671 21437
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21468 19855 21471
rect 19978 21468 19984 21480
rect 19843 21440 19984 21468
rect 19843 21437 19855 21440
rect 19797 21431 19855 21437
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 21928 21468 21956 21508
rect 22077 21505 22089 21508
rect 22123 21505 22135 21539
rect 22077 21499 22135 21505
rect 23400 21480 23428 21576
rect 25148 21536 25176 21632
rect 26329 21539 26387 21545
rect 21836 21440 21956 21468
rect 19153 21403 19211 21409
rect 17144 21372 19104 21400
rect 13538 21332 13544 21344
rect 12820 21304 13544 21332
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 16669 21335 16727 21341
rect 16669 21301 16681 21335
rect 16715 21332 16727 21335
rect 17218 21332 17224 21344
rect 16715 21304 17224 21332
rect 16715 21301 16727 21304
rect 16669 21295 16727 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18046 21292 18052 21344
rect 18104 21292 18110 21344
rect 19076 21332 19104 21372
rect 19153 21369 19165 21403
rect 19199 21369 19211 21403
rect 19153 21363 19211 21369
rect 21545 21403 21603 21409
rect 21545 21369 21557 21403
rect 21591 21400 21603 21403
rect 21836 21400 21864 21440
rect 23382 21428 23388 21480
rect 23440 21428 23446 21480
rect 23658 21428 23664 21480
rect 23716 21428 23722 21480
rect 24302 21428 24308 21480
rect 24360 21468 24366 21480
rect 24780 21468 24808 21522
rect 25148 21508 25820 21536
rect 25130 21468 25136 21480
rect 24360 21440 25136 21468
rect 24360 21428 24366 21440
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 25225 21471 25283 21477
rect 25225 21437 25237 21471
rect 25271 21437 25283 21471
rect 25225 21431 25283 21437
rect 25240 21400 25268 21431
rect 21591 21372 21864 21400
rect 24688 21372 25268 21400
rect 25792 21400 25820 21508
rect 26329 21505 26341 21539
rect 26375 21536 26387 21539
rect 26988 21536 27016 21635
rect 28074 21632 28080 21684
rect 28132 21672 28138 21684
rect 29730 21672 29736 21684
rect 28132 21644 29736 21672
rect 28132 21632 28138 21644
rect 29730 21632 29736 21644
rect 29788 21632 29794 21684
rect 35342 21632 35348 21684
rect 35400 21632 35406 21684
rect 36078 21632 36084 21684
rect 36136 21632 36142 21684
rect 36357 21675 36415 21681
rect 36357 21641 36369 21675
rect 36403 21672 36415 21675
rect 36446 21672 36452 21684
rect 36403 21644 36452 21672
rect 36403 21641 36415 21644
rect 36357 21635 36415 21641
rect 36446 21632 36452 21644
rect 36504 21632 36510 21684
rect 38102 21632 38108 21684
rect 38160 21672 38166 21684
rect 38197 21675 38255 21681
rect 38197 21672 38209 21675
rect 38160 21644 38209 21672
rect 38160 21632 38166 21644
rect 38197 21641 38209 21644
rect 38243 21641 38255 21675
rect 38197 21635 38255 21641
rect 39850 21632 39856 21684
rect 39908 21632 39914 21684
rect 27341 21607 27399 21613
rect 27341 21573 27353 21607
rect 27387 21604 27399 21607
rect 27614 21604 27620 21616
rect 27387 21576 27620 21604
rect 27387 21573 27399 21576
rect 27341 21567 27399 21573
rect 27614 21564 27620 21576
rect 27672 21604 27678 21616
rect 27672 21576 28396 21604
rect 27672 21564 27678 21576
rect 28368 21545 28396 21576
rect 29270 21564 29276 21616
rect 29328 21604 29334 21616
rect 29328 21576 29868 21604
rect 29328 21564 29334 21576
rect 26375 21508 27016 21536
rect 28077 21539 28135 21545
rect 26375 21505 26387 21508
rect 26329 21499 26387 21505
rect 28077 21505 28089 21539
rect 28123 21505 28135 21539
rect 28077 21499 28135 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 28905 21539 28963 21545
rect 28905 21536 28917 21539
rect 28399 21508 28917 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 28905 21505 28917 21508
rect 28951 21505 28963 21539
rect 28905 21499 28963 21505
rect 29549 21539 29607 21545
rect 29549 21505 29561 21539
rect 29595 21536 29607 21539
rect 29638 21536 29644 21548
rect 29595 21508 29644 21536
rect 29595 21505 29607 21508
rect 29549 21499 29607 21505
rect 25869 21471 25927 21477
rect 25869 21437 25881 21471
rect 25915 21468 25927 21471
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 25915 21440 27445 21468
rect 25915 21437 25927 21440
rect 25869 21431 25927 21437
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 27522 21428 27528 21480
rect 27580 21428 27586 21480
rect 28092 21400 28120 21499
rect 29638 21496 29644 21508
rect 29696 21496 29702 21548
rect 29840 21545 29868 21576
rect 35526 21564 35532 21616
rect 35584 21604 35590 21616
rect 35897 21607 35955 21613
rect 35584 21576 35848 21604
rect 35584 21564 35590 21576
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21505 29883 21539
rect 29825 21499 29883 21505
rect 35253 21539 35311 21545
rect 35253 21505 35265 21539
rect 35299 21505 35311 21539
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 35253 21499 35311 21505
rect 35360 21508 35449 21536
rect 28166 21428 28172 21480
rect 28224 21428 28230 21480
rect 28997 21471 29055 21477
rect 28997 21437 29009 21471
rect 29043 21468 29055 21471
rect 29365 21471 29423 21477
rect 29365 21468 29377 21471
rect 29043 21440 29377 21468
rect 29043 21437 29055 21440
rect 28997 21431 29055 21437
rect 29365 21437 29377 21440
rect 29411 21437 29423 21471
rect 29365 21431 29423 21437
rect 28902 21400 28908 21412
rect 25792 21372 28908 21400
rect 21591 21369 21603 21372
rect 21545 21363 21603 21369
rect 23290 21332 23296 21344
rect 19076 21304 23296 21332
rect 23290 21292 23296 21304
rect 23348 21332 23354 21344
rect 24688 21332 24716 21372
rect 28902 21360 28908 21372
rect 28960 21360 28966 21412
rect 29273 21403 29331 21409
rect 29273 21369 29285 21403
rect 29319 21400 29331 21403
rect 35268 21400 35296 21499
rect 35360 21468 35388 21508
rect 35437 21505 35449 21508
rect 35483 21505 35495 21539
rect 35437 21499 35495 21505
rect 35710 21496 35716 21548
rect 35768 21496 35774 21548
rect 35820 21536 35848 21576
rect 35897 21573 35909 21607
rect 35943 21604 35955 21607
rect 35943 21576 36308 21604
rect 35943 21573 35955 21576
rect 35897 21567 35955 21573
rect 35989 21539 36047 21545
rect 35989 21536 36001 21539
rect 35820 21508 36001 21536
rect 35989 21505 36001 21508
rect 36035 21505 36047 21539
rect 35989 21499 36047 21505
rect 36078 21496 36084 21548
rect 36136 21496 36142 21548
rect 36280 21545 36308 21576
rect 36173 21539 36231 21545
rect 36173 21505 36185 21539
rect 36219 21505 36231 21539
rect 36173 21499 36231 21505
rect 36265 21539 36323 21545
rect 36265 21505 36277 21539
rect 36311 21505 36323 21539
rect 36265 21499 36323 21505
rect 35526 21468 35532 21480
rect 35360 21440 35532 21468
rect 35526 21428 35532 21440
rect 35584 21468 35590 21480
rect 36096 21468 36124 21496
rect 35584 21440 36124 21468
rect 35584 21428 35590 21440
rect 29319 21372 35296 21400
rect 29319 21369 29331 21372
rect 29273 21363 29331 21369
rect 23348 21304 24716 21332
rect 23348 21292 23354 21304
rect 28074 21292 28080 21344
rect 28132 21292 28138 21344
rect 28537 21335 28595 21341
rect 28537 21301 28549 21335
rect 28583 21332 28595 21335
rect 28994 21332 29000 21344
rect 28583 21304 29000 21332
rect 28583 21301 28595 21304
rect 28537 21295 28595 21301
rect 28994 21292 29000 21304
rect 29052 21292 29058 21344
rect 35268 21332 35296 21372
rect 35434 21360 35440 21412
rect 35492 21400 35498 21412
rect 36188 21400 36216 21499
rect 36446 21496 36452 21548
rect 36504 21496 36510 21548
rect 39301 21539 39359 21545
rect 39301 21505 39313 21539
rect 39347 21536 39359 21539
rect 39868 21536 39896 21632
rect 39347 21508 39896 21536
rect 39347 21505 39359 21508
rect 39301 21499 39359 21505
rect 38841 21471 38899 21477
rect 38841 21437 38853 21471
rect 38887 21468 38899 21471
rect 38887 21440 38976 21468
rect 38887 21437 38899 21440
rect 38841 21431 38899 21437
rect 38948 21409 38976 21440
rect 39390 21428 39396 21480
rect 39448 21428 39454 21480
rect 35492 21372 36216 21400
rect 38933 21403 38991 21409
rect 35492 21360 35498 21372
rect 38933 21369 38945 21403
rect 38979 21369 38991 21403
rect 38933 21363 38991 21369
rect 35710 21332 35716 21344
rect 35268 21304 35716 21332
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 38838 21292 38844 21344
rect 38896 21332 38902 21344
rect 39482 21332 39488 21344
rect 38896 21304 39488 21332
rect 38896 21292 38902 21304
rect 39482 21292 39488 21304
rect 39540 21292 39546 21344
rect 1104 21242 45172 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 45172 21242
rect 1104 21168 45172 21190
rect 11241 21131 11299 21137
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11422 21128 11428 21140
rect 11287 21100 11428 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 11422 21088 11428 21100
rect 11480 21088 11486 21140
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13814 21128 13820 21140
rect 13771 21100 13820 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 18690 21088 18696 21140
rect 18748 21088 18754 21140
rect 22373 21131 22431 21137
rect 22373 21097 22385 21131
rect 22419 21128 22431 21131
rect 23290 21128 23296 21140
rect 22419 21100 23296 21128
rect 22419 21097 22431 21100
rect 22373 21091 22431 21097
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 24762 21128 24768 21140
rect 23584 21100 24768 21128
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20992 9551 20995
rect 9539 20964 12020 20992
rect 9539 20961 9551 20964
rect 9493 20955 9551 20961
rect 11992 20936 12020 20964
rect 23198 20952 23204 21004
rect 23256 20992 23262 21004
rect 23584 21001 23612 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 32306 21088 32312 21140
rect 32364 21088 32370 21140
rect 39301 21131 39359 21137
rect 39301 21097 39313 21131
rect 39347 21128 39359 21131
rect 39390 21128 39396 21140
rect 39347 21100 39396 21128
rect 39347 21097 39359 21100
rect 39301 21091 39359 21097
rect 23293 20995 23351 21001
rect 23293 20992 23305 20995
rect 23256 20964 23305 20992
rect 23256 20952 23262 20964
rect 23293 20961 23305 20964
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23569 20995 23627 21001
rect 23569 20961 23581 20995
rect 23615 20992 23627 20995
rect 23658 20992 23664 21004
rect 23615 20964 23664 20992
rect 23615 20961 23627 20964
rect 23569 20955 23627 20961
rect 23658 20952 23664 20964
rect 23716 20952 23722 21004
rect 25130 20952 25136 21004
rect 25188 20992 25194 21004
rect 25188 20964 25912 20992
rect 25188 20952 25194 20964
rect 10778 20884 10784 20936
rect 10836 20924 10842 20936
rect 10836 20896 10902 20924
rect 10836 20884 10842 20896
rect 11974 20884 11980 20936
rect 12032 20884 12038 20936
rect 14090 20884 14096 20936
rect 14148 20884 14154 20936
rect 14182 20884 14188 20936
rect 14240 20884 14246 20936
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 17402 20924 17408 20936
rect 17359 20896 17408 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 20714 20884 20720 20936
rect 20772 20884 20778 20936
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 23382 20924 23388 20936
rect 21039 20896 23388 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 23382 20884 23388 20896
rect 23440 20924 23446 20936
rect 24394 20924 24400 20936
rect 23440 20896 24400 20924
rect 23440 20884 23446 20896
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 9766 20816 9772 20868
rect 9824 20816 9830 20868
rect 12250 20816 12256 20868
rect 12308 20816 12314 20868
rect 14200 20856 14228 20884
rect 13478 20828 14228 20856
rect 17580 20859 17638 20865
rect 17580 20825 17592 20859
rect 17626 20856 17638 20859
rect 17770 20856 17776 20868
rect 17626 20828 17776 20856
rect 17626 20825 17638 20828
rect 17580 20819 17638 20825
rect 17770 20816 17776 20828
rect 17828 20816 17834 20868
rect 21238 20859 21296 20865
rect 21238 20856 21250 20859
rect 20916 20828 21250 20856
rect 14458 20748 14464 20800
rect 14516 20788 14522 20800
rect 20916 20797 20944 20828
rect 21238 20825 21250 20828
rect 21284 20825 21296 20859
rect 21238 20819 21296 20825
rect 23845 20859 23903 20865
rect 23845 20825 23857 20859
rect 23891 20856 23903 20859
rect 23891 20828 24624 20856
rect 23891 20825 23903 20828
rect 23845 20819 23903 20825
rect 14737 20791 14795 20797
rect 14737 20788 14749 20791
rect 14516 20760 14749 20788
rect 14516 20748 14522 20760
rect 14737 20757 14749 20760
rect 14783 20757 14795 20791
rect 14737 20751 14795 20757
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 22738 20748 22744 20800
rect 22796 20748 22802 20800
rect 23750 20748 23756 20800
rect 23808 20748 23814 20800
rect 24210 20748 24216 20800
rect 24268 20748 24274 20800
rect 24596 20788 24624 20828
rect 24670 20816 24676 20868
rect 24728 20816 24734 20868
rect 25884 20856 25912 20964
rect 32030 20952 32036 21004
rect 32088 20952 32094 21004
rect 39117 20995 39175 21001
rect 39117 20961 39129 20995
rect 39163 20992 39175 20995
rect 39316 20992 39344 21091
rect 39390 21088 39396 21100
rect 39448 21088 39454 21140
rect 39163 20964 39344 20992
rect 39163 20961 39175 20964
rect 39117 20955 39175 20961
rect 39482 20952 39488 21004
rect 39540 20952 39546 21004
rect 31941 20927 31999 20933
rect 31941 20893 31953 20927
rect 31987 20924 31999 20927
rect 32398 20924 32404 20936
rect 31987 20896 32404 20924
rect 31987 20893 31999 20896
rect 31941 20887 31999 20893
rect 32398 20884 32404 20896
rect 32456 20884 32462 20936
rect 35526 20884 35532 20936
rect 35584 20884 35590 20936
rect 35710 20884 35716 20936
rect 35768 20884 35774 20936
rect 36446 20884 36452 20936
rect 36504 20884 36510 20936
rect 38930 20884 38936 20936
rect 38988 20884 38994 20936
rect 39209 20927 39267 20933
rect 39209 20893 39221 20927
rect 39255 20924 39267 20927
rect 39393 20927 39451 20933
rect 39255 20896 39344 20924
rect 39255 20893 39267 20896
rect 39209 20887 39267 20893
rect 25958 20856 25964 20868
rect 25884 20842 25964 20856
rect 25898 20828 25964 20842
rect 25958 20816 25964 20828
rect 26016 20856 26022 20868
rect 27706 20856 27712 20868
rect 26016 20828 27712 20856
rect 26016 20816 26022 20828
rect 27706 20816 27712 20828
rect 27764 20816 27770 20868
rect 35434 20816 35440 20868
rect 35492 20856 35498 20868
rect 35621 20859 35679 20865
rect 35621 20856 35633 20859
rect 35492 20828 35633 20856
rect 35492 20816 35498 20828
rect 35621 20825 35633 20828
rect 35667 20856 35679 20859
rect 36464 20856 36492 20884
rect 35667 20828 36492 20856
rect 35667 20825 35679 20828
rect 35621 20819 35679 20825
rect 39316 20800 39344 20896
rect 39393 20893 39405 20927
rect 39439 20924 39451 20927
rect 39500 20924 39528 20952
rect 39439 20896 39528 20924
rect 39439 20893 39451 20896
rect 39393 20887 39451 20893
rect 26145 20791 26203 20797
rect 26145 20788 26157 20791
rect 24596 20760 26157 20788
rect 26145 20757 26157 20760
rect 26191 20788 26203 20791
rect 28074 20788 28080 20800
rect 26191 20760 28080 20788
rect 26191 20757 26203 20760
rect 26145 20751 26203 20757
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 38746 20748 38752 20800
rect 38804 20748 38810 20800
rect 39298 20748 39304 20800
rect 39356 20748 39362 20800
rect 1104 20698 45172 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 45172 20698
rect 1104 20624 45172 20646
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 10045 20587 10103 20593
rect 10045 20584 10057 20587
rect 9824 20556 10057 20584
rect 9824 20544 9830 20556
rect 10045 20553 10057 20556
rect 10091 20553 10103 20587
rect 10045 20547 10103 20553
rect 10505 20587 10563 20593
rect 10505 20553 10517 20587
rect 10551 20553 10563 20587
rect 10505 20547 10563 20553
rect 10873 20587 10931 20593
rect 10873 20553 10885 20587
rect 10919 20584 10931 20587
rect 11422 20584 11428 20596
rect 10919 20556 11428 20584
rect 10919 20553 10931 20556
rect 10873 20547 10931 20553
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20448 10287 20451
rect 10520 20448 10548 20547
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 13872 20556 14381 20584
rect 13872 20544 13878 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14369 20547 14427 20553
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 12124 20488 12173 20516
rect 12124 20476 12130 20488
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12161 20479 12219 20485
rect 10275 20420 10548 20448
rect 11885 20451 11943 20457
rect 10275 20417 10287 20420
rect 10229 20411 10287 20417
rect 11885 20417 11897 20451
rect 11931 20448 11943 20451
rect 15565 20451 15623 20457
rect 11931 20420 12434 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11238 20380 11244 20392
rect 11195 20352 11244 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 10980 20312 11008 20343
rect 11238 20340 11244 20352
rect 11296 20340 11302 20392
rect 12250 20340 12256 20392
rect 12308 20340 12314 20392
rect 11882 20312 11888 20324
rect 10980 20284 11888 20312
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 12069 20315 12127 20321
rect 12069 20281 12081 20315
rect 12115 20312 12127 20315
rect 12268 20312 12296 20340
rect 12115 20284 12296 20312
rect 12406 20312 12434 20420
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 15672 20448 15700 20547
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15988 20556 16037 20584
rect 15988 20544 15994 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 17770 20544 17776 20596
rect 17828 20544 17834 20596
rect 18046 20544 18052 20596
rect 18104 20544 18110 20596
rect 18417 20587 18475 20593
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 18690 20584 18696 20596
rect 18463 20556 18696 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 18690 20544 18696 20556
rect 18748 20544 18754 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20901 20587 20959 20593
rect 20901 20584 20913 20587
rect 20772 20556 20913 20584
rect 20772 20544 20778 20556
rect 20901 20553 20913 20556
rect 20947 20553 20959 20587
rect 20901 20547 20959 20553
rect 21266 20544 21272 20596
rect 21324 20584 21330 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 21324 20556 21373 20584
rect 21324 20544 21330 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 21450 20544 21456 20596
rect 21508 20584 21514 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21508 20556 21833 20584
rect 21508 20544 21514 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 22189 20587 22247 20593
rect 22189 20553 22201 20587
rect 22235 20584 22247 20587
rect 22738 20584 22744 20596
rect 22235 20556 22744 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 23750 20544 23756 20596
rect 23808 20584 23814 20596
rect 24029 20587 24087 20593
rect 24029 20584 24041 20587
rect 23808 20556 24041 20584
rect 23808 20544 23814 20556
rect 24029 20553 24041 20556
rect 24075 20553 24087 20587
rect 24029 20547 24087 20553
rect 24210 20544 24216 20596
rect 24268 20544 24274 20596
rect 24305 20587 24363 20593
rect 24305 20553 24317 20587
rect 24351 20584 24363 20587
rect 24670 20584 24676 20596
rect 24351 20556 24676 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 31941 20587 31999 20593
rect 31941 20553 31953 20587
rect 31987 20584 31999 20587
rect 32030 20584 32036 20596
rect 31987 20556 32036 20584
rect 31987 20553 31999 20556
rect 31941 20547 31999 20553
rect 32030 20544 32036 20556
rect 32088 20544 32094 20596
rect 32490 20544 32496 20596
rect 32548 20584 32554 20596
rect 32769 20587 32827 20593
rect 32769 20584 32781 20587
rect 32548 20556 32781 20584
rect 32548 20544 32554 20556
rect 32769 20553 32781 20556
rect 32815 20553 32827 20587
rect 32769 20547 32827 20553
rect 38746 20544 38752 20596
rect 38804 20544 38810 20596
rect 38838 20544 38844 20596
rect 38896 20544 38902 20596
rect 39482 20544 39488 20596
rect 39540 20584 39546 20596
rect 39945 20587 40003 20593
rect 39945 20584 39957 20587
rect 39540 20556 39957 20584
rect 39540 20544 39546 20556
rect 39945 20553 39957 20556
rect 39991 20553 40003 20587
rect 39945 20547 40003 20553
rect 17957 20451 18015 20457
rect 15611 20420 15700 20448
rect 15764 20420 16252 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 13078 20340 13084 20392
rect 13136 20380 13142 20392
rect 13136 20352 14412 20380
rect 13136 20340 13142 20352
rect 14001 20315 14059 20321
rect 14001 20312 14013 20315
rect 12406 20284 14013 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 14001 20281 14013 20284
rect 14047 20281 14059 20315
rect 14384 20312 14412 20352
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 15194 20380 15200 20392
rect 14691 20352 15200 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 15194 20340 15200 20352
rect 15252 20380 15258 20392
rect 15764 20380 15792 20420
rect 15252 20352 15792 20380
rect 15252 20340 15258 20352
rect 16114 20340 16120 20392
rect 16172 20340 16178 20392
rect 16224 20389 16252 20420
rect 17957 20417 17969 20451
rect 18003 20448 18015 20451
rect 18064 20448 18092 20544
rect 20070 20516 20076 20528
rect 19812 20488 20076 20516
rect 18003 20420 18092 20448
rect 18509 20451 18567 20457
rect 18003 20417 18015 20420
rect 17957 20411 18015 20417
rect 18509 20417 18521 20451
rect 18555 20448 18567 20451
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 18555 20420 19165 20448
rect 18555 20417 18567 20420
rect 18509 20411 18567 20417
rect 19153 20417 19165 20420
rect 19199 20448 19211 20451
rect 19610 20448 19616 20460
rect 19199 20420 19616 20448
rect 19199 20417 19211 20420
rect 19153 20411 19211 20417
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19812 20457 19840 20488
rect 20070 20476 20076 20488
rect 20128 20516 20134 20528
rect 20128 20488 23428 20516
rect 20128 20476 20134 20488
rect 19797 20451 19855 20457
rect 19797 20417 19809 20451
rect 19843 20417 19855 20451
rect 19797 20411 19855 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 21315 20420 22661 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23400 20457 23428 20488
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20417 23443 20451
rect 23385 20411 23443 20417
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24228 20448 24256 20544
rect 38764 20516 38792 20544
rect 31588 20488 32536 20516
rect 24167 20420 24256 20448
rect 31205 20451 31263 20457
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 31205 20417 31217 20451
rect 31251 20448 31263 20451
rect 31294 20448 31300 20460
rect 31251 20420 31300 20448
rect 31251 20417 31263 20420
rect 31205 20411 31263 20417
rect 31294 20408 31300 20420
rect 31352 20408 31358 20460
rect 31386 20408 31392 20460
rect 31444 20408 31450 20460
rect 31588 20457 31616 20488
rect 32508 20460 32536 20488
rect 37936 20488 38792 20516
rect 38856 20516 38884 20544
rect 38856 20488 38962 20516
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 31938 20448 31944 20460
rect 31803 20420 31944 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 31938 20408 31944 20420
rect 31996 20408 32002 20460
rect 32125 20451 32183 20457
rect 32125 20417 32137 20451
rect 32171 20448 32183 20451
rect 32214 20448 32220 20460
rect 32171 20420 32220 20448
rect 32171 20417 32183 20420
rect 32125 20411 32183 20417
rect 32214 20408 32220 20420
rect 32272 20408 32278 20460
rect 32398 20408 32404 20460
rect 32456 20408 32462 20460
rect 32490 20408 32496 20460
rect 32548 20408 32554 20460
rect 35802 20408 35808 20460
rect 35860 20448 35866 20460
rect 35989 20451 36047 20457
rect 35989 20448 36001 20451
rect 35860 20420 36001 20448
rect 35860 20408 35866 20420
rect 35989 20417 36001 20420
rect 36035 20417 36047 20451
rect 35989 20411 36047 20417
rect 36173 20451 36231 20457
rect 36173 20417 36185 20451
rect 36219 20448 36231 20451
rect 36446 20448 36452 20460
rect 36219 20420 36452 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 37936 20457 37964 20488
rect 37921 20451 37979 20457
rect 37921 20417 37933 20451
rect 37967 20417 37979 20451
rect 37921 20411 37979 20417
rect 38194 20408 38200 20460
rect 38252 20408 38258 20460
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20349 16267 20383
rect 16209 20343 16267 20349
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18414 20380 18420 20392
rect 17920 20352 18420 20380
rect 17920 20340 17926 20352
rect 18414 20340 18420 20352
rect 18472 20380 18478 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18472 20352 18613 20380
rect 18472 20340 18478 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 18601 20343 18659 20349
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 20036 20352 21465 20380
rect 20036 20340 20042 20352
rect 21453 20349 21465 20352
rect 21499 20380 21511 20383
rect 21726 20380 21732 20392
rect 21499 20352 21732 20380
rect 21499 20349 21511 20352
rect 21453 20343 21511 20349
rect 21726 20340 21732 20352
rect 21784 20380 21790 20392
rect 22281 20383 22339 20389
rect 21784 20352 22094 20380
rect 21784 20340 21790 20352
rect 17954 20312 17960 20324
rect 14384 20284 17960 20312
rect 14001 20275 14059 20281
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 18049 20315 18107 20321
rect 18049 20281 18061 20315
rect 18095 20312 18107 20315
rect 18322 20312 18328 20324
rect 18095 20284 18328 20312
rect 18095 20281 18107 20284
rect 18049 20275 18107 20281
rect 18322 20272 18328 20284
rect 18380 20272 18386 20324
rect 22066 20312 22094 20352
rect 22281 20349 22293 20383
rect 22327 20380 22339 20383
rect 22370 20380 22376 20392
rect 22327 20352 22376 20380
rect 22327 20349 22339 20352
rect 22281 20343 22339 20349
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 31481 20383 31539 20389
rect 31481 20349 31493 20383
rect 31527 20380 31539 20383
rect 31527 20352 31754 20380
rect 31527 20349 31539 20352
rect 31481 20343 31539 20349
rect 22480 20312 22508 20340
rect 22066 20284 22508 20312
rect 31726 20324 31754 20352
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 32585 20383 32643 20389
rect 32585 20349 32597 20383
rect 32631 20380 32643 20383
rect 32766 20380 32772 20392
rect 32631 20352 32772 20380
rect 32631 20349 32643 20352
rect 32585 20343 32643 20349
rect 31726 20284 31760 20324
rect 31754 20272 31760 20284
rect 31812 20312 31818 20324
rect 32600 20312 32628 20343
rect 32766 20340 32772 20352
rect 32824 20340 32830 20392
rect 38473 20383 38531 20389
rect 38473 20380 38485 20383
rect 38120 20352 38485 20380
rect 38120 20321 38148 20352
rect 38473 20349 38485 20352
rect 38519 20349 38531 20383
rect 38473 20343 38531 20349
rect 31812 20284 32628 20312
rect 38105 20315 38163 20321
rect 31812 20272 31818 20284
rect 38105 20281 38117 20315
rect 38151 20281 38163 20315
rect 38105 20275 38163 20281
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13596 20216 13645 20244
rect 13596 20204 13602 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 13633 20207 13691 20213
rect 15378 20204 15384 20256
rect 15436 20204 15442 20256
rect 31205 20247 31263 20253
rect 31205 20213 31217 20247
rect 31251 20244 31263 20247
rect 32582 20244 32588 20256
rect 31251 20216 32588 20244
rect 31251 20213 31263 20216
rect 31205 20207 31263 20213
rect 32582 20204 32588 20216
rect 32640 20204 32646 20256
rect 35989 20247 36047 20253
rect 35989 20213 36001 20247
rect 36035 20244 36047 20247
rect 36814 20244 36820 20256
rect 36035 20216 36820 20244
rect 36035 20213 36047 20216
rect 35989 20207 36047 20213
rect 36814 20204 36820 20216
rect 36872 20204 36878 20256
rect 1104 20154 45172 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 45172 20154
rect 1104 20080 45172 20102
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 13446 20040 13452 20052
rect 12124 20012 13452 20040
rect 12124 20000 12130 20012
rect 13446 20000 13452 20012
rect 13504 20040 13510 20052
rect 19426 20040 19432 20052
rect 13504 20012 19432 20040
rect 13504 20000 13510 20012
rect 19426 20000 19432 20012
rect 19484 20040 19490 20052
rect 28813 20043 28871 20049
rect 28813 20040 28825 20043
rect 19484 20012 22508 20040
rect 19484 20000 19490 20012
rect 13541 19975 13599 19981
rect 13541 19941 13553 19975
rect 13587 19972 13599 19975
rect 14090 19972 14096 19984
rect 13587 19944 14096 19972
rect 13587 19941 13599 19944
rect 13541 19935 13599 19941
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 15102 19932 15108 19984
rect 15160 19932 15166 19984
rect 19245 19975 19303 19981
rect 19245 19972 19257 19975
rect 18892 19944 19257 19972
rect 15197 19907 15255 19913
rect 15197 19873 15209 19907
rect 15243 19904 15255 19907
rect 15470 19904 15476 19916
rect 15243 19876 15476 19904
rect 15243 19873 15255 19876
rect 15197 19867 15255 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15930 19864 15936 19916
rect 15988 19904 15994 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 15988 19876 16957 19904
rect 15988 19864 15994 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 11974 19836 11980 19848
rect 10183 19808 11980 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 11072 19780 11100 19808
rect 11974 19796 11980 19808
rect 12032 19836 12038 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 12032 19808 12173 19836
rect 12032 19796 12038 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 16758 19796 16764 19848
rect 16816 19836 16822 19848
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 16816 19808 17141 19836
rect 16816 19796 16822 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 17678 19796 17684 19848
rect 17736 19796 17742 19848
rect 18892 19845 18920 19944
rect 19245 19941 19257 19944
rect 19291 19941 19303 19975
rect 19245 19935 19303 19941
rect 19610 19932 19616 19984
rect 19668 19932 19674 19984
rect 19628 19845 19656 19932
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 19978 19904 19984 19916
rect 19935 19876 19984 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 21266 19864 21272 19916
rect 21324 19904 21330 19916
rect 22002 19904 22008 19916
rect 21324 19876 22008 19904
rect 21324 19864 21330 19876
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 21910 19796 21916 19848
rect 21968 19836 21974 19848
rect 22480 19845 22508 20012
rect 25516 20012 28825 20040
rect 25516 19916 25544 20012
rect 28813 20009 28825 20012
rect 28859 20040 28871 20043
rect 29178 20040 29184 20052
rect 28859 20012 29184 20040
rect 28859 20009 28871 20012
rect 28813 20003 28871 20009
rect 29178 20000 29184 20012
rect 29236 20000 29242 20052
rect 29273 20043 29331 20049
rect 29273 20009 29285 20043
rect 29319 20040 29331 20043
rect 29454 20040 29460 20052
rect 29319 20012 29460 20040
rect 29319 20009 29331 20012
rect 29273 20003 29331 20009
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 31938 20040 31944 20052
rect 31220 20012 31944 20040
rect 25498 19864 25504 19916
rect 25556 19864 25562 19916
rect 28994 19864 29000 19916
rect 29052 19864 29058 19916
rect 29638 19864 29644 19916
rect 29696 19864 29702 19916
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21968 19808 22109 19836
rect 21968 19796 21974 19808
rect 22097 19805 22109 19808
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 26786 19836 26792 19848
rect 26467 19808 26792 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26786 19796 26792 19808
rect 26844 19796 26850 19848
rect 28718 19796 28724 19848
rect 28776 19836 28782 19848
rect 29089 19839 29147 19845
rect 29089 19836 29101 19839
rect 28776 19808 29101 19836
rect 28776 19796 28782 19808
rect 29089 19805 29101 19808
rect 29135 19836 29147 19839
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29135 19808 29745 19836
rect 29135 19805 29147 19808
rect 29089 19799 29147 19805
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 31018 19796 31024 19848
rect 31076 19796 31082 19848
rect 31220 19845 31248 20012
rect 31938 20000 31944 20012
rect 31996 20000 32002 20052
rect 32214 20000 32220 20052
rect 32272 20000 32278 20052
rect 32398 20000 32404 20052
rect 32456 20040 32462 20052
rect 32677 20043 32735 20049
rect 32677 20040 32689 20043
rect 32456 20012 32689 20040
rect 32456 20000 32462 20012
rect 32677 20009 32689 20012
rect 32723 20009 32735 20043
rect 32677 20003 32735 20009
rect 34701 20043 34759 20049
rect 34701 20009 34713 20043
rect 34747 20009 34759 20043
rect 34701 20003 34759 20009
rect 31386 19932 31392 19984
rect 31444 19972 31450 19984
rect 31444 19944 31800 19972
rect 31444 19932 31450 19944
rect 31662 19864 31668 19916
rect 31720 19864 31726 19916
rect 31772 19913 31800 19944
rect 32490 19932 32496 19984
rect 32548 19972 32554 19984
rect 34716 19972 34744 20003
rect 35618 20000 35624 20052
rect 35676 20040 35682 20052
rect 35897 20043 35955 20049
rect 35897 20040 35909 20043
rect 35676 20012 35909 20040
rect 35676 20000 35682 20012
rect 35897 20009 35909 20012
rect 35943 20009 35955 20043
rect 35897 20003 35955 20009
rect 38841 20043 38899 20049
rect 38841 20009 38853 20043
rect 38887 20040 38899 20043
rect 38930 20040 38936 20052
rect 38887 20012 38936 20040
rect 38887 20009 38899 20012
rect 38841 20003 38899 20009
rect 38930 20000 38936 20012
rect 38988 20000 38994 20052
rect 32548 19944 34744 19972
rect 35253 19975 35311 19981
rect 32548 19932 32554 19944
rect 35253 19941 35265 19975
rect 35299 19972 35311 19975
rect 35802 19972 35808 19984
rect 35299 19944 35808 19972
rect 35299 19941 35311 19944
rect 35253 19935 35311 19941
rect 35802 19932 35808 19944
rect 35860 19932 35866 19984
rect 31757 19907 31815 19913
rect 31757 19873 31769 19907
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 34698 19864 34704 19916
rect 34756 19904 34762 19916
rect 35069 19907 35127 19913
rect 35069 19904 35081 19907
rect 34756 19876 35081 19904
rect 34756 19864 34762 19876
rect 35069 19873 35081 19876
rect 35115 19873 35127 19907
rect 35069 19867 35127 19873
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19904 35219 19907
rect 35621 19907 35679 19913
rect 35621 19904 35633 19907
rect 35207 19876 35633 19904
rect 35207 19873 35219 19876
rect 35161 19867 35219 19873
rect 35621 19873 35633 19876
rect 35667 19873 35679 19907
rect 35621 19867 35679 19873
rect 35894 19864 35900 19916
rect 35952 19904 35958 19916
rect 37185 19907 37243 19913
rect 37185 19904 37197 19907
rect 35952 19876 37197 19904
rect 35952 19864 35958 19876
rect 37185 19873 37197 19876
rect 37231 19873 37243 19907
rect 37185 19867 37243 19873
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19805 31263 19839
rect 31205 19799 31263 19805
rect 31386 19796 31392 19848
rect 31444 19796 31450 19848
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19805 31539 19839
rect 31481 19799 31539 19805
rect 31849 19839 31907 19845
rect 31849 19805 31861 19839
rect 31895 19805 31907 19839
rect 31849 19799 31907 19805
rect 10404 19771 10462 19777
rect 10404 19737 10416 19771
rect 10450 19768 10462 19771
rect 10686 19768 10692 19780
rect 10450 19740 10692 19768
rect 10450 19737 10462 19740
rect 10404 19731 10462 19737
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 11054 19728 11060 19780
rect 11112 19728 11118 19780
rect 12434 19777 12440 19780
rect 12406 19771 12440 19777
rect 12406 19737 12418 19771
rect 12406 19731 12440 19737
rect 12434 19728 12440 19731
rect 12492 19728 12498 19780
rect 15378 19728 15384 19780
rect 15436 19768 15442 19780
rect 15473 19771 15531 19777
rect 15473 19768 15485 19771
rect 15436 19740 15485 19768
rect 15436 19728 15442 19740
rect 15473 19737 15485 19740
rect 15519 19737 15531 19771
rect 15473 19731 15531 19737
rect 16022 19728 16028 19780
rect 16080 19728 16086 19780
rect 16868 19740 22094 19768
rect 11514 19660 11520 19712
rect 11572 19660 11578 19712
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 16868 19700 16896 19740
rect 12124 19672 16896 19700
rect 12124 19660 12130 19672
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19978 19700 19984 19712
rect 19751 19672 19984 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 21542 19660 21548 19712
rect 21600 19660 21606 19712
rect 22066 19700 22094 19740
rect 23934 19728 23940 19780
rect 23992 19768 23998 19780
rect 24029 19771 24087 19777
rect 24029 19768 24041 19771
rect 23992 19740 24041 19768
rect 23992 19728 23998 19740
rect 24029 19737 24041 19740
rect 24075 19768 24087 19771
rect 24394 19768 24400 19780
rect 24075 19740 24400 19768
rect 24075 19737 24087 19740
rect 24029 19731 24087 19737
rect 24394 19728 24400 19740
rect 24452 19768 24458 19780
rect 26970 19768 26976 19780
rect 24452 19740 26976 19768
rect 24452 19728 24458 19740
rect 26970 19728 26976 19740
rect 27028 19728 27034 19780
rect 28813 19771 28871 19777
rect 28813 19737 28825 19771
rect 28859 19768 28871 19771
rect 28902 19768 28908 19780
rect 28859 19740 28908 19768
rect 28859 19737 28871 19740
rect 28813 19731 28871 19737
rect 28902 19728 28908 19740
rect 28960 19728 28966 19780
rect 31294 19768 31300 19780
rect 30116 19740 31300 19768
rect 22462 19700 22468 19712
rect 22066 19672 22468 19700
rect 22462 19660 22468 19672
rect 22520 19660 22526 19712
rect 26605 19703 26663 19709
rect 26605 19669 26617 19703
rect 26651 19700 26663 19703
rect 27154 19700 27160 19712
rect 26651 19672 27160 19700
rect 26651 19669 26663 19672
rect 26605 19663 26663 19669
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 28994 19660 29000 19712
rect 29052 19700 29058 19712
rect 29730 19700 29736 19712
rect 29052 19672 29736 19700
rect 29052 19660 29058 19672
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30116 19709 30144 19740
rect 31294 19728 31300 19740
rect 31352 19768 31358 19780
rect 31496 19768 31524 19799
rect 31864 19768 31892 19799
rect 31938 19796 31944 19848
rect 31996 19836 32002 19848
rect 32033 19839 32091 19845
rect 32033 19836 32045 19839
rect 31996 19808 32045 19836
rect 31996 19796 32002 19808
rect 32033 19805 32045 19808
rect 32079 19805 32091 19839
rect 32033 19799 32091 19805
rect 32306 19796 32312 19848
rect 32364 19796 32370 19848
rect 32493 19839 32551 19845
rect 32493 19805 32505 19839
rect 32539 19836 32551 19839
rect 32582 19836 32588 19848
rect 32539 19808 32588 19836
rect 32539 19805 32551 19808
rect 32493 19799 32551 19805
rect 32582 19796 32588 19808
rect 32640 19796 32646 19848
rect 33689 19839 33747 19845
rect 33689 19836 33701 19839
rect 33060 19808 33701 19836
rect 31352 19740 31892 19768
rect 31352 19728 31358 19740
rect 33060 19712 33088 19808
rect 33689 19805 33701 19808
rect 33735 19805 33747 19839
rect 33689 19799 33747 19805
rect 33965 19839 34023 19845
rect 33965 19805 33977 19839
rect 34011 19805 34023 19839
rect 33965 19799 34023 19805
rect 34149 19839 34207 19845
rect 34149 19805 34161 19839
rect 34195 19836 34207 19839
rect 34977 19839 35035 19845
rect 34977 19836 34989 19839
rect 34195 19808 34989 19836
rect 34195 19805 34207 19808
rect 34149 19799 34207 19805
rect 34977 19805 34989 19808
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 33980 19768 34008 19799
rect 35434 19796 35440 19848
rect 35492 19796 35498 19848
rect 35526 19796 35532 19848
rect 35584 19796 35590 19848
rect 35713 19839 35771 19845
rect 35713 19805 35725 19839
rect 35759 19805 35771 19839
rect 35713 19799 35771 19805
rect 35989 19839 36047 19845
rect 35989 19805 36001 19839
rect 36035 19805 36047 19839
rect 35989 19799 36047 19805
rect 34882 19768 34888 19780
rect 33980 19740 34888 19768
rect 34882 19728 34888 19740
rect 34940 19728 34946 19780
rect 35728 19712 35756 19799
rect 36004 19768 36032 19799
rect 36170 19796 36176 19848
rect 36228 19796 36234 19848
rect 37274 19796 37280 19848
rect 37332 19796 37338 19848
rect 39025 19839 39083 19845
rect 39025 19805 39037 19839
rect 39071 19836 39083 19839
rect 39482 19836 39488 19848
rect 39071 19808 39488 19836
rect 39071 19805 39083 19808
rect 39025 19799 39083 19805
rect 39482 19796 39488 19808
rect 39540 19796 39546 19848
rect 37292 19768 37320 19796
rect 36004 19740 37320 19768
rect 39209 19771 39267 19777
rect 39209 19737 39221 19771
rect 39255 19768 39267 19771
rect 39298 19768 39304 19780
rect 39255 19740 39304 19768
rect 39255 19737 39267 19740
rect 39209 19731 39267 19737
rect 39298 19728 39304 19740
rect 39356 19728 39362 19780
rect 30101 19703 30159 19709
rect 30101 19669 30113 19703
rect 30147 19669 30159 19703
rect 30101 19663 30159 19669
rect 31205 19703 31263 19709
rect 31205 19669 31217 19703
rect 31251 19700 31263 19703
rect 31754 19700 31760 19712
rect 31251 19672 31760 19700
rect 31251 19669 31263 19672
rect 31205 19663 31263 19669
rect 31754 19660 31760 19672
rect 31812 19660 31818 19712
rect 33042 19660 33048 19712
rect 33100 19660 33106 19712
rect 33781 19703 33839 19709
rect 33781 19669 33793 19703
rect 33827 19700 33839 19703
rect 34422 19700 34428 19712
rect 33827 19672 34428 19700
rect 33827 19669 33839 19672
rect 33781 19663 33839 19669
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 35710 19660 35716 19712
rect 35768 19660 35774 19712
rect 35802 19660 35808 19712
rect 35860 19700 35866 19712
rect 36630 19700 36636 19712
rect 35860 19672 36636 19700
rect 35860 19660 35866 19672
rect 36630 19660 36636 19672
rect 36688 19660 36694 19712
rect 36722 19660 36728 19712
rect 36780 19700 36786 19712
rect 36817 19703 36875 19709
rect 36817 19700 36829 19703
rect 36780 19672 36829 19700
rect 36780 19660 36786 19672
rect 36817 19669 36829 19672
rect 36863 19669 36875 19703
rect 36817 19663 36875 19669
rect 36906 19660 36912 19712
rect 36964 19660 36970 19712
rect 1104 19610 45172 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 45172 19610
rect 1104 19536 45172 19558
rect 10686 19456 10692 19508
rect 10744 19456 10750 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 11532 19360 11560 19459
rect 11882 19456 11888 19508
rect 11940 19456 11946 19508
rect 12345 19499 12403 19505
rect 12345 19465 12357 19499
rect 12391 19496 12403 19499
rect 12434 19496 12440 19508
rect 12391 19468 12440 19496
rect 12391 19465 12403 19468
rect 12345 19459 12403 19465
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 12621 19499 12679 19505
rect 12621 19465 12633 19499
rect 12667 19465 12679 19499
rect 12621 19459 12679 19465
rect 12989 19499 13047 19505
rect 12989 19465 13001 19499
rect 13035 19496 13047 19499
rect 14458 19496 14464 19508
rect 13035 19468 14464 19496
rect 13035 19465 13047 19468
rect 12989 19459 13047 19465
rect 10919 19332 11560 19360
rect 11900 19360 11928 19456
rect 12434 19360 12440 19372
rect 11900 19332 12440 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12636 19360 12664 19459
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 14829 19499 14887 19505
rect 14829 19496 14841 19499
rect 14608 19468 14841 19496
rect 14608 19456 14614 19468
rect 14829 19465 14841 19468
rect 14875 19465 14887 19499
rect 14829 19459 14887 19465
rect 14921 19499 14979 19505
rect 14921 19465 14933 19499
rect 14967 19496 14979 19499
rect 15194 19496 15200 19508
rect 14967 19468 15200 19496
rect 14967 19465 14979 19468
rect 14921 19459 14979 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19496 15439 19499
rect 16022 19496 16028 19508
rect 15427 19468 16028 19496
rect 15427 19465 15439 19468
rect 15381 19459 15439 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 16114 19456 16120 19508
rect 16172 19496 16178 19508
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 16172 19468 17049 19496
rect 16172 19456 16178 19468
rect 17037 19465 17049 19468
rect 17083 19465 17095 19499
rect 17037 19459 17095 19465
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17678 19496 17684 19508
rect 17451 19468 17684 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 13078 19388 13084 19440
rect 13136 19388 13142 19440
rect 13538 19428 13544 19440
rect 13464 19400 13544 19428
rect 13464 19369 13492 19400
rect 13538 19388 13544 19400
rect 13596 19428 13602 19440
rect 15470 19428 15476 19440
rect 13596 19400 15476 19428
rect 13596 19388 13602 19400
rect 15470 19388 15476 19400
rect 15528 19388 15534 19440
rect 16758 19428 16764 19440
rect 16316 19400 16764 19428
rect 12575 19332 12664 19360
rect 13449 19363 13507 19369
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 13449 19329 13461 19363
rect 13495 19329 13507 19363
rect 13449 19323 13507 19329
rect 13716 19363 13774 19369
rect 13716 19329 13728 19363
rect 13762 19360 13774 19363
rect 14090 19360 14096 19372
rect 13762 19332 14096 19360
rect 13762 19329 13774 19332
rect 13716 19323 13774 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 16316 19369 16344 19400
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 15160 19332 15301 19360
rect 15160 19320 15166 19332
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19329 17003 19363
rect 17052 19360 17080 19459
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 18690 19456 18696 19508
rect 18748 19456 18754 19508
rect 19705 19499 19763 19505
rect 19705 19465 19717 19499
rect 19751 19496 19763 19499
rect 20070 19496 20076 19508
rect 19751 19468 20076 19496
rect 19751 19465 19763 19468
rect 19705 19459 19763 19465
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20947 19468 22094 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 18592 19431 18650 19437
rect 18592 19397 18604 19431
rect 18638 19428 18650 19431
rect 18708 19428 18736 19456
rect 21174 19428 21180 19440
rect 18638 19400 18736 19428
rect 20640 19400 21180 19428
rect 18638 19397 18650 19400
rect 18592 19391 18650 19397
rect 17497 19363 17555 19369
rect 17497 19360 17509 19363
rect 17052 19332 17509 19360
rect 16945 19323 17003 19329
rect 17497 19329 17509 19332
rect 17543 19329 17555 19363
rect 20640 19360 20668 19400
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 22066 19437 22094 19468
rect 23934 19456 23940 19508
rect 23992 19456 23998 19508
rect 28718 19496 28724 19508
rect 26804 19468 28724 19496
rect 21637 19431 21695 19437
rect 21637 19397 21649 19431
rect 21683 19428 21695 19431
rect 22066 19431 22124 19437
rect 21683 19400 21956 19428
rect 21683 19397 21695 19400
rect 21637 19391 21695 19397
rect 17497 19323 17555 19329
rect 17604 19332 20668 19360
rect 20717 19363 20775 19369
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 12066 19292 12072 19304
rect 12023 19264 12072 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12207 19264 13185 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 13173 19255 13231 19261
rect 15396 19264 15485 19292
rect 13188 19156 13216 19255
rect 15396 19156 15424 19264
rect 15473 19261 15485 19264
rect 15519 19292 15531 19295
rect 16758 19292 16764 19304
rect 15519 19264 16764 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 16960 19292 16988 19323
rect 17604 19292 17632 19332
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 21818 19360 21824 19372
rect 20717 19323 20775 19329
rect 20824 19332 21824 19360
rect 16960 19264 17632 19292
rect 18046 19252 18052 19304
rect 18104 19252 18110 19304
rect 18322 19252 18328 19304
rect 18380 19252 18386 19304
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 20732 19224 20760 19323
rect 20824 19304 20852 19332
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 21928 19360 21956 19400
rect 22066 19397 22078 19431
rect 22112 19397 22124 19431
rect 22066 19391 22124 19397
rect 22370 19388 22376 19440
rect 22428 19428 22434 19440
rect 23198 19428 23204 19440
rect 22428 19400 23204 19428
rect 22428 19388 22434 19400
rect 23198 19388 23204 19400
rect 23256 19388 23262 19440
rect 23952 19428 23980 19456
rect 25958 19428 25964 19440
rect 23860 19400 23980 19428
rect 25346 19400 25964 19428
rect 23382 19360 23388 19372
rect 21928 19332 23388 19360
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 23860 19369 23888 19400
rect 25958 19388 25964 19400
rect 26016 19388 26022 19440
rect 26421 19431 26479 19437
rect 26421 19397 26433 19431
rect 26467 19428 26479 19431
rect 26804 19428 26832 19468
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 29365 19499 29423 19505
rect 29365 19465 29377 19499
rect 29411 19496 29423 19499
rect 29638 19496 29644 19508
rect 29411 19468 29644 19496
rect 29411 19465 29423 19468
rect 29365 19459 29423 19465
rect 29638 19456 29644 19468
rect 29696 19456 29702 19508
rect 29730 19456 29736 19508
rect 29788 19496 29794 19508
rect 29788 19468 30604 19496
rect 29788 19456 29794 19468
rect 26467 19400 26832 19428
rect 26467 19397 26479 19400
rect 26421 19391 26479 19397
rect 27154 19388 27160 19440
rect 27212 19428 27218 19440
rect 27249 19431 27307 19437
rect 27249 19428 27261 19431
rect 27212 19400 27261 19428
rect 27212 19388 27218 19400
rect 27249 19397 27261 19400
rect 27295 19397 27307 19431
rect 27249 19391 27307 19397
rect 27706 19388 27712 19440
rect 27764 19388 27770 19440
rect 29270 19388 29276 19440
rect 29328 19428 29334 19440
rect 30576 19428 30604 19468
rect 31018 19456 31024 19508
rect 31076 19496 31082 19508
rect 31113 19499 31171 19505
rect 31113 19496 31125 19499
rect 31076 19468 31125 19496
rect 31076 19456 31082 19468
rect 31113 19465 31125 19468
rect 31159 19465 31171 19499
rect 31113 19459 31171 19465
rect 31386 19456 31392 19508
rect 31444 19456 31450 19508
rect 31938 19456 31944 19508
rect 31996 19456 32002 19508
rect 34698 19456 34704 19508
rect 34756 19496 34762 19508
rect 34793 19499 34851 19505
rect 34793 19496 34805 19499
rect 34756 19468 34805 19496
rect 34756 19456 34762 19468
rect 34793 19465 34805 19468
rect 34839 19465 34851 19499
rect 34793 19459 34851 19465
rect 34882 19456 34888 19508
rect 34940 19456 34946 19508
rect 35526 19456 35532 19508
rect 35584 19456 35590 19508
rect 36357 19431 36415 19437
rect 29328 19400 30328 19428
rect 29328 19388 29334 19400
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 26329 19363 26387 19369
rect 26329 19360 26341 19363
rect 23845 19323 23903 19329
rect 25332 19332 26341 19360
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 21082 19252 21088 19304
rect 21140 19252 21146 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23768 19264 24133 19292
rect 21450 19224 21456 19236
rect 16080 19196 18368 19224
rect 20732 19196 21456 19224
rect 16080 19184 16086 19196
rect 13188 19128 15424 19156
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15988 19128 16129 19156
rect 15988 19116 15994 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 18340 19156 18368 19196
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 23768 19233 23796 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 23753 19227 23811 19233
rect 23753 19193 23765 19227
rect 23799 19193 23811 19227
rect 23753 19187 23811 19193
rect 21634 19156 21640 19168
rect 18340 19128 21640 19156
rect 16117 19119 16175 19125
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 22520 19128 23213 19156
rect 22520 19116 22526 19128
rect 23201 19125 23213 19128
rect 23247 19156 23259 19159
rect 25332 19156 25360 19332
rect 26329 19329 26341 19332
rect 26375 19329 26387 19363
rect 26329 19323 26387 19329
rect 26786 19320 26792 19372
rect 26844 19320 26850 19372
rect 26970 19320 26976 19372
rect 27028 19320 27034 19372
rect 28905 19363 28963 19369
rect 28905 19329 28917 19363
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 26234 19252 26240 19304
rect 26292 19252 26298 19304
rect 26804 19233 26832 19320
rect 28718 19252 28724 19304
rect 28776 19292 28782 19304
rect 28920 19292 28948 19323
rect 28994 19320 29000 19372
rect 29052 19360 29058 19372
rect 29089 19363 29147 19369
rect 29089 19360 29101 19363
rect 29052 19332 29101 19360
rect 29052 19320 29058 19332
rect 29089 19329 29101 19332
rect 29135 19329 29147 19363
rect 29089 19323 29147 19329
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 30300 19369 30328 19400
rect 30576 19400 30880 19428
rect 30576 19369 30604 19400
rect 30852 19369 30880 19400
rect 31220 19400 31800 19428
rect 31220 19369 31248 19400
rect 29641 19366 29699 19369
rect 29472 19363 29699 19366
rect 29472 19360 29653 19363
rect 29236 19338 29653 19360
rect 29236 19332 29500 19338
rect 29629 19332 29653 19338
rect 29236 19320 29242 19332
rect 29641 19329 29653 19332
rect 29687 19329 29699 19363
rect 29641 19323 29699 19329
rect 30285 19363 30343 19369
rect 30285 19329 30297 19363
rect 30331 19329 30343 19363
rect 30285 19323 30343 19329
rect 30561 19363 30619 19369
rect 30561 19329 30573 19363
rect 30607 19329 30619 19363
rect 30561 19323 30619 19329
rect 30653 19363 30711 19369
rect 30653 19329 30665 19363
rect 30699 19329 30711 19363
rect 30653 19323 30711 19329
rect 30837 19363 30895 19369
rect 30837 19329 30849 19363
rect 30883 19329 30895 19363
rect 30837 19323 30895 19329
rect 31021 19363 31079 19369
rect 31021 19329 31033 19363
rect 31067 19329 31079 19363
rect 31021 19323 31079 19329
rect 31205 19363 31263 19369
rect 31205 19329 31217 19363
rect 31251 19329 31263 19363
rect 31205 19323 31263 19329
rect 29270 19292 29276 19304
rect 28776 19264 29276 19292
rect 28776 19252 28782 19264
rect 29270 19252 29276 19264
rect 29328 19252 29334 19304
rect 29733 19295 29791 19301
rect 29733 19261 29745 19295
rect 29779 19292 29791 19295
rect 30101 19295 30159 19301
rect 30101 19292 30113 19295
rect 29779 19264 30113 19292
rect 29779 19261 29791 19264
rect 29733 19255 29791 19261
rect 30101 19261 30113 19264
rect 30147 19261 30159 19295
rect 30300 19292 30328 19323
rect 30668 19292 30696 19323
rect 30300 19264 30696 19292
rect 31036 19292 31064 19323
rect 31478 19320 31484 19372
rect 31536 19320 31542 19372
rect 31772 19369 31800 19400
rect 34348 19400 35112 19428
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19329 31631 19363
rect 31573 19323 31631 19329
rect 31757 19363 31815 19369
rect 31757 19329 31769 19363
rect 31803 19360 31815 19363
rect 33410 19360 33416 19372
rect 31803 19332 33416 19360
rect 31803 19329 31815 19332
rect 31757 19323 31815 19329
rect 31588 19292 31616 19323
rect 33410 19320 33416 19332
rect 33468 19320 33474 19372
rect 33870 19320 33876 19372
rect 33928 19320 33934 19372
rect 31036 19264 31616 19292
rect 30101 19255 30159 19261
rect 26789 19227 26847 19233
rect 26789 19193 26801 19227
rect 26835 19193 26847 19227
rect 26789 19187 26847 19193
rect 28902 19184 28908 19236
rect 28960 19224 28966 19236
rect 28997 19227 29055 19233
rect 28997 19224 29009 19227
rect 28960 19196 29009 19224
rect 28960 19184 28966 19196
rect 28997 19193 29009 19196
rect 29043 19193 29055 19227
rect 28997 19187 29055 19193
rect 30009 19227 30067 19233
rect 30009 19193 30021 19227
rect 30055 19224 30067 19227
rect 31036 19224 31064 19264
rect 32122 19252 32128 19304
rect 32180 19252 32186 19304
rect 33042 19252 33048 19304
rect 33100 19292 33106 19304
rect 34348 19301 34376 19400
rect 34422 19320 34428 19372
rect 34480 19320 34486 19372
rect 35084 19369 35112 19400
rect 36357 19397 36369 19431
rect 36403 19428 36415 19431
rect 37645 19431 37703 19437
rect 37645 19428 37657 19431
rect 36403 19400 37657 19428
rect 36403 19397 36415 19400
rect 36357 19391 36415 19397
rect 37645 19397 37657 19400
rect 37691 19397 37703 19431
rect 37645 19391 37703 19397
rect 35069 19363 35127 19369
rect 35069 19329 35081 19363
rect 35115 19329 35127 19363
rect 35069 19323 35127 19329
rect 35161 19363 35219 19369
rect 35161 19329 35173 19363
rect 35207 19360 35219 19363
rect 35342 19360 35348 19372
rect 35207 19332 35348 19360
rect 35207 19329 35219 19332
rect 35161 19323 35219 19329
rect 34333 19295 34391 19301
rect 34333 19292 34345 19295
rect 33100 19264 34345 19292
rect 33100 19252 33106 19264
rect 34333 19261 34345 19264
rect 34379 19261 34391 19295
rect 34440 19292 34468 19320
rect 35176 19292 35204 19323
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 35437 19363 35495 19369
rect 35437 19329 35449 19363
rect 35483 19360 35495 19363
rect 35618 19360 35624 19372
rect 35483 19332 35624 19360
rect 35483 19329 35495 19332
rect 35437 19323 35495 19329
rect 35618 19320 35624 19332
rect 35676 19360 35682 19372
rect 35713 19363 35771 19369
rect 35713 19360 35725 19363
rect 35676 19332 35725 19360
rect 35676 19320 35682 19332
rect 35713 19329 35725 19332
rect 35759 19329 35771 19363
rect 35713 19323 35771 19329
rect 35894 19320 35900 19372
rect 35952 19320 35958 19372
rect 36265 19363 36323 19369
rect 36265 19329 36277 19363
rect 36311 19329 36323 19363
rect 36265 19323 36323 19329
rect 34440 19264 35204 19292
rect 34333 19255 34391 19261
rect 36280 19236 36308 19323
rect 36446 19320 36452 19372
rect 36504 19320 36510 19372
rect 36538 19320 36544 19372
rect 36596 19369 36602 19372
rect 36596 19363 36625 19369
rect 36613 19329 36625 19363
rect 36596 19323 36625 19329
rect 36596 19320 36602 19323
rect 36722 19320 36728 19372
rect 36780 19320 36786 19372
rect 36814 19320 36820 19372
rect 36872 19320 36878 19372
rect 36906 19320 36912 19372
rect 36964 19360 36970 19372
rect 37001 19363 37059 19369
rect 37001 19360 37013 19363
rect 36964 19332 37013 19360
rect 36964 19320 36970 19332
rect 37001 19329 37013 19332
rect 37047 19360 37059 19363
rect 37277 19363 37335 19369
rect 37277 19360 37289 19363
rect 37047 19332 37289 19360
rect 37047 19329 37059 19332
rect 37001 19323 37059 19329
rect 37277 19329 37289 19332
rect 37323 19329 37335 19363
rect 37277 19323 37335 19329
rect 37366 19320 37372 19372
rect 37424 19360 37430 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37424 19332 37473 19360
rect 37424 19320 37430 19332
rect 37461 19329 37473 19332
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 30055 19196 31064 19224
rect 30055 19193 30067 19196
rect 30009 19187 30067 19193
rect 23247 19128 25360 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 25498 19116 25504 19168
rect 25556 19156 25562 19168
rect 25593 19159 25651 19165
rect 25593 19156 25605 19159
rect 25556 19128 25605 19156
rect 25556 19116 25562 19128
rect 25593 19125 25605 19128
rect 25639 19125 25651 19159
rect 29012 19156 29040 19187
rect 36262 19184 36268 19236
rect 36320 19224 36326 19236
rect 36909 19227 36967 19233
rect 36909 19224 36921 19227
rect 36320 19196 36921 19224
rect 36320 19184 36326 19196
rect 36909 19193 36921 19196
rect 36955 19193 36967 19227
rect 36909 19187 36967 19193
rect 30469 19159 30527 19165
rect 30469 19156 30481 19159
rect 29012 19128 30481 19156
rect 25593 19119 25651 19125
rect 30469 19125 30481 19128
rect 30515 19125 30527 19159
rect 30469 19119 30527 19125
rect 30742 19116 30748 19168
rect 30800 19116 30806 19168
rect 31754 19116 31760 19168
rect 31812 19156 31818 19168
rect 35345 19159 35403 19165
rect 35345 19156 35357 19159
rect 31812 19128 35357 19156
rect 31812 19116 31818 19128
rect 35345 19125 35357 19128
rect 35391 19156 35403 19159
rect 35894 19156 35900 19168
rect 35391 19128 35900 19156
rect 35391 19125 35403 19128
rect 35345 19119 35403 19125
rect 35894 19116 35900 19128
rect 35952 19116 35958 19168
rect 36081 19159 36139 19165
rect 36081 19125 36093 19159
rect 36127 19156 36139 19159
rect 37274 19156 37280 19168
rect 36127 19128 37280 19156
rect 36127 19125 36139 19128
rect 36081 19119 36139 19125
rect 37274 19116 37280 19128
rect 37332 19116 37338 19168
rect 1104 19066 45172 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 45172 19066
rect 1104 18992 45172 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 1728 18924 10088 18952
rect 1728 18912 1734 18924
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 10060 18893 10088 18924
rect 12434 18912 12440 18964
rect 12492 18912 12498 18964
rect 14090 18912 14096 18964
rect 14148 18912 14154 18964
rect 17037 18955 17095 18961
rect 17037 18921 17049 18955
rect 17083 18952 17095 18955
rect 18046 18952 18052 18964
rect 17083 18924 18052 18952
rect 17083 18921 17095 18924
rect 17037 18915 17095 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19150 18952 19156 18964
rect 18156 18924 19156 18952
rect 9309 18887 9367 18893
rect 9309 18884 9321 18887
rect 1820 18856 9321 18884
rect 1820 18844 1826 18856
rect 9309 18853 9321 18856
rect 9355 18853 9367 18887
rect 9309 18847 9367 18853
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18853 10103 18887
rect 10045 18847 10103 18853
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 18156 18884 18184 18924
rect 19150 18912 19156 18924
rect 19208 18952 19214 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 19208 18924 19257 18952
rect 19208 18912 19214 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 20806 18952 20812 18964
rect 19245 18915 19303 18921
rect 20548 18924 20812 18952
rect 18012 18856 18184 18884
rect 18012 18844 18018 18856
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11572 18788 11805 18816
rect 11572 18776 11578 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 15194 18776 15200 18828
rect 15252 18776 15258 18828
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 20548 18825 20576 18924
rect 20806 18912 20812 18924
rect 20864 18912 20870 18964
rect 21450 18912 21456 18964
rect 21508 18952 21514 18964
rect 22005 18955 22063 18961
rect 22005 18952 22017 18955
rect 21508 18924 22017 18952
rect 21508 18912 21514 18924
rect 22005 18921 22017 18924
rect 22051 18921 22063 18955
rect 23477 18955 23535 18961
rect 23477 18952 23489 18955
rect 22005 18915 22063 18921
rect 23216 18924 23489 18952
rect 21634 18844 21640 18896
rect 21692 18844 21698 18896
rect 21910 18844 21916 18896
rect 21968 18884 21974 18896
rect 21968 18856 23152 18884
rect 21968 18844 21974 18856
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 15528 18788 15669 18816
rect 15528 18776 15534 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 15657 18779 15715 18785
rect 19076 18788 20545 18816
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 15930 18757 15936 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14323 18720 14657 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 15924 18748 15936 18757
rect 15891 18720 15936 18748
rect 14645 18711 14703 18717
rect 15924 18711 15936 18720
rect 15930 18708 15936 18711
rect 15988 18708 15994 18760
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 19076 18757 19104 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 20533 18779 20591 18785
rect 19061 18751 19119 18757
rect 19061 18748 19073 18751
rect 18380 18720 19073 18748
rect 18380 18708 18386 18720
rect 19061 18717 19073 18720
rect 19107 18717 19119 18751
rect 19797 18751 19855 18757
rect 19797 18748 19809 18751
rect 19061 18711 19119 18717
rect 19168 18720 19809 18748
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 9769 18683 9827 18689
rect 9769 18680 9781 18683
rect 9723 18652 9781 18680
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 9769 18649 9781 18652
rect 9815 18680 9827 18683
rect 18816 18683 18874 18689
rect 9815 18652 12434 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 6914 18612 6920 18624
rect 1627 18584 6920 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 9214 18572 9220 18624
rect 9272 18572 9278 18624
rect 10226 18572 10232 18624
rect 10284 18572 10290 18624
rect 12406 18612 12434 18652
rect 18816 18649 18828 18683
rect 18862 18680 18874 18683
rect 18966 18680 18972 18692
rect 18862 18652 18972 18680
rect 18862 18649 18874 18652
rect 18816 18643 18874 18649
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 15102 18612 15108 18624
rect 12406 18584 15108 18612
rect 15102 18572 15108 18584
rect 15160 18572 15166 18624
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 19168 18612 19196 18720
rect 19797 18717 19809 18720
rect 19843 18748 19855 18751
rect 21082 18748 21088 18760
rect 19843 18720 21088 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 21082 18708 21088 18720
rect 21140 18708 21146 18760
rect 20622 18640 20628 18692
rect 20680 18680 20686 18692
rect 20778 18683 20836 18689
rect 20778 18680 20790 18683
rect 20680 18652 20790 18680
rect 20680 18640 20686 18652
rect 20778 18649 20790 18652
rect 20824 18649 20836 18683
rect 21652 18680 21680 18844
rect 22649 18819 22707 18825
rect 22649 18785 22661 18819
rect 22695 18816 22707 18819
rect 22738 18816 22744 18828
rect 22695 18788 22744 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 22554 18680 22560 18692
rect 21652 18652 22560 18680
rect 20778 18643 20836 18649
rect 22554 18640 22560 18652
rect 22612 18680 22618 18692
rect 23014 18680 23020 18692
rect 22612 18652 23020 18680
rect 22612 18640 22618 18652
rect 23014 18640 23020 18652
rect 23072 18640 23078 18692
rect 23124 18680 23152 18856
rect 23216 18757 23244 18924
rect 23477 18921 23489 18924
rect 23523 18921 23535 18955
rect 23477 18915 23535 18921
rect 23566 18912 23572 18964
rect 23624 18952 23630 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 23624 18924 24409 18952
rect 23624 18912 23630 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 25590 18912 25596 18964
rect 25648 18952 25654 18964
rect 33042 18952 33048 18964
rect 25648 18924 28120 18952
rect 25648 18912 25654 18924
rect 23400 18856 24440 18884
rect 23400 18828 23428 18856
rect 23382 18776 23388 18828
rect 23440 18776 23446 18828
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23716 18788 24041 18816
rect 23716 18776 23722 18788
rect 24029 18785 24041 18788
rect 24075 18816 24087 18819
rect 24210 18816 24216 18828
rect 24075 18788 24216 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 24210 18776 24216 18788
rect 24268 18776 24274 18828
rect 24412 18816 24440 18856
rect 24486 18844 24492 18896
rect 24544 18884 24550 18896
rect 26234 18884 26240 18896
rect 24544 18856 26240 18884
rect 24544 18844 24550 18856
rect 24964 18825 24992 18856
rect 26234 18844 26240 18856
rect 26292 18844 26298 18896
rect 24857 18819 24915 18825
rect 24857 18816 24869 18819
rect 24412 18788 24869 18816
rect 24857 18785 24869 18788
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 24949 18819 25007 18825
rect 24949 18785 24961 18819
rect 24995 18785 25007 18819
rect 26252 18816 26280 18844
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 26252 18788 26709 18816
rect 24949 18779 25007 18785
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 28092 18816 28120 18924
rect 31865 18924 33048 18952
rect 28169 18887 28227 18893
rect 28169 18853 28181 18887
rect 28215 18884 28227 18887
rect 28810 18884 28816 18896
rect 28215 18856 28816 18884
rect 28215 18853 28227 18856
rect 28169 18847 28227 18853
rect 28810 18844 28816 18856
rect 28868 18844 28874 18896
rect 31865 18884 31893 18924
rect 33042 18912 33048 18924
rect 33100 18912 33106 18964
rect 33410 18912 33416 18964
rect 33468 18912 33474 18964
rect 34992 18924 35664 18952
rect 32214 18884 32220 18896
rect 29380 18856 31893 18884
rect 31956 18856 32220 18884
rect 28092 18788 28580 18816
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 25590 18748 25596 18760
rect 23891 18720 25596 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 25590 18708 25596 18720
rect 25648 18708 25654 18760
rect 26513 18751 26571 18757
rect 26513 18717 26525 18751
rect 26559 18748 26571 18751
rect 27706 18748 27712 18760
rect 26559 18720 27712 18748
rect 26559 18717 26571 18720
rect 26513 18711 26571 18717
rect 27706 18708 27712 18720
rect 27764 18748 27770 18760
rect 27801 18751 27859 18757
rect 27801 18748 27813 18751
rect 27764 18720 27813 18748
rect 27764 18708 27770 18720
rect 27801 18717 27813 18720
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 27985 18751 28043 18757
rect 27985 18717 27997 18751
rect 28031 18748 28043 18751
rect 28092 18748 28120 18788
rect 28552 18757 28580 18788
rect 28626 18776 28632 18828
rect 28684 18776 28690 18828
rect 29380 18825 29408 18856
rect 29365 18819 29423 18825
rect 29365 18785 29377 18819
rect 29411 18785 29423 18819
rect 29365 18779 29423 18785
rect 30653 18819 30711 18825
rect 30653 18785 30665 18819
rect 30699 18816 30711 18819
rect 31754 18816 31760 18828
rect 30699 18788 31760 18816
rect 30699 18785 30711 18788
rect 30653 18779 30711 18785
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 28031 18720 28120 18748
rect 28537 18751 28595 18757
rect 28031 18717 28043 18720
rect 27985 18711 28043 18717
rect 28537 18717 28549 18751
rect 28583 18717 28595 18751
rect 29641 18751 29699 18757
rect 29641 18748 29653 18751
rect 28537 18711 28595 18717
rect 28966 18720 29653 18748
rect 26605 18683 26663 18689
rect 26605 18680 26617 18683
rect 23124 18652 26617 18680
rect 26605 18649 26617 18652
rect 26651 18649 26663 18683
rect 27816 18680 27844 18711
rect 28966 18680 28994 18720
rect 29641 18717 29653 18720
rect 29687 18717 29699 18751
rect 30742 18748 30748 18760
rect 30314 18720 30748 18748
rect 29641 18711 29699 18717
rect 30742 18708 30748 18720
rect 30800 18708 30806 18760
rect 31956 18757 31984 18856
rect 32214 18844 32220 18856
rect 32272 18844 32278 18896
rect 32398 18844 32404 18896
rect 32456 18884 32462 18896
rect 33137 18887 33195 18893
rect 33137 18884 33149 18887
rect 32456 18856 33149 18884
rect 32456 18844 32462 18856
rect 33137 18853 33149 18856
rect 33183 18853 33195 18887
rect 34992 18884 35020 18924
rect 33137 18847 33195 18853
rect 33244 18856 35020 18884
rect 33244 18816 33272 18856
rect 34701 18819 34759 18825
rect 34701 18816 34713 18819
rect 32692 18788 33272 18816
rect 33888 18788 34713 18816
rect 31941 18751 31999 18757
rect 31850 18729 31908 18735
rect 31850 18695 31862 18729
rect 31896 18695 31908 18729
rect 31941 18717 31953 18751
rect 31987 18717 31999 18751
rect 31941 18711 31999 18717
rect 32306 18708 32312 18760
rect 32364 18708 32370 18760
rect 32692 18748 32720 18788
rect 32416 18720 32720 18748
rect 31850 18692 31908 18695
rect 27816 18652 28994 18680
rect 26605 18643 26663 18649
rect 31846 18640 31852 18692
rect 31904 18640 31910 18692
rect 32030 18640 32036 18692
rect 32088 18640 32094 18692
rect 32171 18683 32229 18689
rect 32171 18649 32183 18683
rect 32217 18680 32229 18683
rect 32416 18680 32444 18720
rect 32766 18708 32772 18760
rect 32824 18748 32830 18760
rect 33888 18757 33916 18788
rect 34701 18785 34713 18788
rect 34747 18785 34759 18819
rect 34701 18779 34759 18785
rect 33045 18751 33103 18757
rect 33045 18748 33057 18751
rect 32824 18720 33057 18748
rect 32824 18708 32830 18720
rect 33045 18717 33057 18720
rect 33091 18717 33103 18751
rect 33045 18711 33103 18717
rect 33229 18751 33287 18757
rect 33229 18717 33241 18751
rect 33275 18717 33287 18751
rect 33229 18711 33287 18717
rect 33505 18751 33563 18757
rect 33505 18717 33517 18751
rect 33551 18748 33563 18751
rect 33873 18751 33931 18757
rect 33551 18720 33640 18748
rect 33551 18717 33563 18720
rect 33505 18711 33563 18717
rect 32217 18652 32444 18680
rect 32217 18649 32229 18652
rect 32171 18643 32229 18649
rect 32490 18640 32496 18692
rect 32548 18680 32554 18692
rect 32953 18683 33011 18689
rect 32953 18680 32965 18683
rect 32548 18652 32965 18680
rect 32548 18640 32554 18652
rect 32953 18649 32965 18652
rect 32999 18680 33011 18683
rect 33244 18680 33272 18711
rect 32999 18652 33272 18680
rect 32999 18649 33011 18652
rect 32953 18643 33011 18649
rect 33612 18624 33640 18720
rect 33873 18717 33885 18751
rect 33919 18717 33931 18751
rect 33873 18711 33931 18717
rect 34330 18708 34336 18760
rect 34388 18708 34394 18760
rect 34606 18708 34612 18760
rect 34664 18748 34670 18760
rect 34882 18748 34888 18760
rect 34664 18720 34888 18748
rect 34664 18708 34670 18720
rect 34882 18708 34888 18720
rect 34940 18708 34946 18760
rect 33965 18683 34023 18689
rect 33965 18649 33977 18683
rect 34011 18649 34023 18683
rect 33965 18643 34023 18649
rect 17727 18584 19196 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 22370 18572 22376 18624
rect 22428 18572 22434 18624
rect 22462 18572 22468 18624
rect 22520 18572 22526 18624
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 23750 18572 23756 18624
rect 23808 18612 23814 18624
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23808 18584 23949 18612
rect 23808 18572 23814 18584
rect 23937 18581 23949 18584
rect 23983 18581 23995 18615
rect 23937 18575 23995 18581
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 25498 18612 25504 18624
rect 24811 18584 25504 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 25498 18572 25504 18584
rect 25556 18572 25562 18624
rect 26142 18572 26148 18624
rect 26200 18572 26206 18624
rect 31665 18615 31723 18621
rect 31665 18581 31677 18615
rect 31711 18612 31723 18615
rect 32398 18612 32404 18624
rect 31711 18584 32404 18612
rect 31711 18581 31723 18584
rect 31665 18575 31723 18581
rect 32398 18572 32404 18584
rect 32456 18572 32462 18624
rect 32582 18572 32588 18624
rect 32640 18572 32646 18624
rect 33594 18572 33600 18624
rect 33652 18572 33658 18624
rect 33686 18572 33692 18624
rect 33744 18572 33750 18624
rect 33980 18612 34008 18643
rect 34054 18640 34060 18692
rect 34112 18640 34118 18692
rect 34195 18683 34253 18689
rect 34195 18649 34207 18683
rect 34241 18680 34253 18683
rect 34992 18680 35020 18856
rect 35526 18844 35532 18896
rect 35584 18844 35590 18896
rect 35636 18884 35664 18924
rect 35710 18912 35716 18964
rect 35768 18912 35774 18964
rect 36081 18955 36139 18961
rect 36081 18921 36093 18955
rect 36127 18952 36139 18955
rect 36170 18952 36176 18964
rect 36127 18924 36176 18952
rect 36127 18921 36139 18924
rect 36081 18915 36139 18921
rect 36170 18912 36176 18924
rect 36228 18912 36234 18964
rect 36538 18912 36544 18964
rect 36596 18912 36602 18964
rect 36556 18884 36584 18912
rect 35636 18856 36584 18884
rect 35544 18816 35572 18844
rect 35084 18788 35572 18816
rect 35084 18757 35112 18788
rect 35069 18751 35127 18757
rect 35069 18717 35081 18751
rect 35115 18717 35127 18751
rect 35069 18711 35127 18717
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18717 35219 18751
rect 35161 18711 35219 18717
rect 34241 18652 35020 18680
rect 35176 18680 35204 18711
rect 35250 18708 35256 18760
rect 35308 18708 35314 18760
rect 35544 18757 35572 18788
rect 37458 18776 37464 18828
rect 37516 18816 37522 18828
rect 37829 18819 37887 18825
rect 37829 18816 37841 18819
rect 37516 18788 37841 18816
rect 37516 18776 37522 18788
rect 37829 18785 37841 18788
rect 37875 18785 37887 18819
rect 37829 18779 37887 18785
rect 35529 18751 35587 18757
rect 35529 18717 35541 18751
rect 35575 18717 35587 18751
rect 35529 18711 35587 18717
rect 35618 18708 35624 18760
rect 35676 18708 35682 18760
rect 35805 18751 35863 18757
rect 35805 18717 35817 18751
rect 35851 18748 35863 18751
rect 35894 18748 35900 18760
rect 35851 18720 35900 18748
rect 35851 18717 35863 18720
rect 35805 18711 35863 18717
rect 35894 18708 35900 18720
rect 35952 18708 35958 18760
rect 36262 18708 36268 18760
rect 36320 18708 36326 18760
rect 35437 18683 35495 18689
rect 35437 18680 35449 18683
rect 35176 18652 35449 18680
rect 34241 18649 34253 18652
rect 34195 18643 34253 18649
rect 35437 18649 35449 18652
rect 35483 18680 35495 18683
rect 36280 18680 36308 18708
rect 35483 18652 36308 18680
rect 37122 18652 37228 18680
rect 35483 18649 35495 18652
rect 35437 18643 35495 18649
rect 35345 18615 35403 18621
rect 35345 18612 35357 18615
rect 33980 18584 35357 18612
rect 35345 18581 35357 18584
rect 35391 18581 35403 18615
rect 37200 18612 37228 18652
rect 37274 18640 37280 18692
rect 37332 18680 37338 18692
rect 37553 18683 37611 18689
rect 37553 18680 37565 18683
rect 37332 18652 37565 18680
rect 37332 18640 37338 18652
rect 37553 18649 37565 18652
rect 37599 18649 37611 18683
rect 37553 18643 37611 18649
rect 38289 18683 38347 18689
rect 38289 18649 38301 18683
rect 38335 18680 38347 18683
rect 38562 18680 38568 18692
rect 38335 18652 38568 18680
rect 38335 18649 38347 18652
rect 38289 18643 38347 18649
rect 38562 18640 38568 18652
rect 38620 18640 38626 18692
rect 38194 18612 38200 18624
rect 37200 18584 38200 18612
rect 35345 18575 35403 18581
rect 38194 18572 38200 18584
rect 38252 18572 38258 18624
rect 1104 18522 45172 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 45172 18522
rect 1104 18448 45172 18470
rect 9214 18368 9220 18420
rect 9272 18368 9278 18420
rect 10226 18368 10232 18420
rect 10284 18368 10290 18420
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 18322 18408 18328 18420
rect 16816 18380 18328 18408
rect 16816 18368 16822 18380
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19024 18380 19809 18408
rect 19024 18368 19030 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 20622 18368 20628 18420
rect 20680 18368 20686 18420
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 21085 18411 21143 18417
rect 21085 18377 21097 18411
rect 21131 18408 21143 18411
rect 21542 18408 21548 18420
rect 21131 18380 21548 18408
rect 21131 18377 21143 18380
rect 21085 18371 21143 18377
rect 9232 18272 9260 18368
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9232 18244 9873 18272
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 10244 18272 10272 18368
rect 15102 18300 15108 18352
rect 15160 18340 15166 18352
rect 15160 18312 19748 18340
rect 15160 18300 15166 18312
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10244 18244 10793 18272
rect 9861 18235 9919 18241
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 19208 18244 19257 18272
rect 19208 18232 19214 18244
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 11698 18164 11704 18216
rect 11756 18164 11762 18216
rect 18322 18164 18328 18216
rect 18380 18164 18386 18216
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 13998 18096 14004 18148
rect 14056 18136 14062 18148
rect 15381 18139 15439 18145
rect 15381 18136 15393 18139
rect 14056 18108 15393 18136
rect 14056 18096 14062 18108
rect 15381 18105 15393 18108
rect 15427 18105 15439 18139
rect 15381 18099 15439 18105
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11422 18068 11428 18080
rect 11011 18040 11428 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 12342 18028 12348 18080
rect 12400 18028 12406 18080
rect 15562 18028 15568 18080
rect 15620 18028 15626 18080
rect 18340 18068 18368 18164
rect 18708 18136 18736 18167
rect 18782 18164 18788 18216
rect 18840 18164 18846 18216
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19536 18204 19564 18235
rect 19015 18176 19564 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19058 18136 19064 18148
rect 18708 18108 19064 18136
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19337 18071 19395 18077
rect 19337 18068 19349 18071
rect 18340 18040 19349 18068
rect 19337 18037 19349 18040
rect 19383 18037 19395 18071
rect 19628 18068 19656 18235
rect 19720 18136 19748 18312
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 20732 18272 20760 18371
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 21726 18368 21732 18420
rect 21784 18408 21790 18420
rect 22738 18408 22744 18420
rect 21784 18380 22744 18408
rect 21784 18368 21790 18380
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23014 18368 23020 18420
rect 23072 18408 23078 18420
rect 23750 18408 23756 18420
rect 23072 18380 23756 18408
rect 23072 18368 23078 18380
rect 23750 18368 23756 18380
rect 23808 18368 23814 18420
rect 23934 18368 23940 18420
rect 23992 18368 23998 18420
rect 25590 18368 25596 18420
rect 25648 18368 25654 18420
rect 28626 18368 28632 18420
rect 28684 18368 28690 18420
rect 32306 18368 32312 18420
rect 32364 18408 32370 18420
rect 32769 18411 32827 18417
rect 32769 18408 32781 18411
rect 32364 18380 32781 18408
rect 32364 18368 32370 18380
rect 32769 18377 32781 18380
rect 32815 18377 32827 18411
rect 32769 18371 32827 18377
rect 34241 18411 34299 18417
rect 34241 18377 34253 18411
rect 34287 18408 34299 18411
rect 34330 18408 34336 18420
rect 34287 18380 34336 18408
rect 34287 18377 34299 18380
rect 34241 18371 34299 18377
rect 34330 18368 34336 18380
rect 34388 18368 34394 18420
rect 35342 18368 35348 18420
rect 35400 18408 35406 18420
rect 35989 18411 36047 18417
rect 35989 18408 36001 18411
rect 35400 18380 36001 18408
rect 35400 18368 35406 18380
rect 35989 18377 36001 18380
rect 36035 18377 36047 18411
rect 35989 18371 36047 18377
rect 36170 18368 36176 18420
rect 36228 18368 36234 18420
rect 38194 18368 38200 18420
rect 38252 18368 38258 18420
rect 39298 18368 39304 18420
rect 39356 18368 39362 18420
rect 20487 18244 20760 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 21174 18164 21180 18216
rect 21232 18164 21238 18216
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18204 21419 18207
rect 21744 18204 21772 18368
rect 21818 18300 21824 18352
rect 21876 18340 21882 18352
rect 23952 18340 23980 18368
rect 26326 18340 26332 18352
rect 21876 18312 23980 18340
rect 25346 18312 26332 18340
rect 21876 18300 21882 18312
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 22388 18281 22416 18312
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18241 22431 18275
rect 22629 18275 22687 18281
rect 22629 18272 22641 18275
rect 22373 18235 22431 18241
rect 22480 18244 22641 18272
rect 22480 18204 22508 18244
rect 22629 18241 22641 18244
rect 22675 18241 22687 18275
rect 22629 18235 22687 18241
rect 23382 18232 23388 18284
rect 23440 18232 23446 18284
rect 23768 18272 23796 18312
rect 26326 18300 26332 18312
rect 26384 18340 26390 18352
rect 26694 18340 26700 18352
rect 26384 18312 26700 18340
rect 26384 18300 26390 18312
rect 26694 18300 26700 18312
rect 26752 18300 26758 18352
rect 27724 18312 28994 18340
rect 27724 18284 27752 18312
rect 23845 18275 23903 18281
rect 23845 18272 23857 18275
rect 23768 18244 23857 18272
rect 23845 18241 23857 18244
rect 23891 18241 23903 18275
rect 23845 18235 23903 18241
rect 26142 18232 26148 18284
rect 26200 18232 26206 18284
rect 27706 18232 27712 18284
rect 27764 18232 27770 18284
rect 28718 18232 28724 18284
rect 28776 18272 28782 18284
rect 28813 18275 28871 18281
rect 28813 18272 28825 18275
rect 28776 18244 28825 18272
rect 28776 18232 28782 18244
rect 28813 18241 28825 18244
rect 28859 18241 28871 18275
rect 28966 18272 28994 18312
rect 31846 18300 31852 18352
rect 31904 18340 31910 18352
rect 32582 18340 32588 18352
rect 31904 18312 32588 18340
rect 31904 18300 31910 18312
rect 32582 18300 32588 18312
rect 32640 18300 32646 18352
rect 29089 18275 29147 18281
rect 29089 18272 29101 18275
rect 28966 18244 29101 18272
rect 28813 18235 28871 18241
rect 29089 18241 29101 18244
rect 29135 18241 29147 18275
rect 29089 18235 29147 18241
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 36081 18275 36139 18281
rect 32088 18244 34100 18272
rect 32088 18232 32094 18244
rect 21407 18176 21772 18204
rect 22296 18176 22508 18204
rect 23400 18204 23428 18232
rect 34072 18216 34100 18244
rect 36081 18241 36093 18275
rect 36127 18272 36139 18275
rect 36188 18272 36216 18368
rect 38212 18340 38240 18368
rect 38212 18312 38318 18340
rect 36127 18244 36216 18272
rect 36127 18241 36139 18244
rect 36081 18235 36139 18241
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23400 18176 24133 18204
rect 21407 18173 21419 18176
rect 21361 18167 21419 18173
rect 21910 18136 21916 18148
rect 19720 18108 21916 18136
rect 21910 18096 21916 18108
rect 21968 18096 21974 18148
rect 22296 18145 22324 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 28994 18164 29000 18216
rect 29052 18164 29058 18216
rect 30926 18164 30932 18216
rect 30984 18204 30990 18216
rect 31478 18204 31484 18216
rect 30984 18176 31484 18204
rect 30984 18164 30990 18176
rect 31478 18164 31484 18176
rect 31536 18204 31542 18216
rect 32125 18207 32183 18213
rect 32125 18204 32137 18207
rect 31536 18176 32137 18204
rect 31536 18164 31542 18176
rect 32125 18173 32137 18176
rect 32171 18173 32183 18207
rect 32125 18167 32183 18173
rect 33594 18164 33600 18216
rect 33652 18164 33658 18216
rect 34054 18164 34060 18216
rect 34112 18204 34118 18216
rect 36354 18204 36360 18216
rect 34112 18176 36360 18204
rect 34112 18164 34118 18176
rect 36354 18164 36360 18176
rect 36412 18164 36418 18216
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 37553 18207 37611 18213
rect 37553 18204 37565 18207
rect 37516 18176 37565 18204
rect 37516 18164 37522 18176
rect 37553 18173 37565 18176
rect 37599 18173 37611 18207
rect 37553 18167 37611 18173
rect 37826 18164 37832 18216
rect 37884 18164 37890 18216
rect 22281 18139 22339 18145
rect 22281 18105 22293 18139
rect 22327 18105 22339 18139
rect 22281 18099 22339 18105
rect 23474 18068 23480 18080
rect 19628 18040 23480 18068
rect 19337 18031 19395 18037
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 26326 18028 26332 18080
rect 26384 18028 26390 18080
rect 1104 17978 45172 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 45172 17978
rect 1104 17904 45172 17926
rect 11517 17867 11575 17873
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 11698 17864 11704 17876
rect 11563 17836 11704 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22189 17867 22247 17873
rect 22189 17864 22201 17867
rect 22152 17836 22201 17864
rect 22152 17824 22158 17836
rect 22189 17833 22201 17836
rect 22235 17833 22247 17867
rect 22189 17827 22247 17833
rect 27706 17824 27712 17876
rect 27764 17824 27770 17876
rect 30926 17824 30932 17876
rect 30984 17824 30990 17876
rect 32214 17824 32220 17876
rect 32272 17864 32278 17876
rect 32769 17867 32827 17873
rect 32272 17836 32628 17864
rect 32272 17824 32278 17836
rect 6914 17756 6920 17808
rect 6972 17756 6978 17808
rect 16301 17799 16359 17805
rect 16301 17765 16313 17799
rect 16347 17796 16359 17799
rect 16347 17768 23888 17796
rect 16347 17765 16359 17768
rect 16301 17759 16359 17765
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 11054 17728 11060 17740
rect 9815 17700 11060 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 11054 17688 11060 17700
rect 11112 17728 11118 17740
rect 11514 17728 11520 17740
rect 11112 17700 11520 17728
rect 11112 17688 11118 17700
rect 11514 17688 11520 17700
rect 11572 17728 11578 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11572 17700 11621 17728
rect 11572 17688 11578 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12342 17728 12348 17740
rect 11931 17700 12348 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 21910 17688 21916 17740
rect 21968 17728 21974 17740
rect 21968 17700 22692 17728
rect 21968 17688 21974 17700
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15620 17632 16129 17660
rect 15620 17620 15626 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 22554 17620 22560 17672
rect 22612 17620 22618 17672
rect 22664 17660 22692 17700
rect 22738 17688 22744 17740
rect 22796 17688 22802 17740
rect 23658 17688 23664 17740
rect 23716 17688 23722 17740
rect 23676 17660 23704 17688
rect 22664 17632 23704 17660
rect 6641 17595 6699 17601
rect 6641 17561 6653 17595
rect 6687 17592 6699 17595
rect 7190 17592 7196 17604
rect 6687 17564 7196 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 10042 17552 10048 17604
rect 10100 17552 10106 17604
rect 10778 17552 10784 17604
rect 10836 17552 10842 17604
rect 23750 17592 23756 17604
rect 12268 17564 12374 17592
rect 13372 17564 23756 17592
rect 12268 17536 12296 17564
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 13372 17533 13400 17564
rect 23750 17552 23756 17564
rect 23808 17552 23814 17604
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 15654 17484 15660 17536
rect 15712 17524 15718 17536
rect 21818 17524 21824 17536
rect 15712 17496 21824 17524
rect 15712 17484 15718 17496
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 22646 17484 22652 17536
rect 22704 17484 22710 17536
rect 23860 17524 23888 17768
rect 23934 17688 23940 17740
rect 23992 17728 23998 17740
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 23992 17700 25973 17728
rect 23992 17688 23998 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 26237 17731 26295 17737
rect 26237 17697 26249 17731
rect 26283 17728 26295 17731
rect 26326 17728 26332 17740
rect 26283 17700 26332 17728
rect 26283 17697 26295 17700
rect 26237 17691 26295 17697
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 32398 17688 32404 17740
rect 32456 17688 32462 17740
rect 32600 17728 32628 17836
rect 32769 17833 32781 17867
rect 32815 17864 32827 17867
rect 33594 17864 33600 17876
rect 32815 17836 33600 17864
rect 32815 17833 32827 17836
rect 32769 17827 32827 17833
rect 33594 17824 33600 17836
rect 33652 17824 33658 17876
rect 32677 17731 32735 17737
rect 32677 17728 32689 17731
rect 32600 17700 32689 17728
rect 32677 17697 32689 17700
rect 32723 17697 32735 17731
rect 32677 17691 32735 17697
rect 33686 17688 33692 17740
rect 33744 17728 33750 17740
rect 34241 17731 34299 17737
rect 34241 17728 34253 17731
rect 33744 17700 34253 17728
rect 33744 17688 33750 17700
rect 34241 17697 34253 17700
rect 34287 17697 34299 17731
rect 34241 17691 34299 17697
rect 34514 17688 34520 17740
rect 34572 17688 34578 17740
rect 28902 17620 28908 17672
rect 28960 17620 28966 17672
rect 26694 17552 26700 17604
rect 26752 17552 26758 17604
rect 32122 17592 32128 17604
rect 31970 17564 32128 17592
rect 32122 17552 32128 17564
rect 32180 17592 32186 17604
rect 32858 17592 32864 17604
rect 32180 17564 32864 17592
rect 32180 17552 32186 17564
rect 32858 17552 32864 17564
rect 32916 17592 32922 17604
rect 32916 17564 33074 17592
rect 32916 17552 32922 17564
rect 35802 17552 35808 17604
rect 35860 17552 35866 17604
rect 27246 17524 27252 17536
rect 23860 17496 27252 17524
rect 27246 17484 27252 17496
rect 27304 17484 27310 17536
rect 28074 17484 28080 17536
rect 28132 17524 28138 17536
rect 28353 17527 28411 17533
rect 28353 17524 28365 17527
rect 28132 17496 28365 17524
rect 28132 17484 28138 17496
rect 28353 17493 28365 17496
rect 28399 17493 28411 17527
rect 28353 17487 28411 17493
rect 37093 17527 37151 17533
rect 37093 17493 37105 17527
rect 37139 17524 37151 17527
rect 37458 17524 37464 17536
rect 37139 17496 37464 17524
rect 37139 17493 37151 17496
rect 37093 17487 37151 17493
rect 37458 17484 37464 17496
rect 37516 17484 37522 17536
rect 1104 17434 45172 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 45172 17434
rect 1104 17360 45172 17382
rect 7098 17280 7104 17332
rect 7156 17280 7162 17332
rect 13265 17323 13323 17329
rect 10796 17292 11928 17320
rect 7116 17184 7144 17280
rect 10796 17264 10824 17292
rect 10778 17212 10784 17264
rect 10836 17212 10842 17264
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11480 17224 11805 17252
rect 11480 17212 11486 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11900 17252 11928 17292
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 15654 17320 15660 17332
rect 13311 17292 15660 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 19797 17323 19855 17329
rect 15795 17292 19380 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 12250 17252 12256 17264
rect 11900 17224 12256 17252
rect 11793 17215 11851 17221
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 15930 17252 15936 17264
rect 15396 17224 15936 17252
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 7116 17156 7481 17184
rect 7469 17153 7481 17156
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 11514 17144 11520 17196
rect 11572 17144 11578 17196
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15120 17116 15148 17147
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 15396 17193 15424 17224
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 19242 17212 19248 17264
rect 19300 17212 19306 17264
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 15470 17144 15476 17196
rect 15528 17144 15534 17196
rect 15838 17144 15844 17196
rect 15896 17144 15902 17196
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 16482 17184 16488 17196
rect 16071 17156 16488 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 19352 17193 19380 17292
rect 19797 17289 19809 17323
rect 19843 17289 19855 17323
rect 19797 17283 19855 17289
rect 19812 17252 19840 17283
rect 19978 17280 19984 17332
rect 20036 17280 20042 17332
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20441 17323 20499 17329
rect 20441 17320 20453 17323
rect 20404 17292 20453 17320
rect 20404 17280 20410 17292
rect 20441 17289 20453 17292
rect 20487 17289 20499 17323
rect 20441 17283 20499 17289
rect 22465 17323 22523 17329
rect 22465 17289 22477 17323
rect 22511 17320 22523 17323
rect 28721 17323 28779 17329
rect 22511 17292 28580 17320
rect 22511 17289 22523 17292
rect 22465 17283 22523 17289
rect 23198 17252 23204 17264
rect 19812 17224 23204 17252
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 26694 17212 26700 17264
rect 26752 17252 26758 17264
rect 27522 17252 27528 17264
rect 26752 17224 27528 17252
rect 26752 17212 26758 17224
rect 27522 17212 27528 17224
rect 27580 17252 27586 17264
rect 28552 17252 28580 17292
rect 28721 17289 28733 17323
rect 28767 17320 28779 17323
rect 28902 17320 28908 17332
rect 28767 17292 28908 17320
rect 28767 17289 28779 17292
rect 28721 17283 28779 17289
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 37826 17280 37832 17332
rect 37884 17320 37890 17332
rect 38105 17323 38163 17329
rect 38105 17320 38117 17323
rect 37884 17292 38117 17320
rect 37884 17280 37890 17292
rect 38105 17289 38117 17292
rect 38151 17289 38163 17323
rect 38105 17283 38163 17289
rect 39114 17280 39120 17332
rect 39172 17320 39178 17332
rect 40586 17320 40592 17332
rect 39172 17292 40592 17320
rect 39172 17280 39178 17292
rect 40586 17280 40592 17292
rect 40644 17280 40650 17332
rect 29641 17255 29699 17261
rect 29641 17252 29653 17255
rect 27580 17224 27738 17252
rect 28552 17224 29653 17252
rect 27580 17212 27586 17224
rect 29641 17221 29653 17224
rect 29687 17221 29699 17255
rect 30926 17252 30932 17264
rect 30866 17224 30932 17252
rect 29641 17215 29699 17221
rect 30926 17212 30932 17224
rect 30984 17252 30990 17264
rect 32122 17252 32128 17264
rect 30984 17224 32128 17252
rect 30984 17212 30990 17224
rect 32122 17212 32128 17224
rect 32180 17212 32186 17264
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 19800 17187 19858 17193
rect 19800 17153 19812 17187
rect 19846 17184 19858 17187
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19846 17156 20177 17184
rect 19846 17153 19858 17156
rect 19800 17147 19858 17153
rect 20165 17153 20177 17156
rect 20211 17184 20223 17187
rect 22370 17184 22376 17196
rect 20211 17156 22376 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 15120 17088 16160 17116
rect 16132 16992 16160 17088
rect 16850 17076 16856 17128
rect 16908 17076 16914 17128
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17116 17095 17119
rect 17586 17116 17592 17128
rect 17083 17088 17592 17116
rect 17083 17085 17095 17088
rect 17037 17079 17095 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17770 17076 17776 17128
rect 17828 17076 17834 17128
rect 17862 17076 17868 17128
rect 17920 17125 17926 17128
rect 17920 17119 17948 17125
rect 17936 17085 17948 17119
rect 17920 17079 17948 17085
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18690 17116 18696 17128
rect 18095 17088 18696 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 17920 17076 17926 17079
rect 16390 17008 16396 17060
rect 16448 17048 16454 17060
rect 17494 17048 17500 17060
rect 16448 17020 17500 17048
rect 16448 17008 16454 17020
rect 17494 17008 17500 17020
rect 17552 17008 17558 17060
rect 7282 16940 7288 16992
rect 7340 16940 7346 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 16025 16983 16083 16989
rect 16025 16980 16037 16983
rect 14332 16952 16037 16980
rect 14332 16940 14338 16952
rect 16025 16949 16037 16952
rect 16071 16949 16083 16983
rect 16025 16943 16083 16949
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 18432 16980 18460 17088
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 18984 17060 19012 17147
rect 19242 17076 19248 17128
rect 19300 17076 19306 17128
rect 18966 17008 18972 17060
rect 19024 17048 19030 17060
rect 19812 17048 19840 17147
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 38010 17144 38016 17196
rect 38068 17144 38074 17196
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17085 20499 17119
rect 20441 17079 20499 17085
rect 19024 17020 19840 17048
rect 20456 17048 20484 17079
rect 21818 17076 21824 17128
rect 21876 17076 21882 17128
rect 26973 17119 27031 17125
rect 26973 17085 26985 17119
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 22922 17048 22928 17060
rect 20456 17020 22928 17048
rect 19024 17008 19030 17020
rect 22922 17008 22928 17020
rect 22980 17008 22986 17060
rect 16172 16952 18460 16980
rect 18693 16983 18751 16989
rect 16172 16940 16178 16952
rect 18693 16949 18705 16983
rect 18739 16980 18751 16983
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18739 16952 19073 16980
rect 18739 16949 18751 16952
rect 18693 16943 18751 16949
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19061 16943 19119 16949
rect 19426 16940 19432 16992
rect 19484 16940 19490 16992
rect 20254 16940 20260 16992
rect 20312 16940 20318 16992
rect 26988 16980 27016 17079
rect 27246 17076 27252 17128
rect 27304 17076 27310 17128
rect 28902 17076 28908 17128
rect 28960 17116 28966 17128
rect 29365 17119 29423 17125
rect 29365 17116 29377 17119
rect 28960 17088 29377 17116
rect 28960 17076 28966 17088
rect 29365 17085 29377 17088
rect 29411 17085 29423 17119
rect 29365 17079 29423 17085
rect 34977 17119 35035 17125
rect 34977 17085 34989 17119
rect 35023 17116 35035 17119
rect 35434 17116 35440 17128
rect 35023 17088 35440 17116
rect 35023 17085 35035 17088
rect 34977 17079 35035 17085
rect 35434 17076 35440 17088
rect 35492 17076 35498 17128
rect 35345 17051 35403 17057
rect 35345 17017 35357 17051
rect 35391 17048 35403 17051
rect 44634 17048 44640 17060
rect 35391 17020 44640 17048
rect 35391 17017 35403 17020
rect 35345 17011 35403 17017
rect 44634 17008 44640 17020
rect 44692 17008 44698 17060
rect 27614 16980 27620 16992
rect 26988 16952 27620 16980
rect 27614 16940 27620 16952
rect 27672 16940 27678 16992
rect 31110 16940 31116 16992
rect 31168 16940 31174 16992
rect 35437 16983 35495 16989
rect 35437 16949 35449 16983
rect 35483 16980 35495 16983
rect 35894 16980 35900 16992
rect 35483 16952 35900 16980
rect 35483 16949 35495 16952
rect 35437 16943 35495 16949
rect 35894 16940 35900 16952
rect 35952 16940 35958 16992
rect 1104 16890 45172 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 45172 16890
rect 1104 16816 45172 16838
rect 15933 16779 15991 16785
rect 14752 16748 15700 16776
rect 7006 16600 7012 16652
rect 7064 16600 7070 16652
rect 7282 16600 7288 16652
rect 7340 16600 7346 16652
rect 8757 16643 8815 16649
rect 8757 16609 8769 16643
rect 8803 16640 8815 16643
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8803 16612 9137 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 14274 16600 14280 16652
rect 14332 16600 14338 16652
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 14752 16649 14780 16748
rect 15672 16708 15700 16748
rect 15933 16745 15945 16779
rect 15979 16776 15991 16779
rect 15979 16748 16804 16776
rect 15979 16745 15991 16748
rect 15933 16739 15991 16745
rect 16776 16708 16804 16748
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 16908 16748 17417 16776
rect 16908 16736 16914 16748
rect 17405 16745 17417 16748
rect 17451 16745 17463 16779
rect 17405 16739 17463 16745
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 17681 16779 17739 16785
rect 17681 16776 17693 16779
rect 17644 16748 17693 16776
rect 17644 16736 17650 16748
rect 17681 16745 17693 16748
rect 17727 16745 17739 16779
rect 17681 16739 17739 16745
rect 18782 16736 18788 16788
rect 18840 16736 18846 16788
rect 20254 16736 20260 16788
rect 20312 16736 20318 16788
rect 27522 16736 27528 16788
rect 27580 16736 27586 16788
rect 27880 16779 27938 16785
rect 27880 16745 27892 16779
rect 27926 16776 27938 16779
rect 28074 16776 28080 16788
rect 27926 16748 28080 16776
rect 27926 16745 27938 16748
rect 27880 16739 27938 16745
rect 28074 16736 28080 16748
rect 28132 16736 28138 16788
rect 35240 16779 35298 16785
rect 35240 16745 35252 16779
rect 35286 16776 35298 16779
rect 35986 16776 35992 16788
rect 35286 16748 35992 16776
rect 35286 16745 35298 16748
rect 35240 16739 35298 16745
rect 35986 16736 35992 16748
rect 36044 16736 36050 16788
rect 37080 16779 37138 16785
rect 37080 16745 37092 16779
rect 37126 16776 37138 16779
rect 37274 16776 37280 16788
rect 37126 16748 37280 16776
rect 37126 16745 37138 16748
rect 37080 16739 37138 16745
rect 37274 16736 37280 16748
rect 37332 16736 37338 16788
rect 20272 16708 20300 16736
rect 15672 16680 16252 16708
rect 16776 16680 20300 16708
rect 23124 16680 25268 16708
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14516 16612 14749 16640
rect 14516 16600 14522 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14826 16600 14832 16652
rect 14884 16640 14890 16652
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 14884 16612 15025 16640
rect 14884 16600 14890 16612
rect 15013 16609 15025 16612
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15335 16612 15885 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 14090 16532 14096 16584
rect 14148 16532 14154 16584
rect 15102 16532 15108 16584
rect 15160 16581 15166 16584
rect 15160 16575 15188 16581
rect 15176 16541 15188 16575
rect 15857 16572 15885 16612
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15988 16612 16037 16640
rect 15988 16600 15994 16612
rect 16025 16609 16037 16612
rect 16071 16609 16083 16643
rect 16025 16603 16083 16609
rect 16114 16600 16120 16652
rect 16172 16600 16178 16652
rect 16224 16640 16252 16680
rect 16390 16640 16396 16652
rect 16224 16612 16396 16640
rect 16132 16572 16160 16600
rect 16224 16581 16252 16612
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 16592 16612 17325 16640
rect 15857 16544 16160 16572
rect 16209 16575 16267 16581
rect 15160 16535 15188 16541
rect 16209 16541 16221 16575
rect 16255 16541 16267 16575
rect 16485 16575 16543 16581
rect 16485 16572 16497 16575
rect 16209 16535 16267 16541
rect 16316 16544 16497 16572
rect 15160 16532 15166 16535
rect 9674 16504 9680 16516
rect 8510 16476 9680 16504
rect 9674 16464 9680 16476
rect 9732 16504 9738 16516
rect 10778 16504 10784 16516
rect 9732 16476 10784 16504
rect 9732 16464 9738 16476
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 15838 16464 15844 16516
rect 15896 16504 15902 16516
rect 16316 16504 16344 16544
rect 16485 16541 16497 16544
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 16592 16504 16620 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 17494 16600 17500 16652
rect 17552 16600 17558 16652
rect 18233 16643 18291 16649
rect 18233 16609 18245 16643
rect 18279 16640 18291 16643
rect 18414 16640 18420 16652
rect 18279 16612 18420 16640
rect 18279 16609 18291 16612
rect 18233 16603 18291 16609
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 23124 16584 23152 16680
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23440 16612 23765 16640
rect 23440 16600 23446 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 25240 16640 25268 16680
rect 25406 16640 25412 16652
rect 23753 16603 23811 16609
rect 23860 16612 25176 16640
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 15896 16476 16344 16504
rect 16408 16476 16620 16504
rect 15896 16464 15902 16476
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 9769 16439 9827 16445
rect 9769 16436 9781 16439
rect 9548 16408 9781 16436
rect 9548 16396 9554 16408
rect 9769 16405 9781 16408
rect 9815 16405 9827 16439
rect 9769 16399 9827 16405
rect 15562 16396 15568 16448
rect 15620 16436 15626 16448
rect 16408 16445 16436 16476
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 15620 16408 16405 16436
rect 15620 16396 15626 16408
rect 16393 16405 16405 16408
rect 16439 16405 16451 16439
rect 16393 16399 16451 16405
rect 17126 16396 17132 16448
rect 17184 16436 17190 16448
rect 17604 16436 17632 16535
rect 18506 16532 18512 16584
rect 18564 16532 18570 16584
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16572 18843 16575
rect 18966 16572 18972 16584
rect 18831 16544 18972 16572
rect 18831 16541 18843 16544
rect 18785 16535 18843 16541
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 23106 16532 23112 16584
rect 23164 16532 23170 16584
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 23860 16581 23888 16612
rect 23661 16575 23719 16581
rect 23661 16572 23673 16575
rect 23624 16544 23673 16572
rect 23624 16532 23630 16544
rect 23661 16541 23673 16544
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16541 23903 16575
rect 23845 16535 23903 16541
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 24544 16544 24869 16572
rect 24544 16532 24550 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 24946 16532 24952 16584
rect 25004 16532 25010 16584
rect 25038 16532 25044 16584
rect 25096 16532 25102 16584
rect 23492 16504 23520 16532
rect 24581 16507 24639 16513
rect 24581 16504 24593 16507
rect 23492 16476 24593 16504
rect 24581 16473 24593 16476
rect 24627 16473 24639 16507
rect 25148 16504 25176 16612
rect 25240 16612 25412 16640
rect 25240 16581 25268 16612
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25332 16504 25360 16532
rect 25148 16476 25360 16504
rect 27540 16504 27568 16736
rect 31938 16668 31944 16720
rect 31996 16708 32002 16720
rect 32677 16711 32735 16717
rect 32677 16708 32689 16711
rect 31996 16680 32689 16708
rect 31996 16668 32002 16680
rect 32677 16677 32689 16680
rect 32723 16677 32735 16711
rect 32677 16671 32735 16677
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 29549 16643 29607 16649
rect 29549 16640 29561 16643
rect 27672 16612 29561 16640
rect 27672 16600 27678 16612
rect 28920 16584 28948 16612
rect 29549 16609 29561 16612
rect 29595 16609 29607 16643
rect 29549 16603 29607 16609
rect 32861 16643 32919 16649
rect 32861 16609 32873 16643
rect 32907 16640 32919 16643
rect 32907 16612 33172 16640
rect 32907 16609 32919 16612
rect 32861 16603 32919 16609
rect 28902 16532 28908 16584
rect 28960 16532 28966 16584
rect 29178 16572 29184 16584
rect 29026 16544 29184 16572
rect 29178 16532 29184 16544
rect 29236 16532 29242 16584
rect 31297 16575 31355 16581
rect 31297 16541 31309 16575
rect 31343 16572 31355 16575
rect 33042 16572 33048 16584
rect 31343 16544 33048 16572
rect 31343 16541 31355 16544
rect 31297 16535 31355 16541
rect 33042 16532 33048 16544
rect 33100 16532 33106 16584
rect 33144 16581 33172 16612
rect 34514 16600 34520 16652
rect 34572 16640 34578 16652
rect 34977 16643 35035 16649
rect 34977 16640 34989 16643
rect 34572 16612 34989 16640
rect 34572 16600 34578 16612
rect 34977 16609 34989 16612
rect 35023 16640 35035 16643
rect 36817 16643 36875 16649
rect 36817 16640 36829 16643
rect 35023 16612 36829 16640
rect 35023 16609 35035 16612
rect 34977 16603 35035 16609
rect 36817 16609 36829 16612
rect 36863 16640 36875 16643
rect 37458 16640 37464 16652
rect 36863 16612 37464 16640
rect 36863 16609 36875 16612
rect 36817 16603 36875 16609
rect 37458 16600 37464 16612
rect 37516 16600 37522 16652
rect 38565 16643 38623 16649
rect 38565 16609 38577 16643
rect 38611 16640 38623 16643
rect 39209 16643 39267 16649
rect 39209 16640 39221 16643
rect 38611 16612 39221 16640
rect 38611 16609 38623 16612
rect 38565 16603 38623 16609
rect 39209 16609 39221 16612
rect 39255 16609 39267 16643
rect 39209 16603 39267 16609
rect 33137 16575 33195 16581
rect 33137 16541 33149 16575
rect 33183 16541 33195 16575
rect 33137 16535 33195 16541
rect 38194 16532 38200 16584
rect 38252 16532 38258 16584
rect 44542 16532 44548 16584
rect 44600 16532 44606 16584
rect 28166 16504 28172 16516
rect 27540 16476 28172 16504
rect 24581 16467 24639 16473
rect 28166 16464 28172 16476
rect 28224 16464 28230 16516
rect 32401 16507 32459 16513
rect 32401 16504 32413 16507
rect 29196 16476 32413 16504
rect 17184 16408 17632 16436
rect 17184 16396 17190 16408
rect 18046 16396 18052 16448
rect 18104 16396 18110 16448
rect 18138 16396 18144 16448
rect 18196 16396 18202 16448
rect 18601 16439 18659 16445
rect 18601 16405 18613 16439
rect 18647 16436 18659 16439
rect 18690 16436 18696 16448
rect 18647 16408 18696 16436
rect 18647 16405 18659 16408
rect 18601 16399 18659 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 23658 16396 23664 16448
rect 23716 16436 23722 16448
rect 29196 16436 29224 16476
rect 32401 16473 32413 16476
rect 32447 16504 32459 16507
rect 36814 16504 36820 16516
rect 32447 16476 35480 16504
rect 36478 16476 36820 16504
rect 32447 16473 32459 16476
rect 32401 16467 32459 16473
rect 35452 16448 35480 16476
rect 36814 16464 36820 16476
rect 36872 16504 36878 16516
rect 36872 16476 37412 16504
rect 36872 16464 36878 16476
rect 23716 16408 29224 16436
rect 23716 16396 23722 16408
rect 29362 16396 29368 16448
rect 29420 16396 29426 16448
rect 32950 16396 32956 16448
rect 33008 16396 33014 16448
rect 35434 16396 35440 16448
rect 35492 16396 35498 16448
rect 36722 16396 36728 16448
rect 36780 16396 36786 16448
rect 37384 16436 37412 16476
rect 38212 16436 38240 16532
rect 37384 16408 38240 16436
rect 38378 16396 38384 16448
rect 38436 16436 38442 16448
rect 38657 16439 38715 16445
rect 38657 16436 38669 16439
rect 38436 16408 38669 16436
rect 38436 16396 38442 16408
rect 38657 16405 38669 16408
rect 38703 16405 38715 16439
rect 38657 16399 38715 16405
rect 44726 16396 44732 16448
rect 44784 16396 44790 16448
rect 1104 16346 45172 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 45172 16346
rect 1104 16272 45172 16294
rect 9674 16192 9680 16244
rect 9732 16192 9738 16244
rect 13446 16192 13452 16244
rect 13504 16192 13510 16244
rect 14090 16192 14096 16244
rect 14148 16232 14154 16244
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 14148 16204 14841 16232
rect 14148 16192 14154 16204
rect 14829 16201 14841 16204
rect 14875 16201 14887 16235
rect 14829 16195 14887 16201
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 15344 16204 15485 16232
rect 15344 16192 15350 16204
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 17034 16232 17040 16244
rect 15473 16195 15531 16201
rect 15580 16204 17040 16232
rect 9490 16124 9496 16176
rect 9548 16124 9554 16176
rect 9692 16164 9720 16192
rect 9692 16136 9982 16164
rect 14734 16124 14740 16176
rect 14792 16124 14798 16176
rect 14918 16124 14924 16176
rect 14976 16164 14982 16176
rect 15580 16164 15608 16204
rect 17034 16192 17040 16204
rect 17092 16232 17098 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17092 16204 17417 16232
rect 17092 16192 17098 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 19705 16235 19763 16241
rect 19705 16232 19717 16235
rect 19484 16204 19717 16232
rect 19484 16192 19490 16204
rect 19705 16201 19717 16204
rect 19751 16201 19763 16235
rect 22278 16232 22284 16244
rect 19705 16195 19763 16201
rect 22066 16204 22284 16232
rect 21913 16167 21971 16173
rect 14976 16136 15608 16164
rect 15948 16136 17356 16164
rect 14976 16124 14982 16136
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 7156 16000 7205 16028
rect 7156 15988 7162 16000
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 8128 16028 8156 16059
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14826 16096 14832 16108
rect 13964 16068 14832 16096
rect 13964 16056 13970 16068
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 15010 16056 15016 16108
rect 15068 16056 15074 16108
rect 15562 16096 15568 16108
rect 15120 16068 15568 16096
rect 7699 16000 8156 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8996 16000 9229 16028
rect 8996 15988 9002 16000
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 1578 15920 1584 15972
rect 1636 15960 1642 15972
rect 7469 15963 7527 15969
rect 7469 15960 7481 15963
rect 1636 15932 7481 15960
rect 1636 15920 1642 15932
rect 7469 15929 7481 15932
rect 7515 15929 7527 15963
rect 7469 15923 7527 15929
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 15120 15892 15148 16068
rect 15562 16056 15568 16068
rect 15620 16096 15626 16108
rect 15948 16105 15976 16136
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15620 16068 15669 16096
rect 15620 16056 15626 16068
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15933 16099 15991 16105
rect 15795 16068 15885 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 15857 16028 15885 16068
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16096 16083 16099
rect 16071 16068 16160 16096
rect 16071 16065 16083 16068
rect 16025 16059 16083 16065
rect 16132 16040 16160 16068
rect 16868 16040 16896 16136
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 15335 16000 15885 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 13596 15864 15148 15892
rect 15197 15895 15255 15901
rect 13596 15852 13602 15864
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15746 15892 15752 15904
rect 15243 15864 15752 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 15857 15892 15885 16000
rect 16114 15988 16120 16040
rect 16172 15988 16178 16040
rect 16850 15988 16856 16040
rect 16908 15988 16914 16040
rect 16022 15920 16028 15972
rect 16080 15960 16086 15972
rect 16960 15960 16988 16059
rect 17034 16056 17040 16108
rect 17092 16056 17098 16108
rect 17218 16056 17224 16108
rect 17276 16056 17282 16108
rect 17328 16105 17356 16136
rect 21913 16133 21925 16167
rect 21959 16164 21971 16167
rect 22066 16164 22094 16204
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 22370 16192 22376 16244
rect 22428 16192 22434 16244
rect 22922 16192 22928 16244
rect 22980 16192 22986 16244
rect 23198 16192 23204 16244
rect 23256 16232 23262 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 23256 16204 24317 16232
rect 23256 16192 23262 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 25130 16192 25136 16244
rect 25188 16192 25194 16244
rect 28166 16192 28172 16244
rect 28224 16232 28230 16244
rect 32950 16232 32956 16244
rect 28224 16204 29224 16232
rect 28224 16192 28230 16204
rect 22388 16164 22416 16192
rect 29196 16176 29224 16204
rect 32600 16204 32956 16232
rect 23014 16164 23020 16176
rect 21959 16136 22094 16164
rect 22296 16136 23020 16164
rect 21959 16133 21971 16136
rect 21913 16127 21971 16133
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17402 16056 17408 16108
rect 17460 16096 17466 16108
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 17460 16068 17601 16096
rect 17460 16056 17466 16068
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 17589 16059 17647 16065
rect 18690 16056 18696 16108
rect 18748 16096 18754 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 18748 16068 19441 16096
rect 18748 16056 18754 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 22296 16105 22324 16136
rect 23014 16124 23020 16136
rect 23072 16124 23078 16176
rect 23566 16164 23572 16176
rect 23216 16136 23572 16164
rect 23216 16108 23244 16136
rect 23566 16124 23572 16136
rect 23624 16164 23630 16176
rect 23845 16167 23903 16173
rect 23845 16164 23857 16167
rect 23624 16136 23857 16164
rect 23624 16124 23630 16136
rect 23845 16133 23857 16136
rect 23891 16164 23903 16167
rect 23891 16136 24900 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21140 16068 22109 16096
rect 21140 16056 21146 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16065 22339 16099
rect 22281 16059 22339 16065
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16096 22799 16099
rect 23109 16099 23167 16105
rect 22787 16068 22968 16096
rect 22787 16065 22799 16068
rect 22741 16059 22799 16065
rect 17862 15988 17868 16040
rect 17920 15988 17926 16040
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 16028 19763 16031
rect 22465 16031 22523 16037
rect 22465 16028 22477 16031
rect 19751 16000 20208 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 16080 15932 16988 15960
rect 17589 15963 17647 15969
rect 16080 15920 16086 15932
rect 17589 15929 17601 15963
rect 17635 15960 17647 15963
rect 17880 15960 17908 15988
rect 17635 15932 17908 15960
rect 17635 15929 17647 15932
rect 17589 15923 17647 15929
rect 20180 15904 20208 16000
rect 21836 16000 22477 16028
rect 21836 15972 21864 16000
rect 22465 15997 22477 16000
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22940 15972 22968 16068
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23124 16028 23152 16059
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 23382 16056 23388 16108
rect 23440 16056 23446 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23523 16068 23704 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23566 16028 23572 16040
rect 23124 16000 23572 16028
rect 23566 15988 23572 16000
rect 23624 15988 23630 16040
rect 21818 15920 21824 15972
rect 21876 15920 21882 15972
rect 22922 15920 22928 15972
rect 22980 15920 22986 15972
rect 23014 15920 23020 15972
rect 23072 15960 23078 15972
rect 23676 15960 23704 16068
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 24544 16000 24716 16028
rect 24544 15988 24550 16000
rect 23072 15932 23704 15960
rect 23072 15920 23078 15932
rect 23750 15920 23756 15972
rect 23808 15960 23814 15972
rect 24688 15960 24716 16000
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 24872 16037 24900 16136
rect 27890 16124 27896 16176
rect 27948 16124 27954 16176
rect 29178 16164 29184 16176
rect 29118 16136 29184 16164
rect 29178 16124 29184 16136
rect 29236 16164 29242 16176
rect 30926 16164 30932 16176
rect 29236 16136 30932 16164
rect 29236 16124 29242 16136
rect 30926 16124 30932 16136
rect 30984 16124 30990 16176
rect 32600 16173 32628 16204
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 35894 16192 35900 16244
rect 35952 16192 35958 16244
rect 35986 16192 35992 16244
rect 36044 16192 36050 16244
rect 36722 16192 36728 16244
rect 36780 16192 36786 16244
rect 38010 16192 38016 16244
rect 38068 16192 38074 16244
rect 41386 16204 41920 16232
rect 32585 16167 32643 16173
rect 32585 16133 32597 16167
rect 32631 16133 32643 16167
rect 32585 16127 32643 16133
rect 32858 16124 32864 16176
rect 32916 16164 32922 16176
rect 32916 16136 33074 16164
rect 32916 16124 32922 16136
rect 34146 16124 34152 16176
rect 34204 16124 34210 16176
rect 25314 16056 25320 16108
rect 25372 16096 25378 16108
rect 25372 16068 26096 16096
rect 25372 16056 25378 16068
rect 26068 16040 26096 16068
rect 27614 16056 27620 16108
rect 27672 16056 27678 16108
rect 29362 16056 29368 16108
rect 29420 16096 29426 16108
rect 30558 16096 30564 16108
rect 29420 16068 30564 16096
rect 29420 16056 29426 16068
rect 30558 16056 30564 16068
rect 30616 16056 30622 16108
rect 30745 16099 30803 16105
rect 30745 16065 30757 16099
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 15997 24915 16031
rect 24857 15991 24915 15997
rect 25406 15988 25412 16040
rect 25464 15988 25470 16040
rect 25501 16031 25559 16037
rect 25501 15997 25513 16031
rect 25547 15997 25559 16031
rect 25501 15991 25559 15997
rect 25516 15960 25544 15991
rect 25590 15988 25596 16040
rect 25648 15988 25654 16040
rect 26050 15988 26056 16040
rect 26108 15988 26114 16040
rect 23808 15932 24624 15960
rect 24688 15932 25544 15960
rect 30760 15960 30788 16059
rect 31110 16056 31116 16108
rect 31168 16056 31174 16108
rect 31202 16056 31208 16108
rect 31260 16096 31266 16108
rect 31662 16105 31668 16108
rect 31389 16099 31447 16105
rect 31389 16096 31401 16099
rect 31260 16068 31401 16096
rect 31260 16056 31266 16068
rect 31389 16065 31401 16068
rect 31435 16065 31447 16099
rect 31389 16059 31447 16065
rect 31658 16059 31668 16105
rect 31720 16096 31726 16108
rect 31720 16068 31758 16096
rect 31662 16056 31668 16059
rect 31720 16056 31726 16068
rect 32214 16056 32220 16108
rect 32272 16096 32278 16108
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 32272 16068 32321 16096
rect 32272 16056 32278 16068
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 35912 16096 35940 16192
rect 36173 16099 36231 16105
rect 36173 16096 36185 16099
rect 35912 16068 36185 16096
rect 32309 16059 32367 16065
rect 36173 16065 36185 16068
rect 36219 16065 36231 16099
rect 36740 16096 36768 16192
rect 37458 16124 37464 16176
rect 37516 16164 37522 16176
rect 41386 16164 41414 16204
rect 41892 16176 41920 16204
rect 37516 16136 41414 16164
rect 37516 16124 37522 16136
rect 41874 16124 41880 16176
rect 41932 16124 41938 16176
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 36740 16068 37289 16096
rect 36173 16059 36231 16065
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 37826 16056 37832 16108
rect 37884 16096 37890 16108
rect 38473 16099 38531 16105
rect 38473 16096 38485 16099
rect 37884 16068 38485 16096
rect 37884 16056 37890 16068
rect 38473 16065 38485 16068
rect 38519 16065 38531 16099
rect 38473 16059 38531 16065
rect 31128 16028 31156 16056
rect 31478 16028 31484 16040
rect 31128 16000 31484 16028
rect 31478 15988 31484 16000
rect 31536 15988 31542 16040
rect 33042 15988 33048 16040
rect 33100 16028 33106 16040
rect 33100 16000 35664 16028
rect 33100 15988 33106 16000
rect 30760 15932 31708 15960
rect 23808 15920 23814 15932
rect 16758 15892 16764 15904
rect 15857 15864 16764 15892
rect 16758 15852 16764 15864
rect 16816 15852 16822 15904
rect 17221 15895 17279 15901
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17770 15892 17776 15904
rect 17267 15864 17776 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 19518 15852 19524 15904
rect 19576 15852 19582 15904
rect 20162 15852 20168 15904
rect 20220 15852 20226 15904
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 22557 15895 22615 15901
rect 22557 15892 22569 15895
rect 21784 15864 22569 15892
rect 21784 15852 21790 15864
rect 22557 15861 22569 15864
rect 22603 15861 22615 15895
rect 22557 15855 22615 15861
rect 22649 15895 22707 15901
rect 22649 15861 22661 15895
rect 22695 15892 22707 15895
rect 23658 15892 23664 15904
rect 22695 15864 23664 15892
rect 22695 15861 22707 15864
rect 22649 15855 22707 15861
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 24121 15895 24179 15901
rect 24121 15861 24133 15895
rect 24167 15892 24179 15895
rect 24486 15892 24492 15904
rect 24167 15864 24492 15892
rect 24167 15861 24179 15864
rect 24121 15855 24179 15861
rect 24486 15852 24492 15864
rect 24544 15852 24550 15904
rect 24596 15892 24624 15932
rect 28994 15892 29000 15904
rect 24596 15864 29000 15892
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 29362 15852 29368 15904
rect 29420 15852 29426 15904
rect 30742 15852 30748 15904
rect 30800 15852 30806 15904
rect 31680 15901 31708 15932
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 31754 15892 31760 15904
rect 31711 15864 31760 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 31846 15852 31852 15904
rect 31904 15852 31910 15904
rect 34054 15852 34060 15904
rect 34112 15852 34118 15904
rect 35636 15901 35664 16000
rect 41598 15988 41604 16040
rect 41656 16028 41662 16040
rect 42981 16031 43039 16037
rect 42981 16028 42993 16031
rect 41656 16000 42993 16028
rect 41656 15988 41662 16000
rect 42981 15997 42993 16000
rect 43027 15997 43039 16031
rect 42981 15991 43039 15997
rect 43533 16031 43591 16037
rect 43533 15997 43545 16031
rect 43579 16028 43591 16031
rect 44358 16028 44364 16040
rect 43579 16000 44364 16028
rect 43579 15997 43591 16000
rect 43533 15991 43591 15997
rect 44358 15988 44364 16000
rect 44416 15988 44422 16040
rect 43806 15920 43812 15972
rect 43864 15920 43870 15972
rect 35621 15895 35679 15901
rect 35621 15861 35633 15895
rect 35667 15892 35679 15895
rect 35802 15892 35808 15904
rect 35667 15864 35808 15892
rect 35667 15861 35679 15864
rect 35621 15855 35679 15861
rect 35802 15852 35808 15864
rect 35860 15892 35866 15904
rect 37182 15892 37188 15904
rect 35860 15864 37188 15892
rect 35860 15852 35866 15864
rect 37182 15852 37188 15864
rect 37240 15852 37246 15904
rect 37918 15852 37924 15904
rect 37976 15852 37982 15904
rect 38378 15852 38384 15904
rect 38436 15852 38442 15904
rect 38562 15852 38568 15904
rect 38620 15892 38626 15904
rect 39758 15892 39764 15904
rect 38620 15864 39764 15892
rect 38620 15852 38626 15864
rect 39758 15852 39764 15864
rect 39816 15852 39822 15904
rect 42242 15852 42248 15904
rect 42300 15892 42306 15904
rect 42429 15895 42487 15901
rect 42429 15892 42441 15895
rect 42300 15864 42441 15892
rect 42300 15852 42306 15864
rect 42429 15861 42441 15864
rect 42475 15861 42487 15895
rect 42429 15855 42487 15861
rect 43990 15852 43996 15904
rect 44048 15852 44054 15904
rect 1104 15802 45172 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 45172 15802
rect 1104 15728 45172 15750
rect 8294 15648 8300 15700
rect 8352 15648 8358 15700
rect 10686 15648 10692 15700
rect 10744 15648 10750 15700
rect 14274 15688 14280 15700
rect 12636 15660 14280 15688
rect 8312 15552 8340 15648
rect 12636 15629 12664 15660
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 15102 15688 15108 15700
rect 14599 15660 15108 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 17862 15688 17868 15700
rect 15304 15660 17868 15688
rect 12621 15623 12679 15629
rect 12621 15589 12633 15623
rect 12667 15589 12679 15623
rect 12621 15583 12679 15589
rect 13538 15580 13544 15632
rect 13596 15620 13602 15632
rect 14185 15623 14243 15629
rect 13596 15592 13676 15620
rect 13596 15580 13602 15592
rect 9217 15555 9275 15561
rect 9217 15552 9229 15555
rect 8312 15524 9229 15552
rect 9217 15521 9229 15524
rect 9263 15521 9275 15555
rect 9217 15515 9275 15521
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 13170 15552 13176 15564
rect 12115 15524 13176 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 13648 15561 13676 15592
rect 14185 15589 14197 15623
rect 14231 15620 14243 15623
rect 15304 15620 15332 15660
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18046 15648 18052 15700
rect 18104 15648 18110 15700
rect 20530 15648 20536 15700
rect 20588 15648 20594 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21082 15688 21088 15700
rect 21039 15660 21088 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 21269 15691 21327 15697
rect 21269 15688 21281 15691
rect 21232 15660 21281 15688
rect 21232 15648 21238 15660
rect 21269 15657 21281 15660
rect 21315 15657 21327 15691
rect 21269 15651 21327 15657
rect 22462 15648 22468 15700
rect 22520 15688 22526 15700
rect 23014 15688 23020 15700
rect 22520 15660 23020 15688
rect 22520 15648 22526 15660
rect 15654 15620 15660 15632
rect 14231 15592 15332 15620
rect 15396 15592 15660 15620
rect 14231 15589 14243 15592
rect 14185 15583 14243 15589
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 13311 15524 13369 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13357 15521 13369 15524
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15552 14427 15555
rect 14918 15552 14924 15564
rect 14415 15524 14924 15552
rect 14415 15521 14427 15524
rect 14369 15515 14427 15521
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 15286 15512 15292 15564
rect 15344 15512 15350 15564
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8938 15484 8944 15496
rect 8444 15456 8944 15484
rect 8444 15444 8450 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 12158 15444 12164 15496
rect 12216 15493 12222 15496
rect 12216 15487 12265 15493
rect 12216 15453 12219 15487
rect 12253 15453 12265 15487
rect 12216 15447 12265 15453
rect 12216 15444 12222 15447
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 9674 15376 9680 15428
rect 9732 15376 9738 15428
rect 11422 15376 11428 15428
rect 11480 15376 11486 15428
rect 13556 15348 13584 15447
rect 13630 15376 13636 15428
rect 13688 15416 13694 15428
rect 13740 15416 13768 15447
rect 13814 15444 13820 15496
rect 13872 15444 13878 15496
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 13688 15388 13768 15416
rect 13688 15376 13694 15388
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14108 15416 14136 15447
rect 14056 15388 14136 15416
rect 14369 15419 14427 15425
rect 14056 15376 14062 15388
rect 14369 15385 14381 15419
rect 14415 15416 14427 15419
rect 14476 15416 14504 15447
rect 14415 15388 14504 15416
rect 14660 15416 14688 15447
rect 15194 15444 15200 15496
rect 15252 15444 15258 15496
rect 15396 15493 15424 15592
rect 15654 15580 15660 15592
rect 15712 15620 15718 15632
rect 18064 15620 18092 15648
rect 15712 15592 18092 15620
rect 19613 15623 19671 15629
rect 15712 15580 15718 15592
rect 19613 15589 19625 15623
rect 19659 15620 19671 15623
rect 20622 15620 20628 15632
rect 19659 15592 20628 15620
rect 19659 15589 19671 15592
rect 19613 15583 19671 15589
rect 20622 15580 20628 15592
rect 20680 15580 20686 15632
rect 21818 15620 21824 15632
rect 21468 15592 21824 15620
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 15746 15552 15752 15564
rect 15611 15524 15752 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 15746 15512 15752 15524
rect 15804 15552 15810 15564
rect 15804 15524 17540 15552
rect 15804 15512 15810 15524
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15838 15484 15844 15496
rect 15703 15456 15844 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15286 15416 15292 15428
rect 14660 15388 15292 15416
rect 14415 15385 14427 15388
rect 14369 15379 14427 15385
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 15488 15416 15516 15447
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16672 15465 16730 15471
rect 16040 15416 16068 15444
rect 16672 15431 16684 15465
rect 16718 15431 16730 15465
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 16872 15487 16930 15493
rect 16872 15453 16884 15487
rect 16918 15484 16930 15487
rect 17402 15484 17408 15496
rect 16918 15456 17408 15484
rect 16918 15453 16930 15456
rect 16872 15447 16930 15453
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 17512 15484 17540 15524
rect 17586 15512 17592 15564
rect 17644 15552 17650 15564
rect 17644 15524 21036 15552
rect 17644 15512 17650 15524
rect 19889 15487 19947 15493
rect 19889 15484 19901 15487
rect 17512 15456 18184 15484
rect 16672 15428 16730 15431
rect 15488 15388 16068 15416
rect 16666 15376 16672 15428
rect 16724 15376 16730 15428
rect 16776 15416 16804 15444
rect 18156 15428 18184 15456
rect 18340 15456 19901 15484
rect 16955 15419 17013 15425
rect 16955 15416 16967 15419
rect 16776 15388 16967 15416
rect 16955 15385 16967 15388
rect 17001 15416 17013 15419
rect 17001 15388 17540 15416
rect 17001 15385 17013 15388
rect 16955 15379 17013 15385
rect 14642 15348 14648 15360
rect 13556 15320 14648 15348
rect 14642 15308 14648 15320
rect 14700 15348 14706 15360
rect 16761 15351 16819 15357
rect 16761 15348 16773 15351
rect 14700 15320 16773 15348
rect 14700 15308 14706 15320
rect 16761 15317 16773 15320
rect 16807 15348 16819 15351
rect 17402 15348 17408 15360
rect 16807 15320 17408 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17512 15348 17540 15388
rect 18138 15376 18144 15428
rect 18196 15376 18202 15428
rect 18340 15360 18368 15456
rect 19889 15453 19901 15456
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 20487 15456 20668 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 20640 15416 20668 15456
rect 20714 15444 20720 15496
rect 20772 15444 20778 15496
rect 21008 15493 21036 15524
rect 21468 15493 21496 15592
rect 21818 15580 21824 15592
rect 21876 15580 21882 15632
rect 22005 15623 22063 15629
rect 22005 15589 22017 15623
rect 22051 15620 22063 15623
rect 22738 15620 22744 15632
rect 22051 15592 22744 15620
rect 22051 15589 22063 15592
rect 22005 15583 22063 15589
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 21634 15512 21640 15564
rect 21692 15512 21698 15564
rect 21726 15512 21732 15564
rect 21784 15512 21790 15564
rect 21836 15552 21864 15580
rect 22370 15552 22376 15564
rect 21836 15524 22376 15552
rect 22370 15512 22376 15524
rect 22428 15512 22434 15564
rect 22940 15552 22968 15660
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 23106 15648 23112 15700
rect 23164 15688 23170 15700
rect 23164 15660 23888 15688
rect 23164 15648 23170 15660
rect 23860 15552 23888 15660
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 24213 15691 24271 15697
rect 24213 15688 24225 15691
rect 24084 15660 24225 15688
rect 24084 15648 24090 15660
rect 24213 15657 24225 15660
rect 24259 15657 24271 15691
rect 24213 15651 24271 15657
rect 24302 15648 24308 15700
rect 24360 15688 24366 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 24360 15660 24409 15688
rect 24360 15648 24366 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 24397 15651 24455 15657
rect 24670 15648 24676 15700
rect 24728 15648 24734 15700
rect 25038 15648 25044 15700
rect 25096 15688 25102 15700
rect 25317 15691 25375 15697
rect 25317 15688 25329 15691
rect 25096 15660 25329 15688
rect 25096 15648 25102 15660
rect 25317 15657 25329 15660
rect 25363 15657 25375 15691
rect 25317 15651 25375 15657
rect 26510 15648 26516 15700
rect 26568 15688 26574 15700
rect 27157 15691 27215 15697
rect 27157 15688 27169 15691
rect 26568 15660 27169 15688
rect 26568 15648 26574 15660
rect 27157 15657 27169 15660
rect 27203 15657 27215 15691
rect 27157 15651 27215 15657
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 30006 15697 30012 15700
rect 29963 15691 30012 15697
rect 29963 15688 29975 15691
rect 29052 15660 29975 15688
rect 29052 15648 29058 15660
rect 29963 15657 29975 15660
rect 30009 15657 30012 15691
rect 29963 15651 30012 15657
rect 30006 15648 30012 15651
rect 30064 15648 30070 15700
rect 30558 15648 30564 15700
rect 30616 15648 30622 15700
rect 34054 15648 34060 15700
rect 34112 15648 34118 15700
rect 37458 15688 37464 15700
rect 35820 15660 37464 15688
rect 24688 15620 24716 15648
rect 25961 15623 26019 15629
rect 25961 15620 25973 15623
rect 24688 15592 25973 15620
rect 23937 15555 23995 15561
rect 23937 15552 23949 15555
rect 22940 15524 23244 15552
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15484 21235 15487
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 21223 15456 21465 15484
rect 21223 15453 21235 15456
rect 21177 15447 21235 15453
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 20806 15416 20812 15428
rect 19352 15388 20576 15416
rect 20640 15388 20812 15416
rect 19352 15360 19380 15388
rect 18322 15348 18328 15360
rect 17512 15320 18328 15348
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 19334 15308 19340 15360
rect 19392 15308 19398 15360
rect 19702 15308 19708 15360
rect 19760 15348 19766 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19760 15320 19809 15348
rect 19760 15308 19766 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 19978 15308 19984 15360
rect 20036 15308 20042 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20165 15351 20223 15357
rect 20165 15348 20177 15351
rect 20128 15320 20177 15348
rect 20128 15308 20134 15320
rect 20165 15317 20177 15320
rect 20211 15317 20223 15351
rect 20548 15348 20576 15388
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 20901 15419 20959 15425
rect 20901 15385 20913 15419
rect 20947 15416 20959 15419
rect 21560 15416 21588 15447
rect 21910 15444 21916 15496
rect 21968 15444 21974 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 22152 15456 22201 15484
rect 22152 15444 22158 15456
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 22462 15484 22468 15496
rect 22189 15447 22247 15453
rect 22296 15456 22468 15484
rect 20947 15388 21588 15416
rect 20947 15385 20959 15388
rect 20901 15379 20959 15385
rect 21818 15376 21824 15428
rect 21876 15416 21882 15428
rect 22296 15425 22324 15456
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 22554 15444 22560 15496
rect 22612 15444 22618 15496
rect 22646 15444 22652 15496
rect 22704 15444 22710 15496
rect 22833 15487 22891 15493
rect 22833 15486 22845 15487
rect 22756 15458 22845 15486
rect 22281 15419 22339 15425
rect 22281 15416 22293 15419
rect 21876 15388 22293 15416
rect 21876 15376 21882 15388
rect 22281 15385 22293 15388
rect 22327 15385 22339 15419
rect 22281 15379 22339 15385
rect 22373 15419 22431 15425
rect 22373 15385 22385 15419
rect 22419 15416 22431 15419
rect 22664 15416 22692 15444
rect 22419 15388 22692 15416
rect 22419 15385 22431 15388
rect 22373 15379 22431 15385
rect 22756 15360 22784 15458
rect 22833 15453 22845 15458
rect 22879 15453 22891 15487
rect 22833 15447 22891 15453
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 22940 15360 22968 15447
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23216 15493 23244 15524
rect 23308 15524 23612 15552
rect 23860 15524 23949 15552
rect 23308 15493 23336 15524
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 23072 15456 23121 15484
rect 23072 15444 23078 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 23382 15376 23388 15428
rect 23440 15376 23446 15428
rect 23584 15416 23612 15524
rect 23937 15521 23949 15524
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 24949 15555 25007 15561
rect 24949 15552 24961 15555
rect 24176 15524 24961 15552
rect 24176 15512 24182 15524
rect 24949 15521 24961 15524
rect 24995 15521 25007 15555
rect 24949 15515 25007 15521
rect 23750 15444 23756 15496
rect 23808 15444 23814 15496
rect 25424 15493 25452 15592
rect 25961 15589 25973 15592
rect 26007 15589 26019 15623
rect 25961 15583 26019 15589
rect 30101 15623 30159 15629
rect 30101 15589 30113 15623
rect 30147 15589 30159 15623
rect 30576 15620 30604 15648
rect 31662 15620 31668 15632
rect 30576 15592 31668 15620
rect 30101 15583 30159 15589
rect 25866 15512 25872 15564
rect 25924 15552 25930 15564
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 25924 15524 26525 15552
rect 25924 15512 25930 15524
rect 26513 15521 26525 15524
rect 26559 15521 26571 15555
rect 26513 15515 26571 15521
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 27249 15555 27307 15561
rect 27249 15552 27261 15555
rect 26844 15524 27261 15552
rect 26844 15512 26850 15524
rect 27249 15521 27261 15524
rect 27295 15521 27307 15555
rect 27249 15515 27307 15521
rect 29638 15512 29644 15564
rect 29696 15552 29702 15564
rect 30116 15552 30144 15583
rect 31662 15580 31668 15592
rect 31720 15620 31726 15632
rect 31720 15592 32260 15620
rect 31720 15580 31726 15592
rect 29696 15524 30144 15552
rect 30193 15555 30251 15561
rect 29696 15512 29702 15524
rect 30193 15521 30205 15555
rect 30239 15552 30251 15555
rect 31573 15555 31631 15561
rect 31573 15552 31585 15555
rect 30239 15524 30512 15552
rect 30239 15521 30251 15524
rect 30193 15515 30251 15521
rect 30484 15496 30512 15524
rect 31312 15524 31585 15552
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 24029 15487 24087 15493
rect 24029 15453 24041 15487
rect 24075 15484 24087 15487
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24075 15456 24624 15484
rect 24075 15453 24087 15456
rect 24029 15447 24087 15453
rect 23860 15416 23888 15447
rect 24486 15416 24492 15428
rect 23584 15388 24492 15416
rect 24486 15376 24492 15388
rect 24544 15376 24550 15428
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 20548 15320 22661 15348
rect 20165 15311 20223 15317
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 22738 15308 22744 15360
rect 22796 15308 22802 15360
rect 22922 15308 22928 15360
rect 22980 15348 22986 15360
rect 23842 15348 23848 15360
rect 22980 15320 23848 15348
rect 22980 15308 22986 15320
rect 23842 15308 23848 15320
rect 23900 15348 23906 15360
rect 24118 15348 24124 15360
rect 23900 15320 24124 15348
rect 23900 15308 23906 15320
rect 24118 15308 24124 15320
rect 24176 15308 24182 15360
rect 24596 15348 24624 15456
rect 24688 15456 25237 15484
rect 24688 15428 24716 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 29362 15444 29368 15496
rect 29420 15484 29426 15496
rect 29825 15487 29883 15493
rect 29825 15484 29837 15487
rect 29420 15456 29837 15484
rect 29420 15444 29426 15456
rect 29825 15453 29837 15456
rect 29871 15484 29883 15487
rect 30282 15484 30288 15496
rect 29871 15456 30288 15484
rect 29871 15453 29883 15456
rect 29825 15447 29883 15453
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 30466 15444 30472 15496
rect 30524 15444 30530 15496
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15484 31079 15487
rect 31202 15484 31208 15496
rect 31067 15456 31208 15484
rect 31067 15453 31079 15456
rect 31021 15447 31079 15453
rect 31202 15444 31208 15456
rect 31260 15444 31266 15496
rect 31312 15493 31340 15524
rect 31573 15521 31585 15524
rect 31619 15521 31631 15555
rect 31573 15515 31631 15521
rect 31297 15487 31355 15493
rect 31297 15453 31309 15487
rect 31343 15453 31355 15487
rect 31297 15447 31355 15453
rect 31478 15444 31484 15496
rect 31536 15444 31542 15496
rect 31754 15444 31760 15496
rect 31812 15444 31818 15496
rect 32232 15493 32260 15592
rect 34072 15552 34100 15648
rect 35820 15629 35848 15660
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 37918 15688 37924 15700
rect 37660 15660 37924 15688
rect 35805 15623 35863 15629
rect 35805 15589 35817 15623
rect 35851 15589 35863 15623
rect 35805 15583 35863 15589
rect 34701 15555 34759 15561
rect 34701 15552 34713 15555
rect 34072 15524 34713 15552
rect 34701 15521 34713 15524
rect 34747 15521 34759 15555
rect 34701 15515 34759 15521
rect 35989 15555 36047 15561
rect 35989 15521 36001 15555
rect 36035 15521 36047 15555
rect 35989 15515 36047 15521
rect 37461 15555 37519 15561
rect 37461 15521 37473 15555
rect 37507 15552 37519 15555
rect 37660 15552 37688 15660
rect 37918 15648 37924 15660
rect 37976 15648 37982 15700
rect 41598 15648 41604 15700
rect 41656 15648 41662 15700
rect 43625 15691 43683 15697
rect 43625 15657 43637 15691
rect 43671 15688 43683 15691
rect 43806 15688 43812 15700
rect 43671 15660 43812 15688
rect 43671 15657 43683 15660
rect 43625 15651 43683 15657
rect 43806 15648 43812 15660
rect 43864 15648 43870 15700
rect 37507 15524 37688 15552
rect 37752 15592 39896 15620
rect 37507 15521 37519 15524
rect 37461 15515 37519 15521
rect 32033 15487 32091 15493
rect 32033 15453 32045 15487
rect 32079 15453 32091 15487
rect 32033 15447 32091 15453
rect 32217 15487 32275 15493
rect 32217 15453 32229 15487
rect 32263 15453 32275 15487
rect 36004 15484 36032 15515
rect 37752 15496 37780 15592
rect 39114 15512 39120 15564
rect 39172 15512 39178 15564
rect 39868 15561 39896 15592
rect 39853 15555 39911 15561
rect 39853 15521 39865 15555
rect 39899 15552 39911 15555
rect 40678 15552 40684 15564
rect 39899 15524 40684 15552
rect 39899 15521 39911 15524
rect 39853 15515 39911 15521
rect 40678 15512 40684 15524
rect 40736 15552 40742 15564
rect 41877 15555 41935 15561
rect 41877 15552 41889 15555
rect 40736 15524 41889 15552
rect 40736 15512 40742 15524
rect 41877 15521 41889 15524
rect 41923 15521 41935 15555
rect 41877 15515 41935 15521
rect 42153 15555 42211 15561
rect 42153 15521 42165 15555
rect 42199 15552 42211 15555
rect 42242 15552 42248 15564
rect 42199 15524 42248 15552
rect 42199 15521 42211 15524
rect 42153 15515 42211 15521
rect 42242 15512 42248 15524
rect 42300 15512 42306 15564
rect 32217 15447 32275 15453
rect 32416 15456 36032 15484
rect 24670 15376 24676 15428
rect 24728 15376 24734 15428
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 24946 15416 24952 15428
rect 24811 15388 24952 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 24946 15376 24952 15388
rect 25004 15416 25010 15428
rect 26789 15419 26847 15425
rect 26789 15416 26801 15419
rect 25004 15388 26801 15416
rect 25004 15376 25010 15388
rect 26789 15385 26801 15388
rect 26835 15385 26847 15419
rect 31570 15416 31576 15428
rect 26789 15379 26847 15385
rect 30484 15388 31576 15416
rect 24857 15351 24915 15357
rect 24857 15348 24869 15351
rect 24596 15320 24869 15348
rect 24857 15317 24869 15320
rect 24903 15348 24915 15351
rect 25130 15348 25136 15360
rect 24903 15320 25136 15348
rect 24903 15317 24915 15320
rect 24857 15311 24915 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 26326 15308 26332 15360
rect 26384 15308 26390 15360
rect 26421 15351 26479 15357
rect 26421 15317 26433 15351
rect 26467 15348 26479 15351
rect 26878 15348 26884 15360
rect 26467 15320 26884 15348
rect 26467 15317 26479 15320
rect 26421 15311 26479 15317
rect 26878 15308 26884 15320
rect 26936 15308 26942 15360
rect 30484 15357 30512 15388
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 30469 15351 30527 15357
rect 30469 15317 30481 15351
rect 30515 15317 30527 15351
rect 30469 15311 30527 15317
rect 30558 15308 30564 15360
rect 30616 15348 30622 15360
rect 30837 15351 30895 15357
rect 30837 15348 30849 15351
rect 30616 15320 30849 15348
rect 30616 15308 30622 15320
rect 30837 15317 30849 15320
rect 30883 15317 30895 15351
rect 31772 15348 31800 15444
rect 32048 15416 32076 15447
rect 32306 15416 32312 15428
rect 32048 15388 32312 15416
rect 32306 15376 32312 15388
rect 32364 15376 32370 15428
rect 32416 15348 32444 15456
rect 37734 15444 37740 15496
rect 37792 15444 37798 15496
rect 39485 15487 39543 15493
rect 38488 15456 39068 15484
rect 35434 15376 35440 15428
rect 35492 15376 35498 15428
rect 36814 15376 36820 15428
rect 36872 15376 36878 15428
rect 31772 15320 32444 15348
rect 30837 15311 30895 15317
rect 35342 15308 35348 15360
rect 35400 15308 35406 15360
rect 35894 15308 35900 15360
rect 35952 15308 35958 15360
rect 38488 15357 38516 15456
rect 38654 15425 38660 15428
rect 38632 15419 38660 15425
rect 38632 15385 38644 15419
rect 38632 15379 38660 15385
rect 38654 15376 38660 15379
rect 38712 15376 38718 15428
rect 39040 15416 39068 15456
rect 39485 15453 39497 15487
rect 39531 15453 39543 15487
rect 39485 15447 39543 15453
rect 39500 15416 39528 15447
rect 40129 15419 40187 15425
rect 40129 15416 40141 15419
rect 39040 15388 39528 15416
rect 39684 15388 40141 15416
rect 38473 15351 38531 15357
rect 38473 15317 38485 15351
rect 38519 15317 38531 15351
rect 38473 15311 38531 15317
rect 38746 15308 38752 15360
rect 38804 15308 38810 15360
rect 38841 15351 38899 15357
rect 38841 15317 38853 15351
rect 38887 15348 38899 15351
rect 39022 15348 39028 15360
rect 38887 15320 39028 15348
rect 38887 15317 38899 15320
rect 38841 15311 38899 15317
rect 39022 15308 39028 15320
rect 39080 15308 39086 15360
rect 39684 15357 39712 15388
rect 40129 15385 40141 15388
rect 40175 15385 40187 15419
rect 41354 15388 42642 15416
rect 40129 15379 40187 15385
rect 39669 15351 39727 15357
rect 39669 15317 39681 15351
rect 39715 15317 39727 15351
rect 39669 15311 39727 15317
rect 39758 15308 39764 15360
rect 39816 15348 39822 15360
rect 41432 15348 41460 15388
rect 39816 15320 41460 15348
rect 39816 15308 39822 15320
rect 1104 15258 45172 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 45172 15258
rect 1104 15184 45172 15206
rect 12158 15104 12164 15156
rect 12216 15104 12222 15156
rect 12713 15147 12771 15153
rect 12713 15113 12725 15147
rect 12759 15144 12771 15147
rect 13078 15144 13084 15156
rect 12759 15116 13084 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13170 15104 13176 15156
rect 13228 15144 13234 15156
rect 13228 15116 13952 15144
rect 13228 15104 13234 15116
rect 13446 15076 13452 15088
rect 10152 15048 13452 15076
rect 10152 15020 10180 15048
rect 13446 15036 13452 15048
rect 13504 15036 13510 15088
rect 13814 15036 13820 15088
rect 13872 15036 13878 15088
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 8386 15008 8392 15020
rect 7064 14980 8392 15008
rect 7064 14968 7070 14980
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 8812 14912 10793 14940
rect 8812 14900 8818 14912
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 11716 14940 11744 14971
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12158 15008 12164 15020
rect 12023 14980 12164 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 12308 14980 12357 15008
rect 12308 14968 12314 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 13170 15017 13176 15020
rect 12989 15014 13047 15017
rect 12912 15011 13047 15014
rect 12912 14986 13001 15011
rect 11716 14912 12434 14940
rect 10781 14903 10839 14909
rect 10226 14764 10232 14816
rect 10284 14764 10290 14816
rect 12406 14804 12434 14912
rect 12912 14872 12940 14986
rect 12989 14977 13001 14986
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13167 14971 13176 15017
rect 13228 15008 13234 15020
rect 13228 14980 13267 15008
rect 13170 14968 13176 14971
rect 13228 14968 13234 14980
rect 13832 14940 13860 15036
rect 13924 15017 13952 15116
rect 14458 15104 14464 15156
rect 14516 15104 14522 15156
rect 14550 15104 14556 15156
rect 14608 15104 14614 15156
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 16945 15147 17003 15153
rect 15252 15116 16344 15144
rect 15252 15104 15258 15116
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 13194 14912 13860 14940
rect 13924 14940 13952 14971
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 15008 14427 15011
rect 14476 15008 14504 15104
rect 16316 15088 16344 15116
rect 16945 15113 16957 15147
rect 16991 15144 17003 15147
rect 17034 15144 17040 15156
rect 16991 15116 17040 15144
rect 16991 15113 17003 15116
rect 16945 15107 17003 15113
rect 17034 15104 17040 15116
rect 17092 15144 17098 15156
rect 17310 15144 17316 15156
rect 17092 15116 17316 15144
rect 17092 15104 17098 15116
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 18506 15144 18512 15156
rect 18003 15116 18512 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 18598 15104 18604 15156
rect 18656 15144 18662 15156
rect 20533 15147 20591 15153
rect 18656 15116 20484 15144
rect 18656 15104 18662 15116
rect 16298 15036 16304 15088
rect 16356 15036 16362 15088
rect 16853 15079 16911 15085
rect 16853 15045 16865 15079
rect 16899 15076 16911 15079
rect 17494 15076 17500 15088
rect 16899 15048 17500 15076
rect 16899 15045 16911 15048
rect 16853 15039 16911 15045
rect 17494 15036 17500 15048
rect 17552 15076 17558 15088
rect 18046 15076 18052 15088
rect 17552 15048 18052 15076
rect 17552 15036 17558 15048
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 19797 15079 19855 15085
rect 19797 15045 19809 15079
rect 19843 15076 19855 15079
rect 20456 15076 20484 15116
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20806 15144 20812 15156
rect 20579 15116 20812 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20806 15104 20812 15116
rect 20864 15144 20870 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20864 15116 20913 15144
rect 20864 15104 20870 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22612 15116 22661 15144
rect 22612 15104 22618 15116
rect 22649 15113 22661 15116
rect 22695 15113 22707 15147
rect 22649 15107 22707 15113
rect 22738 15104 22744 15156
rect 22796 15144 22802 15156
rect 23658 15144 23664 15156
rect 22796 15116 23664 15144
rect 22796 15104 22802 15116
rect 23658 15104 23664 15116
rect 23716 15144 23722 15156
rect 25593 15147 25651 15153
rect 25593 15144 25605 15147
rect 23716 15116 25605 15144
rect 23716 15104 23722 15116
rect 25593 15113 25605 15116
rect 25639 15113 25651 15147
rect 25593 15107 25651 15113
rect 26973 15147 27031 15153
rect 26973 15113 26985 15147
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 19843 15048 20300 15076
rect 20456 15048 21128 15076
rect 19843 15045 19855 15048
rect 19797 15039 19855 15045
rect 14415 14980 14504 15008
rect 14415 14977 14427 14980
rect 14369 14971 14427 14977
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16666 15008 16672 15020
rect 15804 14980 16672 15008
rect 15804 14968 15810 14980
rect 16666 14968 16672 14980
rect 16724 15008 16730 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16724 14980 16773 15008
rect 16724 14968 16730 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17589 15011 17647 15017
rect 17589 15008 17601 15011
rect 17267 14980 17601 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17589 14977 17601 14980
rect 17635 15008 17647 15011
rect 18506 15008 18512 15020
rect 17635 14980 18512 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 18656 14980 19625 15008
rect 18656 14968 18662 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 19978 15008 19984 15020
rect 19613 14971 19671 14977
rect 19720 14980 19984 15008
rect 16942 14940 16948 14952
rect 13924 14912 16948 14940
rect 13194 14881 13222 14912
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17497 14943 17555 14949
rect 17497 14940 17509 14943
rect 17331 14912 17509 14940
rect 13173 14875 13231 14881
rect 12912 14844 13124 14872
rect 12894 14804 12900 14816
rect 12406 14776 12900 14804
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13096 14804 13124 14844
rect 13173 14841 13185 14875
rect 13219 14841 13231 14875
rect 13173 14835 13231 14841
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 14185 14875 14243 14881
rect 14185 14872 14197 14875
rect 13872 14844 14197 14872
rect 13872 14832 13878 14844
rect 14185 14841 14197 14844
rect 14231 14841 14243 14875
rect 14185 14835 14243 14841
rect 14274 14832 14280 14884
rect 14332 14832 14338 14884
rect 14366 14804 14372 14816
rect 13096 14776 14372 14804
rect 14366 14764 14372 14776
rect 14424 14804 14430 14816
rect 15562 14804 15568 14816
rect 14424 14776 15568 14804
rect 14424 14764 14430 14776
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17034 14804 17040 14816
rect 16816 14776 17040 14804
rect 16816 14764 16822 14776
rect 17034 14764 17040 14776
rect 17092 14804 17098 14816
rect 17129 14807 17187 14813
rect 17129 14804 17141 14807
rect 17092 14776 17141 14804
rect 17092 14764 17098 14776
rect 17129 14773 17141 14776
rect 17175 14773 17187 14807
rect 17129 14767 17187 14773
rect 17221 14807 17279 14813
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17331 14804 17359 14912
rect 17497 14909 17509 14912
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 17678 14900 17684 14952
rect 17736 14900 17742 14952
rect 17770 14900 17776 14952
rect 17828 14900 17834 14952
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14940 19487 14943
rect 19720 14940 19748 14980
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20162 14968 20168 15020
rect 20220 14968 20226 15020
rect 20272 15008 20300 15048
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20272 14980 20453 15008
rect 20441 14977 20453 14980
rect 20487 15008 20499 15011
rect 20530 15008 20536 15020
rect 20487 14980 20536 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20680 14980 20729 15008
rect 20680 14968 20686 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 20806 14968 20812 15020
rect 20864 14968 20870 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21100 15008 21128 15048
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 23293 15079 23351 15085
rect 23293 15076 23305 15079
rect 21968 15048 23305 15076
rect 21968 15036 21974 15048
rect 23293 15045 23305 15048
rect 23339 15045 23351 15079
rect 23474 15076 23480 15088
rect 23293 15039 23351 15045
rect 23400 15048 23480 15076
rect 21100 14980 21956 15008
rect 19475 14912 19748 14940
rect 19889 14943 19947 14949
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 19889 14909 19901 14943
rect 19935 14940 19947 14943
rect 20070 14940 20076 14952
rect 19935 14912 20076 14940
rect 19935 14909 19947 14912
rect 19889 14903 19947 14909
rect 19150 14832 19156 14884
rect 19208 14872 19214 14884
rect 19352 14872 19380 14903
rect 19208 14844 19380 14872
rect 19208 14832 19214 14844
rect 17267 14776 17359 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 19444 14804 19472 14903
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 20180 14872 20208 14968
rect 21928 14949 21956 14980
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22520 14980 22845 15008
rect 22520 14968 22526 14980
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 23198 15008 23204 15020
rect 23155 14980 23204 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 23400 15017 23428 15048
rect 23474 15036 23480 15048
rect 23532 15076 23538 15088
rect 26988 15076 27016 15107
rect 30742 15104 30748 15156
rect 30800 15104 30806 15156
rect 34514 15104 34520 15156
rect 34572 15104 34578 15156
rect 35894 15104 35900 15156
rect 35952 15104 35958 15156
rect 37274 15104 37280 15156
rect 37332 15104 37338 15156
rect 43990 15104 43996 15156
rect 44048 15104 44054 15156
rect 44269 15147 44327 15153
rect 44269 15113 44281 15147
rect 44315 15144 44327 15147
rect 44542 15144 44548 15156
rect 44315 15116 44548 15144
rect 44315 15113 44327 15116
rect 44269 15107 44327 15113
rect 44542 15104 44548 15116
rect 44600 15104 44606 15156
rect 23532 15048 27016 15076
rect 29457 15079 29515 15085
rect 23532 15036 23538 15048
rect 29457 15045 29469 15079
rect 29503 15076 29515 15079
rect 30760 15076 30788 15104
rect 29503 15048 30696 15076
rect 30760 15048 31340 15076
rect 29503 15045 29515 15048
rect 29457 15039 29515 15045
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 25590 14968 25596 15020
rect 25648 14968 25654 15020
rect 25958 14968 25964 15020
rect 26016 14968 26022 15020
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 15008 26111 15011
rect 26099 14980 26372 15008
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14940 20407 14943
rect 21913 14943 21971 14949
rect 20395 14912 21864 14940
rect 20395 14909 20407 14912
rect 20349 14903 20407 14909
rect 20180 14844 20392 14872
rect 20364 14816 20392 14844
rect 20714 14832 20720 14884
rect 20772 14832 20778 14884
rect 21836 14872 21864 14912
rect 21913 14909 21925 14943
rect 21959 14909 21971 14943
rect 21913 14903 21971 14909
rect 25608 14872 25636 14968
rect 26344 14952 26372 14980
rect 26878 14968 26884 15020
rect 26936 15008 26942 15020
rect 27341 15011 27399 15017
rect 27341 15008 27353 15011
rect 26936 14980 27353 15008
rect 26936 14968 26942 14980
rect 27341 14977 27353 14980
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 29365 15011 29423 15017
rect 29365 15008 29377 15011
rect 29052 14980 29377 15008
rect 29052 14968 29058 14980
rect 29365 14977 29377 14980
rect 29411 14977 29423 15011
rect 29549 15011 29607 15017
rect 29549 15008 29561 15011
rect 29365 14971 29423 14977
rect 29472 14980 29561 15008
rect 25866 14900 25872 14952
rect 25924 14940 25930 14952
rect 26145 14943 26203 14949
rect 26145 14940 26157 14943
rect 25924 14912 26157 14940
rect 25924 14900 25930 14912
rect 26145 14909 26157 14912
rect 26191 14909 26203 14943
rect 26145 14903 26203 14909
rect 21836 14844 25636 14872
rect 26160 14872 26188 14903
rect 26326 14900 26332 14952
rect 26384 14900 26390 14952
rect 27062 14900 27068 14952
rect 27120 14940 27126 14952
rect 27433 14943 27491 14949
rect 27433 14940 27445 14943
rect 27120 14912 27445 14940
rect 27120 14900 27126 14912
rect 27433 14909 27445 14912
rect 27479 14909 27491 14943
rect 27433 14903 27491 14909
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 27540 14872 27568 14903
rect 26160 14844 27568 14872
rect 29472 14816 29500 14980
rect 29549 14977 29561 14980
rect 29595 15008 29607 15011
rect 29638 15008 29644 15020
rect 29595 14980 29644 15008
rect 29595 14977 29607 14980
rect 29549 14971 29607 14977
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 29840 14940 29868 14971
rect 30006 14968 30012 15020
rect 30064 15008 30070 15020
rect 30101 15011 30159 15017
rect 30101 15008 30113 15011
rect 30064 14980 30113 15008
rect 30064 14968 30070 14980
rect 30101 14977 30113 14980
rect 30147 14977 30159 15011
rect 30101 14971 30159 14977
rect 30282 14968 30288 15020
rect 30340 15008 30346 15020
rect 30377 15011 30435 15017
rect 30377 15008 30389 15011
rect 30340 14980 30389 15008
rect 30340 14968 30346 14980
rect 30377 14977 30389 14980
rect 30423 14977 30435 15011
rect 30377 14971 30435 14977
rect 30466 14968 30472 15020
rect 30524 14968 30530 15020
rect 30558 14968 30564 15020
rect 30616 14968 30622 15020
rect 30668 15017 30696 15048
rect 31312 15017 31340 15048
rect 34422 15036 34428 15088
rect 34480 15036 34486 15088
rect 34532 15076 34560 15104
rect 34532 15048 35204 15076
rect 30653 15011 30711 15017
rect 30653 14977 30665 15011
rect 30699 14977 30711 15011
rect 30653 14971 30711 14977
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 15008 30803 15011
rect 31113 15011 31171 15017
rect 31113 15008 31125 15011
rect 30791 14980 31125 15008
rect 30791 14977 30803 14980
rect 30745 14971 30803 14977
rect 31113 14977 31125 14980
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 31297 15011 31355 15017
rect 31297 14977 31309 15011
rect 31343 14977 31355 15011
rect 31297 14971 31355 14977
rect 31386 14968 31392 15020
rect 31444 14968 31450 15020
rect 31478 14968 31484 15020
rect 31536 15008 31542 15020
rect 35176 15017 35204 15048
rect 35342 15036 35348 15088
rect 35400 15036 35406 15088
rect 31573 15011 31631 15017
rect 31573 15008 31585 15011
rect 31536 14980 31585 15008
rect 31536 14968 31542 14980
rect 31573 14977 31585 14980
rect 31619 14977 31631 15011
rect 31573 14971 31631 14977
rect 31665 15011 31723 15017
rect 31665 14977 31677 15011
rect 31711 14977 31723 15011
rect 31665 14971 31723 14977
rect 35161 15011 35219 15017
rect 35161 14977 35173 15011
rect 35207 14977 35219 15011
rect 35161 14971 35219 14977
rect 30576 14940 30604 14968
rect 29840 14912 30604 14940
rect 31202 14900 31208 14952
rect 31260 14940 31266 14952
rect 31680 14940 31708 14971
rect 33413 14943 33471 14949
rect 33413 14940 33425 14943
rect 31260 14912 33425 14940
rect 31260 14900 31266 14912
rect 33413 14909 33425 14912
rect 33459 14909 33471 14943
rect 33413 14903 33471 14909
rect 34885 14943 34943 14949
rect 34885 14909 34897 14943
rect 34931 14940 34943 14943
rect 35360 14940 35388 15036
rect 35437 15011 35495 15017
rect 35437 14977 35449 15011
rect 35483 15008 35495 15011
rect 35912 15008 35940 15104
rect 35483 14980 35940 15008
rect 44008 15008 44036 15104
rect 44085 15011 44143 15017
rect 44085 15008 44097 15011
rect 44008 14980 44097 15008
rect 35483 14977 35495 14980
rect 35437 14971 35495 14977
rect 44085 14977 44097 14980
rect 44131 14977 44143 15011
rect 44085 14971 44143 14977
rect 34931 14912 35388 14940
rect 34931 14909 34943 14912
rect 34885 14903 34943 14909
rect 35710 14900 35716 14952
rect 35768 14900 35774 14952
rect 37826 14900 37832 14952
rect 37884 14900 37890 14952
rect 17644 14776 19472 14804
rect 17644 14764 17650 14776
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19668 14776 19993 14804
rect 19668 14764 19674 14776
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 19981 14767 20039 14773
rect 20346 14764 20352 14816
rect 20404 14764 20410 14816
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 20806 14804 20812 14816
rect 20496 14776 20812 14804
rect 20496 14764 20502 14776
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 22554 14764 22560 14816
rect 22612 14764 22618 14816
rect 23017 14807 23075 14813
rect 23017 14773 23029 14807
rect 23063 14804 23075 14807
rect 23750 14804 23756 14816
rect 23063 14776 23756 14804
rect 23063 14773 23075 14776
rect 23017 14767 23075 14773
rect 23750 14764 23756 14776
rect 23808 14804 23814 14816
rect 26142 14804 26148 14816
rect 23808 14776 26148 14804
rect 23808 14764 23814 14776
rect 26142 14764 26148 14776
rect 26200 14764 26206 14816
rect 29454 14764 29460 14816
rect 29512 14764 29518 14816
rect 30282 14764 30288 14816
rect 30340 14764 30346 14816
rect 30929 14807 30987 14813
rect 30929 14773 30941 14807
rect 30975 14804 30987 14807
rect 31478 14804 31484 14816
rect 30975 14776 31484 14804
rect 30975 14773 30987 14776
rect 30929 14767 30987 14773
rect 31478 14764 31484 14776
rect 31536 14764 31542 14816
rect 35253 14807 35311 14813
rect 35253 14773 35265 14807
rect 35299 14804 35311 14807
rect 35342 14804 35348 14816
rect 35299 14776 35348 14804
rect 35299 14773 35311 14776
rect 35253 14767 35311 14773
rect 35342 14764 35348 14776
rect 35400 14764 35406 14816
rect 36265 14807 36323 14813
rect 36265 14773 36277 14807
rect 36311 14804 36323 14807
rect 36354 14804 36360 14816
rect 36311 14776 36360 14804
rect 36311 14773 36323 14776
rect 36265 14767 36323 14773
rect 36354 14764 36360 14776
rect 36412 14764 36418 14816
rect 1104 14714 45172 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 45172 14714
rect 1104 14640 45172 14662
rect 7006 14560 7012 14612
rect 7064 14560 7070 14612
rect 8754 14560 8760 14612
rect 8812 14560 8818 14612
rect 10226 14560 10232 14612
rect 10284 14560 10290 14612
rect 11974 14560 11980 14612
rect 12032 14560 12038 14612
rect 12158 14560 12164 14612
rect 12216 14560 12222 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 13814 14600 13820 14612
rect 12584 14572 13820 14600
rect 12584 14560 12590 14572
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14148 14572 14841 14600
rect 14148 14560 14154 14572
rect 14829 14569 14841 14572
rect 14875 14569 14887 14603
rect 14829 14563 14887 14569
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 15344 14572 15485 14600
rect 15344 14560 15350 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 15473 14563 15531 14569
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 15896 14572 16865 14600
rect 15896 14560 15902 14572
rect 16853 14569 16865 14572
rect 16899 14600 16911 14603
rect 16899 14572 17359 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 7024 14473 7052 14560
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 8938 14464 8944 14476
rect 7055 14436 8944 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9217 14467 9275 14473
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 10244 14464 10272 14560
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13630 14532 13636 14544
rect 11848 14504 13636 14532
rect 11848 14492 11854 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 13832 14532 13860 14560
rect 14921 14535 14979 14541
rect 14921 14532 14933 14535
rect 13832 14504 14933 14532
rect 14921 14501 14933 14504
rect 14967 14501 14979 14535
rect 16758 14532 16764 14544
rect 14921 14495 14979 14501
rect 15304 14504 16764 14532
rect 9263 14436 10272 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 11422 14424 11428 14476
rect 11480 14424 11486 14476
rect 15304 14473 15332 14504
rect 16758 14492 16764 14504
rect 16816 14492 16822 14544
rect 17221 14535 17279 14541
rect 17221 14501 17233 14535
rect 17267 14501 17279 14535
rect 17331 14532 17359 14572
rect 17402 14560 17408 14612
rect 17460 14560 17466 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17512 14572 17877 14600
rect 17512 14532 17540 14572
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 17865 14563 17923 14569
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 19337 14603 19395 14609
rect 19337 14600 19349 14603
rect 18196 14572 19349 14600
rect 18196 14560 18202 14572
rect 19337 14569 19349 14572
rect 19383 14600 19395 14603
rect 20438 14600 20444 14612
rect 19383 14572 20444 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20625 14603 20683 14609
rect 20625 14569 20637 14603
rect 20671 14600 20683 14603
rect 20806 14600 20812 14612
rect 20671 14572 20812 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 22554 14560 22560 14612
rect 22612 14560 22618 14612
rect 23198 14560 23204 14612
rect 23256 14600 23262 14612
rect 23382 14600 23388 14612
rect 23256 14572 23388 14600
rect 23256 14560 23262 14572
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 25130 14560 25136 14612
rect 25188 14560 25194 14612
rect 26142 14560 26148 14612
rect 26200 14560 26206 14612
rect 26970 14560 26976 14612
rect 27028 14600 27034 14612
rect 27065 14603 27123 14609
rect 27065 14600 27077 14603
rect 27028 14572 27077 14600
rect 27028 14560 27034 14572
rect 27065 14569 27077 14572
rect 27111 14569 27123 14603
rect 27065 14563 27123 14569
rect 29362 14560 29368 14612
rect 29420 14600 29426 14612
rect 29549 14603 29607 14609
rect 29549 14600 29561 14603
rect 29420 14572 29561 14600
rect 29420 14560 29426 14572
rect 29549 14569 29561 14572
rect 29595 14569 29607 14603
rect 29549 14563 29607 14569
rect 30282 14560 30288 14612
rect 30340 14560 30346 14612
rect 31570 14560 31576 14612
rect 31628 14600 31634 14612
rect 31941 14603 31999 14609
rect 31941 14600 31953 14603
rect 31628 14572 31953 14600
rect 31628 14560 31634 14572
rect 31941 14569 31953 14572
rect 31987 14569 31999 14603
rect 31941 14563 31999 14569
rect 35710 14560 35716 14612
rect 35768 14600 35774 14612
rect 36449 14603 36507 14609
rect 36449 14600 36461 14603
rect 35768 14572 36461 14600
rect 35768 14560 35774 14572
rect 36449 14569 36461 14572
rect 36495 14569 36507 14603
rect 36449 14563 36507 14569
rect 17331 14504 17540 14532
rect 17773 14535 17831 14541
rect 17221 14495 17279 14501
rect 17773 14501 17785 14535
rect 17819 14532 17831 14535
rect 17819 14504 19104 14532
rect 17819 14501 17831 14504
rect 17773 14495 17831 14501
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 15289 14467 15347 14473
rect 14599 14436 15246 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 11900 14368 12081 14396
rect 7282 14288 7288 14340
rect 7340 14288 7346 14340
rect 9674 14328 9680 14340
rect 8510 14300 9680 14328
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 11900 14272 11928 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 14645 14399 14703 14405
rect 12299 14368 13216 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 13188 14272 13216 14368
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14660 14328 14688 14359
rect 15102 14356 15108 14408
rect 15160 14356 15166 14408
rect 15218 14396 15246 14436
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15620 14436 15761 14464
rect 15620 14424 15626 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 16482 14424 16488 14476
rect 16540 14424 16546 14476
rect 16666 14424 16672 14476
rect 16724 14424 16730 14476
rect 16942 14424 16948 14476
rect 17000 14424 17006 14476
rect 17236 14464 17264 14495
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17236 14436 17601 14464
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18138 14464 18144 14476
rect 18012 14436 18144 14464
rect 18012 14424 18018 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 19076 14464 19104 14504
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 19610 14532 19616 14544
rect 19300 14504 19616 14532
rect 19300 14492 19306 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 22572 14532 22600 14560
rect 22572 14504 27292 14532
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19076 14436 20177 14464
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 20349 14467 20407 14473
rect 20349 14433 20361 14467
rect 20395 14464 20407 14467
rect 20533 14467 20591 14473
rect 20533 14464 20545 14467
rect 20395 14436 20545 14464
rect 20395 14433 20407 14436
rect 20349 14427 20407 14433
rect 20533 14433 20545 14436
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14464 20683 14467
rect 21818 14464 21824 14476
rect 20671 14436 21824 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 15381 14399 15439 14405
rect 15218 14368 15332 14396
rect 15304 14328 15332 14368
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15427 14368 15853 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15746 14328 15752 14340
rect 14660 14300 15240 14328
rect 15304 14300 15752 14328
rect 10686 14220 10692 14272
rect 10744 14220 10750 14272
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 11606 14220 11612 14272
rect 11664 14220 11670 14272
rect 11882 14220 11888 14272
rect 11940 14220 11946 14272
rect 13170 14220 13176 14272
rect 13228 14220 13234 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 14185 14263 14243 14269
rect 14185 14260 14197 14263
rect 13412 14232 14197 14260
rect 13412 14220 13418 14232
rect 14185 14229 14197 14232
rect 14231 14229 14243 14263
rect 14185 14223 14243 14229
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 15102 14260 15108 14272
rect 14608 14232 15108 14260
rect 14608 14220 14614 14232
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 15212 14260 15240 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 15856 14328 15884 14359
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 16393 14399 16451 14405
rect 16393 14396 16405 14399
rect 16080 14368 16405 14396
rect 16080 14356 16086 14368
rect 16393 14365 16405 14368
rect 16439 14365 16451 14399
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 16393 14359 16451 14365
rect 16500 14368 16865 14396
rect 16500 14328 16528 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 15856 14300 16528 14328
rect 16669 14331 16727 14337
rect 16408 14272 16436 14300
rect 16669 14297 16681 14331
rect 16715 14297 16727 14331
rect 16960 14328 16988 14424
rect 17034 14356 17040 14408
rect 17092 14356 17098 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17494 14396 17500 14408
rect 17368 14368 17500 14396
rect 17368 14356 17374 14368
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17604 14368 17693 14396
rect 17604 14328 17632 14368
rect 17681 14365 17693 14368
rect 17727 14396 17739 14399
rect 17727 14368 17816 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 16960 14300 17632 14328
rect 17788 14328 17816 14368
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 17954 14328 17960 14340
rect 17788 14300 17960 14328
rect 16669 14291 16727 14297
rect 15378 14260 15384 14272
rect 15212 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14260 15442 14272
rect 15930 14260 15936 14272
rect 15436 14232 15936 14260
rect 15436 14220 15442 14232
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 16684 14260 16712 14291
rect 17954 14288 17960 14300
rect 18012 14288 18018 14340
rect 18616 14328 18644 14359
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19208 14368 19257 14396
rect 19208 14356 19214 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19245 14359 19303 14365
rect 19352 14368 19533 14396
rect 19352 14328 19380 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 19815 14405 19932 14406
rect 19815 14399 19947 14405
rect 19815 14378 19901 14399
rect 18156 14300 18644 14328
rect 18708 14300 19380 14328
rect 19815 14328 19843 14378
rect 19889 14365 19901 14378
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19978 14356 19984 14408
rect 20036 14356 20042 14408
rect 20070 14356 20076 14408
rect 20128 14356 20134 14408
rect 20438 14356 20444 14408
rect 20496 14356 20502 14408
rect 20530 14328 20536 14340
rect 19815 14300 20536 14328
rect 18156 14260 18184 14300
rect 18708 14269 18736 14300
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 16684 14232 18184 14260
rect 18233 14263 18291 14269
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18279 14232 18705 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 18966 14220 18972 14272
rect 19024 14260 19030 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 19024 14232 19073 14260
rect 19024 14220 19030 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 19061 14223 19119 14229
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19484 14232 19625 14260
rect 19484 14220 19490 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 20640 14260 20668 14427
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 25777 14467 25835 14473
rect 25777 14433 25789 14467
rect 25823 14464 25835 14467
rect 25866 14464 25872 14476
rect 25823 14436 25872 14464
rect 25823 14433 25835 14436
rect 25777 14427 25835 14433
rect 25866 14424 25872 14436
rect 25924 14464 25930 14476
rect 26697 14467 26755 14473
rect 26697 14464 26709 14467
rect 25924 14436 26709 14464
rect 25924 14424 25930 14436
rect 26697 14433 26709 14436
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 26786 14424 26792 14476
rect 26844 14464 26850 14476
rect 26844 14436 27016 14464
rect 26844 14424 26850 14436
rect 26988 14405 27016 14436
rect 26973 14399 27031 14405
rect 26973 14365 26985 14399
rect 27019 14365 27031 14399
rect 27157 14399 27215 14405
rect 27157 14396 27169 14399
rect 26973 14359 27031 14365
rect 27080 14368 27169 14396
rect 20809 14331 20867 14337
rect 20809 14297 20821 14331
rect 20855 14328 20867 14331
rect 21726 14328 21732 14340
rect 20855 14300 21732 14328
rect 20855 14297 20867 14300
rect 20809 14291 20867 14297
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 25501 14331 25559 14337
rect 25501 14297 25513 14331
rect 25547 14328 25559 14331
rect 25547 14300 26648 14328
rect 25547 14297 25559 14300
rect 25501 14291 25559 14297
rect 20312 14232 20668 14260
rect 20312 14220 20318 14232
rect 25590 14220 25596 14272
rect 25648 14220 25654 14272
rect 26510 14220 26516 14272
rect 26568 14220 26574 14272
rect 26620 14269 26648 14300
rect 27080 14272 27108 14368
rect 27157 14365 27169 14368
rect 27203 14365 27215 14399
rect 27157 14359 27215 14365
rect 27264 14328 27292 14504
rect 30006 14424 30012 14476
rect 30064 14464 30070 14476
rect 30101 14467 30159 14473
rect 30101 14464 30113 14467
rect 30064 14436 30113 14464
rect 30064 14424 30070 14436
rect 30101 14433 30113 14436
rect 30147 14433 30159 14467
rect 30101 14427 30159 14433
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14396 30251 14399
rect 30300 14396 30328 14560
rect 31754 14424 31760 14476
rect 31812 14464 31818 14476
rect 31812 14436 32260 14464
rect 31812 14424 31818 14436
rect 30239 14368 30328 14396
rect 30239 14365 30251 14368
rect 30193 14359 30251 14365
rect 30374 14356 30380 14408
rect 30432 14396 30438 14408
rect 30837 14399 30895 14405
rect 30837 14396 30849 14399
rect 30432 14368 30849 14396
rect 30432 14356 30438 14368
rect 30837 14365 30849 14368
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 31726 14368 32076 14396
rect 31726 14328 31754 14368
rect 27264 14300 31754 14328
rect 31846 14288 31852 14340
rect 31904 14328 31910 14340
rect 31941 14331 31999 14337
rect 31941 14328 31953 14331
rect 31904 14300 31953 14328
rect 31904 14288 31910 14300
rect 31941 14297 31953 14300
rect 31987 14297 31999 14331
rect 32048 14328 32076 14368
rect 32122 14356 32128 14408
rect 32180 14356 32186 14408
rect 32232 14405 32260 14436
rect 34514 14424 34520 14476
rect 34572 14464 34578 14476
rect 34701 14467 34759 14473
rect 34701 14464 34713 14467
rect 34572 14436 34713 14464
rect 34572 14424 34578 14436
rect 34701 14433 34713 14436
rect 34747 14433 34759 14467
rect 34701 14427 34759 14433
rect 34977 14467 35035 14473
rect 34977 14433 34989 14467
rect 35023 14464 35035 14467
rect 35342 14464 35348 14476
rect 35023 14436 35348 14464
rect 35023 14433 35035 14436
rect 34977 14427 35035 14433
rect 35342 14424 35348 14436
rect 35400 14424 35406 14476
rect 32217 14399 32275 14405
rect 32217 14365 32229 14399
rect 32263 14365 32275 14399
rect 32217 14359 32275 14365
rect 35986 14356 35992 14408
rect 36044 14396 36050 14408
rect 36814 14396 36820 14408
rect 36044 14368 36820 14396
rect 36044 14356 36050 14368
rect 36814 14356 36820 14368
rect 36872 14356 36878 14408
rect 38654 14356 38660 14408
rect 38712 14356 38718 14408
rect 33134 14328 33140 14340
rect 32048 14300 33140 14328
rect 31941 14291 31999 14297
rect 33134 14288 33140 14300
rect 33192 14288 33198 14340
rect 26605 14263 26663 14269
rect 26605 14229 26617 14263
rect 26651 14260 26663 14263
rect 26694 14260 26700 14272
rect 26651 14232 26700 14260
rect 26651 14229 26663 14232
rect 26605 14223 26663 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 27062 14220 27068 14272
rect 27120 14220 27126 14272
rect 32401 14263 32459 14269
rect 32401 14229 32413 14263
rect 32447 14260 32459 14263
rect 38672 14260 38700 14356
rect 32447 14232 38700 14260
rect 32447 14229 32459 14232
rect 32401 14223 32459 14229
rect 1104 14170 45172 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 45172 14170
rect 1104 14096 45172 14118
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 7377 14059 7435 14065
rect 7377 14056 7389 14059
rect 7340 14028 7389 14056
rect 7340 14016 7346 14028
rect 7377 14025 7389 14028
rect 7423 14025 7435 14059
rect 7377 14019 7435 14025
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 11572 14028 12357 14056
rect 11572 14016 11578 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 14090 14056 14096 14068
rect 12345 14019 12403 14025
rect 12636 14028 14096 14056
rect 7190 13880 7196 13932
rect 7248 13880 7254 13932
rect 11974 13880 11980 13932
rect 12032 13880 12038 13932
rect 12526 13880 12532 13932
rect 12584 13880 12590 13932
rect 12636 13929 12664 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14332 14028 14473 14056
rect 14332 14016 14338 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 14734 14016 14740 14068
rect 14792 14016 14798 14068
rect 15286 14016 15292 14068
rect 15344 14016 15350 14068
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 17770 14056 17776 14068
rect 17727 14028 17776 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 12851 13991 12909 13997
rect 12851 13957 12863 13991
rect 12897 13988 12909 13991
rect 13354 13988 13360 14000
rect 12897 13960 13360 13988
rect 12897 13957 12909 13960
rect 12851 13951 12909 13957
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 14752 13988 14780 14016
rect 13872 13960 14780 13988
rect 15304 13988 15332 14016
rect 16224 13988 16252 14019
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 20438 14056 20444 14068
rect 19107 14028 20444 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 24302 14016 24308 14068
rect 24360 14016 24366 14068
rect 24581 14059 24639 14065
rect 24581 14025 24593 14059
rect 24627 14056 24639 14059
rect 24854 14056 24860 14068
rect 24627 14028 24860 14056
rect 24627 14025 24639 14028
rect 24581 14019 24639 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 25038 14016 25044 14068
rect 25096 14016 25102 14068
rect 25133 14059 25191 14065
rect 25133 14025 25145 14059
rect 25179 14056 25191 14059
rect 26142 14056 26148 14068
rect 25179 14028 26148 14056
rect 25179 14025 25191 14028
rect 25133 14019 25191 14025
rect 26142 14016 26148 14028
rect 26200 14056 26206 14068
rect 26602 14056 26608 14068
rect 26200 14028 26608 14056
rect 26200 14016 26206 14028
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 26694 14016 26700 14068
rect 26752 14056 26758 14068
rect 27246 14056 27252 14068
rect 26752 14028 27252 14056
rect 26752 14016 26758 14028
rect 27246 14016 27252 14028
rect 27304 14016 27310 14068
rect 28902 14016 28908 14068
rect 28960 14056 28966 14068
rect 31941 14059 31999 14065
rect 28960 14028 31754 14056
rect 28960 14016 28966 14028
rect 15304 13960 16068 13988
rect 16224 13960 18184 13988
rect 13872 13948 13878 13960
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 11992 13852 12020 13880
rect 12728 13852 12756 13883
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13136 13892 14105 13920
rect 13136 13880 13142 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14274 13880 14280 13932
rect 14332 13880 14338 13932
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14642 13880 14648 13932
rect 14700 13880 14706 13932
rect 14826 13880 14832 13932
rect 14884 13880 14890 13932
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 11992 13824 12756 13852
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13852 13047 13855
rect 13814 13852 13820 13864
rect 13035 13824 13820 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13998 13812 14004 13864
rect 14056 13812 14062 13864
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14568 13852 14596 13880
rect 14240 13824 14596 13852
rect 14660 13852 14688 13880
rect 15194 13852 15200 13864
rect 14660 13824 15200 13852
rect 14240 13812 14246 13824
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 15580 13852 15608 13883
rect 15654 13880 15660 13932
rect 15712 13880 15718 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15804 13892 15853 13920
rect 15804 13880 15810 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 15930 13880 15936 13932
rect 15988 13880 15994 13932
rect 16040 13929 16068 13960
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13889 16083 13923
rect 16025 13883 16083 13889
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16448 13892 17417 13920
rect 16448 13880 16454 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 18156 13920 18184 13960
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 18693 13991 18751 13997
rect 18693 13988 18705 13991
rect 18564 13960 18705 13988
rect 18564 13948 18570 13960
rect 18693 13957 18705 13960
rect 18739 13957 18751 13991
rect 18693 13951 18751 13957
rect 18782 13948 18788 14000
rect 18840 13988 18846 14000
rect 18893 13991 18951 13997
rect 18893 13988 18905 13991
rect 18840 13960 18905 13988
rect 18840 13948 18846 13960
rect 18893 13957 18905 13960
rect 18939 13957 18951 13991
rect 18893 13951 18951 13957
rect 20070 13948 20076 14000
rect 20128 13948 20134 14000
rect 24504 13960 28948 13988
rect 20088 13920 20116 13948
rect 18156 13892 20116 13920
rect 17405 13883 17463 13889
rect 20714 13880 20720 13932
rect 20772 13880 20778 13932
rect 24504 13929 24532 13960
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13889 24363 13923
rect 24305 13883 24363 13889
rect 24489 13923 24547 13929
rect 24489 13889 24501 13923
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 16574 13852 16580 13864
rect 15580 13824 16580 13852
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 16666 13812 16672 13864
rect 16724 13812 16730 13864
rect 17310 13812 17316 13864
rect 17368 13812 17374 13864
rect 17494 13812 17500 13864
rect 17552 13852 17558 13864
rect 17681 13855 17739 13861
rect 17681 13852 17693 13855
rect 17552 13824 17693 13852
rect 17552 13812 17558 13824
rect 17681 13821 17693 13824
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 20732 13852 20760 13880
rect 19208 13824 20760 13852
rect 19208 13812 19214 13824
rect 11256 13756 22094 13784
rect 11256 13728 11284 13756
rect 11238 13676 11244 13728
rect 11296 13676 11302 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 13998 13716 14004 13728
rect 11388 13688 14004 13716
rect 11388 13676 11394 13688
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 14734 13676 14740 13728
rect 14792 13716 14798 13728
rect 16298 13716 16304 13728
rect 14792 13688 16304 13716
rect 14792 13676 14798 13688
rect 16298 13676 16304 13688
rect 16356 13716 16362 13728
rect 17034 13716 17040 13728
rect 16356 13688 17040 13716
rect 16356 13676 16362 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 17276 13688 17509 13716
rect 17276 13676 17282 13688
rect 17497 13685 17509 13688
rect 17543 13716 17555 13719
rect 17586 13716 17592 13728
rect 17543 13688 17592 13716
rect 17543 13685 17555 13688
rect 17497 13679 17555 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18877 13719 18935 13725
rect 18877 13685 18889 13719
rect 18923 13716 18935 13719
rect 18966 13716 18972 13728
rect 18923 13688 18972 13716
rect 18923 13685 18935 13688
rect 18877 13679 18935 13685
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 22066 13716 22094 13756
rect 24118 13744 24124 13796
rect 24176 13784 24182 13796
rect 24320 13784 24348 13883
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 24728 13892 24869 13920
rect 24728 13880 24734 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13920 25283 13923
rect 25590 13920 25596 13932
rect 25271 13892 25596 13920
rect 25271 13889 25283 13892
rect 25225 13883 25283 13889
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 28920 13929 28948 13960
rect 30834 13948 30840 14000
rect 30892 13988 30898 14000
rect 31386 13988 31392 14000
rect 30892 13960 31392 13988
rect 30892 13948 30898 13960
rect 31386 13948 31392 13960
rect 31444 13988 31450 14000
rect 31481 13991 31539 13997
rect 31481 13988 31493 13991
rect 31444 13960 31493 13988
rect 31444 13948 31450 13960
rect 31481 13957 31493 13960
rect 31527 13957 31539 13991
rect 31726 13988 31754 14028
rect 31941 14025 31953 14059
rect 31987 14056 31999 14059
rect 32122 14056 32128 14068
rect 31987 14028 32128 14056
rect 31987 14025 31999 14028
rect 31941 14019 31999 14025
rect 32122 14016 32128 14028
rect 32180 14016 32186 14068
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37332 14028 39896 14056
rect 37332 14016 37338 14028
rect 31726 13960 32904 13988
rect 31481 13951 31539 13957
rect 28905 13923 28963 13929
rect 28905 13889 28917 13923
rect 28951 13920 28963 13923
rect 31018 13920 31024 13932
rect 28951 13892 31024 13920
rect 28951 13889 28963 13892
rect 28905 13883 28963 13889
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 31757 13923 31815 13929
rect 31757 13920 31769 13923
rect 31128 13892 31769 13920
rect 24578 13812 24584 13864
rect 24636 13852 24642 13864
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 24636 13824 24777 13852
rect 24636 13812 24642 13824
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 28721 13855 28779 13861
rect 28721 13852 28733 13855
rect 24765 13815 24823 13821
rect 24872 13824 28733 13852
rect 24872 13784 24900 13824
rect 28721 13821 28733 13824
rect 28767 13852 28779 13855
rect 28767 13824 28994 13852
rect 28767 13821 28779 13824
rect 28721 13815 28779 13821
rect 24176 13756 24900 13784
rect 24176 13744 24182 13756
rect 24946 13744 24952 13796
rect 25004 13784 25010 13796
rect 26786 13784 26792 13796
rect 25004 13756 26792 13784
rect 25004 13744 25010 13756
rect 26786 13744 26792 13756
rect 26844 13744 26850 13796
rect 28966 13784 28994 13824
rect 29086 13812 29092 13864
rect 29144 13812 29150 13864
rect 31128 13784 31156 13892
rect 31757 13889 31769 13892
rect 31803 13920 31815 13923
rect 31938 13920 31944 13932
rect 31803 13892 31944 13920
rect 31803 13889 31815 13892
rect 31757 13883 31815 13889
rect 31938 13880 31944 13892
rect 31996 13880 32002 13932
rect 32876 13929 32904 13960
rect 33134 13948 33140 14000
rect 33192 13948 33198 14000
rect 35986 13948 35992 14000
rect 36044 13948 36050 14000
rect 36354 13948 36360 14000
rect 36412 13988 36418 14000
rect 36449 13991 36507 13997
rect 36449 13988 36461 13991
rect 36412 13960 36461 13988
rect 36412 13948 36418 13960
rect 36449 13957 36461 13960
rect 36495 13957 36507 13991
rect 36449 13951 36507 13957
rect 36814 13948 36820 14000
rect 36872 13988 36878 14000
rect 39868 13997 39896 14028
rect 39853 13991 39911 13997
rect 36872 13960 38594 13988
rect 36872 13948 36878 13960
rect 39853 13957 39865 13991
rect 39899 13957 39911 13991
rect 39853 13951 39911 13957
rect 32861 13923 32919 13929
rect 32861 13889 32873 13923
rect 32907 13889 32919 13923
rect 34422 13920 34428 13932
rect 34270 13892 34428 13920
rect 32861 13883 32919 13889
rect 34422 13880 34428 13892
rect 34480 13920 34486 13932
rect 36725 13923 36783 13929
rect 34480 13892 35112 13920
rect 34480 13880 34486 13892
rect 31665 13855 31723 13861
rect 31665 13821 31677 13855
rect 31711 13852 31723 13855
rect 34977 13855 35035 13861
rect 34977 13852 34989 13855
rect 31711 13824 34989 13852
rect 31711 13821 31723 13824
rect 31665 13815 31723 13821
rect 34977 13821 34989 13824
rect 35023 13821 35035 13855
rect 35084 13852 35112 13892
rect 36725 13889 36737 13923
rect 36771 13920 36783 13923
rect 37734 13920 37740 13932
rect 36771 13892 37740 13920
rect 36771 13889 36783 13892
rect 36725 13883 36783 13889
rect 37734 13880 37740 13892
rect 37792 13920 37798 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 37792 13892 37841 13920
rect 37792 13880 37798 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 35986 13852 35992 13864
rect 35084 13824 35992 13852
rect 34977 13815 35035 13821
rect 35986 13812 35992 13824
rect 36044 13812 36050 13864
rect 28966 13756 31156 13784
rect 39500 13756 40632 13784
rect 30926 13716 30932 13728
rect 22066 13688 30932 13716
rect 30926 13676 30932 13688
rect 30984 13676 30990 13728
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 31481 13719 31539 13725
rect 31481 13716 31493 13719
rect 31168 13688 31493 13716
rect 31168 13676 31174 13688
rect 31481 13685 31493 13688
rect 31527 13685 31539 13719
rect 31481 13679 31539 13685
rect 34606 13676 34612 13728
rect 34664 13676 34670 13728
rect 38092 13719 38150 13725
rect 38092 13685 38104 13719
rect 38138 13716 38150 13719
rect 39500 13716 39528 13756
rect 38138 13688 39528 13716
rect 38138 13685 38150 13688
rect 38092 13679 38150 13685
rect 39574 13676 39580 13728
rect 39632 13676 39638 13728
rect 40604 13716 40632 13756
rect 40678 13744 40684 13796
rect 40736 13784 40742 13796
rect 41141 13787 41199 13793
rect 41141 13784 41153 13787
rect 40736 13756 41153 13784
rect 40736 13744 40742 13756
rect 41141 13753 41153 13756
rect 41187 13784 41199 13787
rect 41230 13784 41236 13796
rect 41187 13756 41236 13784
rect 41187 13753 41199 13756
rect 41141 13747 41199 13753
rect 41230 13744 41236 13756
rect 41288 13744 41294 13796
rect 43622 13784 43628 13796
rect 41386 13756 43628 13784
rect 41386 13716 41414 13756
rect 43622 13744 43628 13756
rect 43680 13744 43686 13796
rect 40604 13688 41414 13716
rect 1104 13626 45172 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 45172 13626
rect 1104 13552 45172 13574
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7190 13512 7196 13524
rect 7147 13484 7196 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 11330 13512 11336 13524
rect 8864 13484 11336 13512
rect 6914 13404 6920 13456
rect 6972 13404 6978 13456
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 7006 13376 7012 13388
rect 6687 13348 7012 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 7006 13336 7012 13348
rect 7064 13376 7070 13388
rect 8864 13376 8892 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 12342 13512 12348 13524
rect 11931 13484 12348 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12584 13484 12817 13512
rect 12584 13472 12590 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 24946 13512 24952 13524
rect 14056 13484 24952 13512
rect 14056 13472 14062 13484
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 26602 13472 26608 13524
rect 26660 13472 26666 13524
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 34146 13512 34152 13524
rect 26844 13484 34152 13512
rect 26844 13472 26850 13484
rect 34146 13472 34152 13484
rect 34204 13472 34210 13524
rect 36909 13515 36967 13521
rect 36909 13481 36921 13515
rect 36955 13512 36967 13515
rect 37826 13512 37832 13524
rect 36955 13484 37832 13512
rect 36955 13481 36967 13484
rect 36909 13475 36967 13481
rect 37826 13472 37832 13484
rect 37884 13472 37890 13524
rect 10689 13447 10747 13453
rect 10689 13413 10701 13447
rect 10735 13444 10747 13447
rect 16666 13444 16672 13456
rect 10735 13416 16672 13444
rect 10735 13413 10747 13416
rect 10689 13407 10747 13413
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 22005 13447 22063 13453
rect 22005 13413 22017 13447
rect 22051 13444 22063 13447
rect 22278 13444 22284 13456
rect 22051 13416 22284 13444
rect 22051 13413 22063 13416
rect 22005 13407 22063 13413
rect 22278 13404 22284 13416
rect 22336 13404 22342 13456
rect 24118 13404 24124 13456
rect 24176 13404 24182 13456
rect 25317 13447 25375 13453
rect 25317 13413 25329 13447
rect 25363 13444 25375 13447
rect 25590 13444 25596 13456
rect 25363 13416 25596 13444
rect 25363 13413 25375 13416
rect 25317 13407 25375 13413
rect 25590 13404 25596 13416
rect 25648 13404 25654 13456
rect 26050 13404 26056 13456
rect 26108 13404 26114 13456
rect 26421 13447 26479 13453
rect 26421 13413 26433 13447
rect 26467 13413 26479 13447
rect 26421 13407 26479 13413
rect 26712 13416 27016 13444
rect 7064 13348 8892 13376
rect 7064 13336 7070 13348
rect 8938 13336 8944 13388
rect 8996 13336 9002 13388
rect 11790 13376 11796 13388
rect 11532 13348 11796 13376
rect 11532 13317 11560 13348
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12912 13376 13032 13384
rect 14734 13376 14740 13388
rect 12912 13374 14740 13376
rect 12897 13368 14740 13374
rect 12897 13334 12909 13368
rect 12943 13356 14740 13368
rect 12943 13334 12955 13356
rect 13004 13348 14740 13356
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 19334 13376 19340 13388
rect 15160 13348 19340 13376
rect 15160 13336 15166 13348
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 21910 13336 21916 13388
rect 21968 13336 21974 13388
rect 22646 13336 22652 13388
rect 22704 13336 22710 13388
rect 23014 13336 23020 13388
rect 23072 13376 23078 13388
rect 24854 13376 24860 13388
rect 23072 13348 24860 13376
rect 23072 13336 23078 13348
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 26145 13379 26203 13385
rect 25087 13348 26096 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 12897 13328 12955 13334
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 11348 13280 11437 13308
rect 9214 13200 9220 13252
rect 9272 13200 9278 13252
rect 9950 13200 9956 13252
rect 10008 13200 10014 13252
rect 11348 13184 11376 13280
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 11716 13240 11744 13271
rect 11440 13212 11744 13240
rect 12636 13240 12664 13271
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13078 13308 13084 13320
rect 13035 13280 13084 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 12894 13240 12900 13252
rect 12636 13212 12900 13240
rect 11440 13184 11468 13212
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 11330 13132 11336 13184
rect 11388 13132 11394 13184
rect 11422 13132 11428 13184
rect 11480 13132 11486 13184
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 13004 13172 13032 13271
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 15470 13308 15476 13320
rect 13688 13280 15476 13308
rect 13688 13268 13694 13280
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16632 13280 17908 13308
rect 16632 13268 16638 13280
rect 13722 13200 13728 13252
rect 13780 13240 13786 13252
rect 16666 13240 16672 13252
rect 13780 13212 16672 13240
rect 13780 13200 13786 13212
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 17880 13240 17908 13280
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 19150 13308 19156 13320
rect 18012 13280 19156 13308
rect 18012 13268 18018 13280
rect 19150 13268 19156 13280
rect 19208 13308 19214 13320
rect 20806 13308 20812 13320
rect 19208 13280 20812 13308
rect 19208 13268 19214 13280
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 22094 13268 22100 13320
rect 22152 13268 22158 13320
rect 22188 13289 22246 13295
rect 22188 13255 22200 13289
rect 22234 13255 22246 13289
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 24394 13268 24400 13320
rect 24452 13308 24458 13320
rect 24673 13311 24731 13317
rect 24673 13308 24685 13311
rect 24452 13280 24685 13308
rect 24452 13268 24458 13280
rect 24673 13277 24685 13280
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 24946 13268 24952 13320
rect 25004 13268 25010 13320
rect 25866 13268 25872 13320
rect 25924 13268 25930 13320
rect 25961 13311 26019 13317
rect 25961 13277 25973 13311
rect 26007 13277 26019 13311
rect 26068 13308 26096 13348
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 26436 13376 26464 13407
rect 26712 13385 26740 13416
rect 26191 13348 26464 13376
rect 26697 13379 26755 13385
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 26697 13345 26709 13379
rect 26743 13345 26755 13379
rect 26881 13379 26939 13385
rect 26881 13376 26893 13379
rect 26697 13339 26755 13345
rect 26804 13348 26893 13376
rect 26804 13320 26832 13348
rect 26881 13345 26893 13348
rect 26927 13345 26939 13379
rect 26881 13339 26939 13345
rect 26988 13320 27016 13416
rect 27246 13404 27252 13456
rect 27304 13404 27310 13456
rect 31018 13404 31024 13456
rect 31076 13404 31082 13456
rect 31202 13404 31208 13456
rect 31260 13444 31266 13456
rect 31570 13444 31576 13456
rect 31260 13416 31576 13444
rect 31260 13404 31266 13416
rect 31570 13404 31576 13416
rect 31628 13404 31634 13456
rect 31665 13447 31723 13453
rect 31665 13413 31677 13447
rect 31711 13444 31723 13447
rect 31846 13444 31852 13456
rect 31711 13416 31852 13444
rect 31711 13413 31723 13416
rect 31665 13407 31723 13413
rect 31846 13404 31852 13416
rect 31904 13404 31910 13456
rect 32217 13447 32275 13453
rect 32217 13444 32229 13447
rect 31956 13416 32229 13444
rect 27065 13379 27123 13385
rect 27065 13345 27077 13379
rect 27111 13376 27123 13379
rect 27706 13376 27712 13388
rect 27111 13348 27712 13376
rect 27111 13345 27123 13348
rect 27065 13339 27123 13345
rect 27706 13336 27712 13348
rect 27764 13336 27770 13388
rect 27801 13379 27859 13385
rect 27801 13345 27813 13379
rect 27847 13376 27859 13379
rect 28629 13379 28687 13385
rect 28629 13376 28641 13379
rect 27847 13348 28641 13376
rect 27847 13345 27859 13348
rect 27801 13339 27859 13345
rect 26602 13308 26608 13320
rect 26068 13280 26608 13308
rect 25961 13271 26019 13277
rect 22188 13252 22246 13255
rect 18230 13240 18236 13252
rect 17880 13212 18236 13240
rect 18230 13200 18236 13212
rect 18288 13240 18294 13252
rect 18288 13212 19334 13240
rect 18288 13200 18294 13212
rect 19306 13184 19334 13212
rect 20254 13200 20260 13252
rect 20312 13240 20318 13252
rect 22186 13240 22192 13252
rect 20312 13212 22192 13240
rect 20312 13200 20318 13212
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 23874 13212 24532 13240
rect 12676 13144 13032 13172
rect 12676 13132 12682 13144
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 15930 13172 15936 13184
rect 13136 13144 15936 13172
rect 13136 13132 13142 13144
rect 15930 13132 15936 13144
rect 15988 13172 15994 13184
rect 16758 13172 16764 13184
rect 15988 13144 16764 13172
rect 15988 13132 15994 13144
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 19306 13144 19340 13184
rect 19334 13132 19340 13144
rect 19392 13172 19398 13184
rect 20622 13172 20628 13184
rect 19392 13144 20628 13172
rect 19392 13132 19398 13144
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 24504 13181 24532 13212
rect 25774 13200 25780 13252
rect 25832 13240 25838 13252
rect 25976 13240 26004 13271
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 26786 13268 26792 13320
rect 26844 13268 26850 13320
rect 26970 13268 26976 13320
rect 27028 13308 27034 13320
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 27028 13280 27169 13308
rect 27028 13268 27034 13280
rect 27157 13277 27169 13280
rect 27203 13308 27215 13311
rect 27816 13308 27844 13339
rect 27203 13280 27844 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 26881 13243 26939 13249
rect 26881 13240 26893 13243
rect 25832 13212 26893 13240
rect 25832 13200 25838 13212
rect 26881 13209 26893 13212
rect 26927 13209 26939 13243
rect 28460 13240 28488 13348
rect 28629 13345 28641 13348
rect 28675 13345 28687 13379
rect 31036 13376 31064 13404
rect 31956 13376 31984 13416
rect 32217 13413 32229 13416
rect 32263 13444 32275 13447
rect 42337 13447 42395 13453
rect 42337 13444 42349 13447
rect 32263 13416 37688 13444
rect 32263 13413 32275 13416
rect 32217 13407 32275 13413
rect 37660 13385 37688 13416
rect 41064 13416 42349 13444
rect 31036 13348 31984 13376
rect 32401 13379 32459 13385
rect 28629 13339 28687 13345
rect 32401 13345 32413 13379
rect 32447 13345 32459 13379
rect 32401 13339 32459 13345
rect 36265 13379 36323 13385
rect 36265 13345 36277 13379
rect 36311 13376 36323 13379
rect 36633 13379 36691 13385
rect 36633 13376 36645 13379
rect 36311 13348 36645 13376
rect 36311 13345 36323 13348
rect 36265 13339 36323 13345
rect 36633 13345 36645 13348
rect 36679 13345 36691 13379
rect 36633 13339 36691 13345
rect 37645 13379 37703 13385
rect 37645 13345 37657 13379
rect 37691 13376 37703 13379
rect 38746 13376 38752 13388
rect 37691 13348 38752 13376
rect 37691 13345 37703 13348
rect 37645 13339 37703 13345
rect 28537 13311 28595 13317
rect 28537 13277 28549 13311
rect 28583 13308 28595 13311
rect 29270 13308 29276 13320
rect 28583 13280 29276 13308
rect 28583 13277 28595 13280
rect 28537 13271 28595 13277
rect 29270 13268 29276 13280
rect 29328 13268 29334 13320
rect 30926 13268 30932 13320
rect 30984 13308 30990 13320
rect 31481 13311 31539 13317
rect 31481 13308 31493 13311
rect 30984 13280 31493 13308
rect 30984 13268 30990 13280
rect 31481 13277 31493 13280
rect 31527 13308 31539 13311
rect 31662 13308 31668 13320
rect 31527 13280 31668 13308
rect 31527 13277 31539 13280
rect 31481 13271 31539 13277
rect 31662 13268 31668 13280
rect 31720 13268 31726 13320
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 32122 13308 32128 13320
rect 31812 13280 32128 13308
rect 31812 13268 31818 13280
rect 32122 13268 32128 13280
rect 32180 13308 32186 13320
rect 32416 13308 32444 13339
rect 38746 13336 38752 13348
rect 38804 13336 38810 13388
rect 39574 13336 39580 13388
rect 39632 13376 39638 13388
rect 39853 13379 39911 13385
rect 39853 13376 39865 13379
rect 39632 13348 39865 13376
rect 39632 13336 39638 13348
rect 39853 13345 39865 13348
rect 39899 13345 39911 13379
rect 39853 13339 39911 13345
rect 32674 13308 32680 13320
rect 32180 13280 32680 13308
rect 32180 13268 32186 13280
rect 32674 13268 32680 13280
rect 32732 13268 32738 13320
rect 34146 13268 34152 13320
rect 34204 13268 34210 13320
rect 34606 13268 34612 13320
rect 34664 13308 34670 13320
rect 35618 13308 35624 13320
rect 34664 13280 35624 13308
rect 34664 13268 34670 13280
rect 35618 13268 35624 13280
rect 35676 13268 35682 13320
rect 36078 13268 36084 13320
rect 36136 13308 36142 13320
rect 36541 13311 36599 13317
rect 36541 13308 36553 13311
rect 36136 13280 36553 13308
rect 36136 13268 36142 13280
rect 36541 13277 36553 13280
rect 36587 13277 36599 13311
rect 36541 13271 36599 13277
rect 29089 13243 29147 13249
rect 29089 13240 29101 13243
rect 26881 13203 26939 13209
rect 26988 13212 28120 13240
rect 28460 13212 29101 13240
rect 24489 13175 24547 13181
rect 24489 13141 24501 13175
rect 24535 13172 24547 13175
rect 26234 13172 26240 13184
rect 24535 13144 26240 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 26510 13132 26516 13184
rect 26568 13172 26574 13184
rect 26988 13172 27016 13212
rect 26568 13144 27016 13172
rect 26568 13132 26574 13144
rect 27614 13132 27620 13184
rect 27672 13132 27678 13184
rect 28092 13181 28120 13212
rect 29089 13209 29101 13212
rect 29135 13209 29147 13243
rect 29089 13203 29147 13209
rect 29840 13212 31754 13240
rect 28077 13175 28135 13181
rect 28077 13141 28089 13175
rect 28123 13141 28135 13175
rect 28077 13135 28135 13141
rect 28442 13132 28448 13184
rect 28500 13132 28506 13184
rect 28902 13132 28908 13184
rect 28960 13132 28966 13184
rect 28994 13132 29000 13184
rect 29052 13172 29058 13184
rect 29840 13172 29868 13212
rect 29052 13144 29868 13172
rect 29052 13132 29058 13144
rect 29914 13132 29920 13184
rect 29972 13172 29978 13184
rect 31297 13175 31355 13181
rect 31297 13172 31309 13175
rect 29972 13144 31309 13172
rect 29972 13132 29978 13144
rect 31297 13141 31309 13144
rect 31343 13141 31355 13175
rect 31726 13172 31754 13212
rect 31938 13200 31944 13252
rect 31996 13200 32002 13252
rect 34164 13240 34192 13268
rect 34793 13243 34851 13249
rect 34793 13240 34805 13243
rect 34164 13212 34805 13240
rect 34793 13209 34805 13212
rect 34839 13240 34851 13243
rect 36556 13240 36584 13271
rect 36722 13268 36728 13320
rect 36780 13268 36786 13320
rect 37001 13311 37059 13317
rect 37001 13308 37013 13311
rect 36832 13280 37013 13308
rect 36832 13240 36860 13280
rect 37001 13277 37013 13280
rect 37047 13277 37059 13311
rect 37001 13271 37059 13277
rect 37090 13268 37096 13320
rect 37148 13308 37154 13320
rect 37277 13311 37335 13317
rect 37277 13308 37289 13311
rect 37148 13280 37289 13308
rect 37148 13268 37154 13280
rect 37277 13277 37289 13280
rect 37323 13277 37335 13311
rect 37277 13271 37335 13277
rect 37458 13268 37464 13320
rect 37516 13308 37522 13320
rect 37918 13308 37924 13320
rect 37516 13280 37924 13308
rect 37516 13268 37522 13280
rect 37918 13268 37924 13280
rect 37976 13268 37982 13320
rect 39022 13268 39028 13320
rect 39080 13308 39086 13320
rect 40589 13311 40647 13317
rect 40589 13308 40601 13311
rect 39080 13280 40601 13308
rect 39080 13268 39086 13280
rect 40589 13277 40601 13280
rect 40635 13277 40647 13311
rect 41064 13308 41092 13416
rect 42337 13413 42349 13416
rect 42383 13413 42395 13447
rect 42337 13407 42395 13413
rect 41230 13336 41236 13388
rect 41288 13376 41294 13388
rect 44085 13379 44143 13385
rect 44085 13376 44097 13379
rect 41288 13348 44097 13376
rect 41288 13336 41294 13348
rect 44085 13345 44097 13348
rect 44131 13345 44143 13379
rect 44085 13339 44143 13345
rect 41141 13311 41199 13317
rect 41141 13308 41153 13311
rect 41064 13280 41153 13308
rect 40589 13271 40647 13277
rect 41141 13277 41153 13280
rect 41187 13277 41199 13311
rect 41141 13271 41199 13277
rect 41322 13268 41328 13320
rect 41380 13308 41386 13320
rect 41380 13280 42734 13308
rect 41380 13268 41386 13280
rect 34839 13212 36492 13240
rect 36556 13212 36860 13240
rect 38626 13212 41414 13240
rect 34839 13209 34851 13212
rect 34793 13203 34851 13209
rect 34698 13172 34704 13184
rect 31726 13144 34704 13172
rect 31297 13135 31355 13141
rect 34698 13132 34704 13144
rect 34756 13132 34762 13184
rect 34882 13132 34888 13184
rect 34940 13172 34946 13184
rect 35434 13172 35440 13184
rect 34940 13144 35440 13172
rect 34940 13132 34946 13144
rect 35434 13132 35440 13144
rect 35492 13132 35498 13184
rect 36464 13172 36492 13212
rect 38626 13172 38654 13212
rect 36464 13144 38654 13172
rect 40494 13132 40500 13184
rect 40552 13132 40558 13184
rect 41386 13172 41414 13212
rect 43806 13200 43812 13252
rect 43864 13200 43870 13252
rect 44358 13172 44364 13184
rect 41386 13144 44364 13172
rect 44358 13132 44364 13144
rect 44416 13132 44422 13184
rect 1104 13082 45172 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 45172 13082
rect 1104 13008 45172 13030
rect 7929 12971 7987 12977
rect 7929 12937 7941 12971
rect 7975 12968 7987 12971
rect 9214 12968 9220 12980
rect 7975 12940 9220 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11698 12928 11704 12980
rect 11756 12928 11762 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12937 12311 12971
rect 12253 12931 12311 12937
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 7006 12900 7012 12912
rect 6871 12872 7012 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 9677 12903 9735 12909
rect 9677 12869 9689 12903
rect 9723 12900 9735 12903
rect 12066 12900 12072 12912
rect 9723 12872 12072 12900
rect 9723 12869 9735 12872
rect 9677 12863 9735 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11195 12804 11284 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7760 12764 7788 12795
rect 7331 12736 7788 12764
rect 11256 12764 11284 12804
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11606 12832 11612 12844
rect 11388 12804 11612 12832
rect 11388 12792 11394 12804
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11698 12835 11756 12841
rect 11698 12801 11710 12835
rect 11744 12832 11756 12835
rect 11974 12832 11980 12844
rect 11744 12804 11980 12832
rect 11744 12801 11756 12804
rect 11698 12795 11756 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12268 12832 12296 12931
rect 13078 12928 13084 12980
rect 13136 12928 13142 12980
rect 13179 12971 13237 12977
rect 13179 12937 13191 12971
rect 13225 12968 13237 12971
rect 13354 12968 13360 12980
rect 13225 12940 13360 12968
rect 13225 12937 13237 12940
rect 13179 12931 13237 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 14826 12968 14832 12980
rect 14783 12940 14832 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 15838 12968 15844 12980
rect 15212 12940 15844 12968
rect 13096 12900 13124 12928
rect 14844 12900 14872 12928
rect 12360 12872 12664 12900
rect 13096 12872 13216 12900
rect 14844 12872 15148 12900
rect 12360 12844 12388 12872
rect 12207 12804 12296 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12342 12792 12348 12844
rect 12400 12792 12406 12844
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 12636 12841 12664 12872
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13078 12832 13084 12844
rect 12759 12804 13084 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 12437 12767 12495 12773
rect 11256 12736 12388 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 1578 12656 1584 12708
rect 1636 12696 1642 12708
rect 7101 12699 7159 12705
rect 7101 12696 7113 12699
rect 1636 12668 7113 12696
rect 1636 12656 1642 12668
rect 7101 12665 7113 12668
rect 7147 12665 7159 12699
rect 7101 12659 7159 12665
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11379 12668 12081 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 12069 12665 12081 12668
rect 12115 12665 12127 12699
rect 12360 12696 12388 12736
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 13188 12764 13216 12872
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 12483 12736 13216 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12986 12696 12992 12708
rect 12360 12668 12992 12696
rect 12069 12659 12127 12665
rect 12986 12656 12992 12668
rect 13044 12696 13050 12708
rect 13280 12696 13308 12795
rect 13354 12792 13360 12844
rect 13412 12792 13418 12844
rect 15120 12841 15148 12872
rect 15212 12844 15240 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16482 12968 16488 12980
rect 16255 12940 16488 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 17497 12971 17555 12977
rect 16724 12940 16988 12968
rect 16724 12928 16730 12940
rect 15764 12872 16068 12900
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14476 12804 14657 12832
rect 13044 12668 13308 12696
rect 14476 12696 14504 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15105 12835 15163 12841
rect 14875 12804 15056 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14608 12736 14933 12764
rect 14608 12724 14614 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 15028 12696 15056 12804
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15427 12804 15700 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15672 12776 15700 12804
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15470 12764 15476 12776
rect 15335 12736 15476 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 15764 12696 15792 12872
rect 16040 12841 16068 12872
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 16816 12872 16896 12900
rect 16816 12860 16822 12872
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 14476 12668 14872 12696
rect 15028 12668 15792 12696
rect 13044 12656 13050 12668
rect 14844 12640 14872 12668
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 9950 12628 9956 12640
rect 9631 12600 9956 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 12434 12628 12440 12640
rect 11664 12600 12440 12628
rect 11664 12588 11670 12600
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13722 12628 13728 12640
rect 12584 12600 13728 12628
rect 12584 12588 12590 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15856 12628 15884 12795
rect 16040 12764 16068 12795
rect 16666 12792 16672 12844
rect 16724 12792 16730 12844
rect 16868 12841 16896 12872
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16960 12832 16988 12940
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 18782 12968 18788 12980
rect 17543 12940 18788 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 19484 12940 19625 12968
rect 19484 12928 19490 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 19889 12971 19947 12977
rect 19889 12937 19901 12971
rect 19935 12968 19947 12971
rect 20162 12968 20168 12980
rect 19935 12940 20168 12968
rect 19935 12937 19947 12940
rect 19889 12931 19947 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21910 12968 21916 12980
rect 21131 12940 21916 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22741 12971 22799 12977
rect 22741 12968 22753 12971
rect 22152 12940 22753 12968
rect 22152 12928 22158 12940
rect 22741 12937 22753 12940
rect 22787 12937 22799 12971
rect 22741 12931 22799 12937
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 25317 12971 25375 12977
rect 25317 12968 25329 12971
rect 23256 12940 25329 12968
rect 23256 12928 23262 12940
rect 25317 12937 25329 12940
rect 25363 12937 25375 12971
rect 25317 12931 25375 12937
rect 25774 12928 25780 12980
rect 25832 12928 25838 12980
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 27246 12968 27252 12980
rect 26292 12940 27252 12968
rect 26292 12928 26298 12940
rect 27246 12928 27252 12940
rect 27304 12928 27310 12980
rect 28902 12928 28908 12980
rect 28960 12928 28966 12980
rect 29270 12928 29276 12980
rect 29328 12968 29334 12980
rect 29457 12971 29515 12977
rect 29457 12968 29469 12971
rect 29328 12940 29469 12968
rect 29328 12928 29334 12940
rect 29457 12937 29469 12940
rect 29503 12937 29515 12971
rect 31846 12968 31852 12980
rect 29457 12931 29515 12937
rect 31036 12940 31852 12968
rect 17773 12903 17831 12909
rect 17773 12869 17785 12903
rect 17819 12900 17831 12903
rect 18325 12903 18383 12909
rect 18325 12900 18337 12903
rect 17819 12872 18000 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 17635 12835 17693 12841
rect 17635 12832 17647 12835
rect 16960 12804 17647 12832
rect 16853 12795 16911 12801
rect 17635 12801 17647 12804
rect 17681 12801 17693 12835
rect 17635 12795 17693 12801
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 16040 12736 16712 12764
rect 16684 12640 16712 12736
rect 17972 12696 18000 12872
rect 18064 12872 18337 12900
rect 18064 12841 18092 12872
rect 18325 12869 18337 12872
rect 18371 12869 18383 12903
rect 18325 12863 18383 12869
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19208 12872 19809 12900
rect 19208 12860 19214 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 23569 12903 23627 12909
rect 23569 12900 23581 12903
rect 19797 12863 19855 12869
rect 19996 12872 20668 12900
rect 18048 12835 18106 12841
rect 18048 12801 18060 12835
rect 18094 12801 18106 12835
rect 18048 12795 18106 12801
rect 18141 12835 18199 12841
rect 18141 12801 18153 12835
rect 18187 12832 18199 12835
rect 18230 12832 18236 12844
rect 18187 12804 18236 12832
rect 18187 12801 18199 12804
rect 18141 12795 18199 12801
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 18598 12832 18604 12844
rect 18463 12804 18604 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 19518 12792 19524 12844
rect 19576 12792 19582 12844
rect 18690 12724 18696 12776
rect 18748 12764 18754 12776
rect 19150 12764 19156 12776
rect 18748 12736 19156 12764
rect 18748 12724 18754 12736
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19996 12764 20024 12872
rect 20254 12792 20260 12844
rect 20312 12792 20318 12844
rect 20530 12792 20536 12844
rect 20588 12792 20594 12844
rect 20640 12841 20668 12872
rect 22066 12872 23581 12900
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20806 12792 20812 12844
rect 20864 12792 20870 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 19812 12736 20024 12764
rect 18322 12696 18328 12708
rect 17972 12668 18328 12696
rect 18322 12656 18328 12668
rect 18380 12696 18386 12708
rect 19812 12705 19840 12736
rect 20070 12724 20076 12776
rect 20128 12724 20134 12776
rect 20165 12767 20223 12773
rect 20165 12733 20177 12767
rect 20211 12733 20223 12767
rect 20165 12727 20223 12733
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12764 20407 12767
rect 22066 12764 22094 12872
rect 23569 12869 23581 12872
rect 23615 12869 23627 12903
rect 23569 12863 23627 12869
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 23808 12872 23980 12900
rect 23808 12860 23814 12872
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 20395 12736 22094 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 19797 12699 19855 12705
rect 18380 12668 18828 12696
rect 18380 12656 18386 12668
rect 18800 12640 18828 12668
rect 19797 12665 19809 12699
rect 19843 12665 19855 12699
rect 20180 12696 20208 12727
rect 20438 12696 20444 12708
rect 20180 12668 20444 12696
rect 19797 12659 19855 12665
rect 20438 12656 20444 12668
rect 20496 12656 20502 12708
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 22296 12696 22324 12795
rect 23014 12792 23020 12844
rect 23072 12832 23078 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 23072 12804 23121 12832
rect 23072 12792 23078 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 23842 12792 23848 12844
rect 23900 12792 23906 12844
rect 23952 12841 23980 12872
rect 24946 12860 24952 12912
rect 25004 12860 25010 12912
rect 25222 12860 25228 12912
rect 25280 12900 25286 12912
rect 25685 12903 25743 12909
rect 25685 12900 25697 12903
rect 25280 12872 25697 12900
rect 25280 12860 25286 12872
rect 25685 12869 25697 12872
rect 25731 12900 25743 12903
rect 27709 12903 27767 12909
rect 27709 12900 27721 12903
rect 25731 12872 27721 12900
rect 25731 12869 25743 12872
rect 25685 12863 25743 12869
rect 27709 12869 27721 12872
rect 27755 12869 27767 12903
rect 27709 12863 27767 12869
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 24026 12792 24032 12844
rect 24084 12792 24090 12844
rect 24213 12835 24271 12841
rect 24213 12801 24225 12835
rect 24259 12832 24271 12835
rect 24302 12832 24308 12844
rect 24259 12804 24308 12832
rect 24259 12801 24271 12804
rect 24213 12795 24271 12801
rect 23382 12724 23388 12776
rect 23440 12724 23446 12776
rect 24228 12696 24256 12795
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 24964 12832 24992 12860
rect 27154 12832 27160 12844
rect 24964 12804 27160 12832
rect 27154 12792 27160 12804
rect 27212 12832 27218 12844
rect 27433 12835 27491 12841
rect 27433 12832 27445 12835
rect 27212 12804 27445 12832
rect 27212 12792 27218 12804
rect 27433 12801 27445 12804
rect 27479 12801 27491 12835
rect 27433 12795 27491 12801
rect 25038 12724 25044 12776
rect 25096 12724 25102 12776
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 25866 12764 25872 12776
rect 25464 12736 25872 12764
rect 25464 12724 25470 12736
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 27709 12767 27767 12773
rect 27709 12733 27721 12767
rect 27755 12764 27767 12767
rect 28920 12764 28948 12928
rect 29638 12792 29644 12844
rect 29696 12792 29702 12844
rect 31036 12841 31064 12940
rect 31846 12928 31852 12940
rect 31904 12928 31910 12980
rect 34698 12928 34704 12980
rect 34756 12968 34762 12980
rect 35342 12968 35348 12980
rect 34756 12940 35348 12968
rect 34756 12928 34762 12940
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 35618 12928 35624 12980
rect 35676 12968 35682 12980
rect 37090 12968 37096 12980
rect 35676 12940 37096 12968
rect 35676 12928 35682 12940
rect 37090 12928 37096 12940
rect 37148 12928 37154 12980
rect 37918 12928 37924 12980
rect 37976 12968 37982 12980
rect 38933 12971 38991 12977
rect 38933 12968 38945 12971
rect 37976 12940 38945 12968
rect 37976 12928 37982 12940
rect 38933 12937 38945 12940
rect 38979 12937 38991 12971
rect 38933 12931 38991 12937
rect 40494 12928 40500 12980
rect 40552 12928 40558 12980
rect 43533 12971 43591 12977
rect 43533 12937 43545 12971
rect 43579 12968 43591 12971
rect 43806 12968 43812 12980
rect 43579 12940 43812 12968
rect 43579 12937 43591 12940
rect 43533 12931 43591 12937
rect 43806 12928 43812 12940
rect 43864 12928 43870 12980
rect 31754 12900 31760 12912
rect 31128 12872 31340 12900
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12801 31079 12835
rect 31021 12795 31079 12801
rect 27755 12736 28948 12764
rect 27755 12733 27767 12736
rect 27709 12727 27767 12733
rect 29822 12724 29828 12776
rect 29880 12724 29886 12776
rect 30466 12724 30472 12776
rect 30524 12764 30530 12776
rect 31128 12764 31156 12872
rect 31312 12841 31340 12872
rect 31496 12872 31760 12900
rect 31496 12841 31524 12872
rect 31754 12860 31760 12872
rect 31812 12860 31818 12912
rect 35360 12900 35388 12928
rect 40405 12903 40463 12909
rect 32140 12872 32904 12900
rect 35360 12886 39238 12900
rect 35360 12872 39252 12886
rect 31205 12835 31263 12841
rect 31205 12801 31217 12835
rect 31251 12801 31263 12835
rect 31205 12795 31263 12801
rect 31297 12835 31355 12841
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 31481 12835 31539 12841
rect 31481 12801 31493 12835
rect 31527 12801 31539 12835
rect 31846 12832 31852 12844
rect 31481 12795 31539 12801
rect 31588 12804 31852 12832
rect 30524 12736 31156 12764
rect 31220 12764 31248 12795
rect 31588 12764 31616 12804
rect 31846 12792 31852 12804
rect 31904 12832 31910 12844
rect 32140 12832 32168 12872
rect 31904 12804 32168 12832
rect 32217 12835 32275 12841
rect 31904 12792 31910 12804
rect 32217 12801 32229 12835
rect 32263 12801 32275 12835
rect 32217 12795 32275 12801
rect 32401 12835 32459 12841
rect 32401 12801 32413 12835
rect 32447 12832 32459 12835
rect 32490 12832 32496 12844
rect 32447 12804 32496 12832
rect 32447 12801 32459 12804
rect 32401 12795 32459 12801
rect 31220 12736 31616 12764
rect 30524 12724 30530 12736
rect 31754 12724 31760 12776
rect 31812 12764 31818 12776
rect 32232 12764 32260 12795
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 32674 12792 32680 12844
rect 32732 12792 32738 12844
rect 32876 12841 32904 12872
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12801 32827 12835
rect 32769 12795 32827 12801
rect 32861 12835 32919 12841
rect 32861 12801 32873 12835
rect 32907 12801 32919 12835
rect 32861 12795 32919 12801
rect 31812 12736 32260 12764
rect 31812 12724 31818 12736
rect 21416 12668 24256 12696
rect 21416 12656 21422 12668
rect 24394 12656 24400 12708
rect 24452 12656 24458 12708
rect 24486 12656 24492 12708
rect 24544 12696 24550 12708
rect 25056 12696 25084 12724
rect 28994 12696 29000 12708
rect 24544 12668 25084 12696
rect 27448 12668 29000 12696
rect 24544 12656 24550 12668
rect 16114 12628 16120 12640
rect 14884 12600 16120 12628
rect 14884 12588 14890 12600
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 17034 12588 17040 12640
rect 17092 12588 17098 12640
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 19518 12628 19524 12640
rect 18840 12600 19524 12628
rect 18840 12588 18846 12600
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 22462 12628 22468 12640
rect 20588 12600 22468 12628
rect 20588 12588 20594 12600
rect 22462 12588 22468 12600
rect 22520 12588 22526 12640
rect 24412 12628 24440 12656
rect 27448 12628 27476 12668
rect 28994 12656 29000 12668
rect 29052 12656 29058 12708
rect 30837 12699 30895 12705
rect 30837 12665 30849 12699
rect 30883 12696 30895 12699
rect 31294 12696 31300 12708
rect 30883 12668 31300 12696
rect 30883 12665 30895 12668
rect 30837 12659 30895 12665
rect 31294 12656 31300 12668
rect 31352 12696 31358 12708
rect 31665 12699 31723 12705
rect 31665 12696 31677 12699
rect 31352 12668 31677 12696
rect 31352 12656 31358 12668
rect 31665 12665 31677 12668
rect 31711 12665 31723 12699
rect 31665 12659 31723 12665
rect 24412 12600 27476 12628
rect 27525 12631 27583 12637
rect 27525 12597 27537 12631
rect 27571 12628 27583 12631
rect 27614 12628 27620 12640
rect 27571 12600 27620 12628
rect 27571 12597 27583 12600
rect 27525 12591 27583 12597
rect 27614 12588 27620 12600
rect 27672 12628 27678 12640
rect 30742 12628 30748 12640
rect 27672 12600 30748 12628
rect 27672 12588 27678 12600
rect 30742 12588 30748 12600
rect 30800 12588 30806 12640
rect 31570 12588 31576 12640
rect 31628 12628 31634 12640
rect 31754 12628 31760 12640
rect 31628 12600 31760 12628
rect 31628 12588 31634 12600
rect 31754 12588 31760 12600
rect 31812 12628 31818 12640
rect 32784 12628 32812 12795
rect 34698 12792 34704 12844
rect 34756 12832 34762 12844
rect 34882 12832 34888 12844
rect 34756 12804 34888 12832
rect 34756 12792 34762 12804
rect 34882 12792 34888 12804
rect 34940 12792 34946 12844
rect 39224 12764 39252 12872
rect 40405 12869 40417 12903
rect 40451 12900 40463 12903
rect 40512 12900 40540 12928
rect 40451 12872 40540 12900
rect 40451 12869 40463 12872
rect 40405 12863 40463 12869
rect 44358 12860 44364 12912
rect 44416 12860 44422 12912
rect 43349 12835 43407 12841
rect 43349 12801 43361 12835
rect 43395 12832 43407 12835
rect 43395 12804 43944 12832
rect 43395 12801 43407 12804
rect 43349 12795 43407 12801
rect 39224 12736 40632 12764
rect 40604 12696 40632 12736
rect 40678 12724 40684 12776
rect 40736 12724 40742 12776
rect 43916 12773 43944 12804
rect 43901 12767 43959 12773
rect 43901 12733 43913 12767
rect 43947 12733 43959 12767
rect 43901 12727 43959 12733
rect 41322 12696 41328 12708
rect 40604 12668 41328 12696
rect 41322 12656 41328 12668
rect 41380 12656 41386 12708
rect 44085 12699 44143 12705
rect 44085 12665 44097 12699
rect 44131 12696 44143 12699
rect 44634 12696 44640 12708
rect 44131 12668 44640 12696
rect 44131 12665 44143 12668
rect 44085 12659 44143 12665
rect 44634 12656 44640 12668
rect 44692 12656 44698 12708
rect 31812 12600 32812 12628
rect 31812 12588 31818 12600
rect 1104 12538 45172 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 45172 12538
rect 1104 12464 45172 12486
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12250 12424 12256 12436
rect 11931 12396 12256 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 13078 12424 13084 12436
rect 12360 12396 13084 12424
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 12360 12356 12388 12396
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13228 12396 13645 12424
rect 13228 12384 13234 12396
rect 13633 12393 13645 12396
rect 13679 12424 13691 12427
rect 13998 12424 14004 12436
rect 13679 12396 14004 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14918 12424 14924 12436
rect 14148 12396 14924 12424
rect 14148 12384 14154 12396
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 15102 12384 15108 12436
rect 15160 12384 15166 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 15344 12396 15393 12424
rect 15344 12384 15350 12396
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 15381 12387 15439 12393
rect 12032 12328 12388 12356
rect 12032 12316 12038 12328
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 13722 12356 13728 12368
rect 12492 12328 13728 12356
rect 12492 12316 12498 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 14369 12359 14427 12365
rect 14369 12325 14381 12359
rect 14415 12356 14427 12359
rect 15194 12356 15200 12368
rect 14415 12328 15200 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 15396 12356 15424 12387
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 17405 12427 17463 12433
rect 15528 12396 17356 12424
rect 15528 12384 15534 12396
rect 15396 12328 15516 12356
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12299 12260 12664 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 11839 12192 12081 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 12069 12189 12081 12192
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12526 12220 12532 12232
rect 12391 12192 12532 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 11517 12155 11575 12161
rect 11517 12121 11529 12155
rect 11563 12152 11575 12155
rect 11606 12152 11612 12164
rect 11563 12124 11612 12152
rect 11563 12121 11575 12124
rect 11517 12115 11575 12121
rect 11606 12112 11612 12124
rect 11664 12112 11670 12164
rect 11701 12155 11759 12161
rect 11701 12121 11713 12155
rect 11747 12152 11759 12155
rect 11882 12152 11888 12164
rect 11747 12124 11888 12152
rect 11747 12121 11759 12124
rect 11701 12115 11759 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 12084 12152 12112 12183
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 12636 12229 12664 12260
rect 14936 12260 15424 12288
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 12667 12192 12848 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 12820 12152 12848 12192
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 12952 12192 13400 12220
rect 12952 12180 12958 12192
rect 12084 12124 12572 12152
rect 12820 12124 12940 12152
rect 12544 12096 12572 12124
rect 12912 12096 12940 12124
rect 13372 12096 13400 12192
rect 13464 12192 13553 12220
rect 13464 12096 13492 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 13998 12220 14004 12232
rect 13771 12192 14004 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 14274 12220 14280 12232
rect 14231 12192 14280 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 14642 12180 14648 12232
rect 14700 12180 14706 12232
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 14936 12229 14964 12260
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 14844 12152 14872 12183
rect 14476 12124 14872 12152
rect 14936 12152 14964 12183
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 15396 12229 15424 12260
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15102 12152 15108 12164
rect 14936 12124 15108 12152
rect 14476 12096 14504 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15488 12152 15516 12328
rect 15654 12316 15660 12368
rect 15712 12316 15718 12368
rect 15764 12328 16160 12356
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15672 12220 15700 12316
rect 15764 12297 15792 12328
rect 16132 12300 16160 12328
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17221 12359 17279 12365
rect 17221 12356 17233 12359
rect 17092 12328 17233 12356
rect 17092 12316 17098 12328
rect 17221 12325 17233 12328
rect 17267 12325 17279 12359
rect 17328 12356 17356 12396
rect 17405 12393 17417 12427
rect 17451 12424 17463 12427
rect 20809 12427 20867 12433
rect 17451 12396 17954 12424
rect 17451 12393 17463 12396
rect 17405 12387 17463 12393
rect 17497 12359 17555 12365
rect 17497 12356 17509 12359
rect 17328 12328 17509 12356
rect 17221 12319 17279 12325
rect 17497 12325 17509 12328
rect 17543 12325 17555 12359
rect 17497 12319 17555 12325
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16114 12248 16120 12300
rect 16172 12248 16178 12300
rect 17310 12288 17316 12300
rect 16500 12260 17316 12288
rect 16500 12232 16528 12260
rect 17310 12248 17316 12260
rect 17368 12288 17374 12300
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 17368 12260 17417 12288
rect 17368 12248 17374 12260
rect 17405 12257 17417 12260
rect 17451 12257 17463 12291
rect 17926 12288 17954 12396
rect 20809 12393 20821 12427
rect 20855 12424 20867 12427
rect 20898 12424 20904 12436
rect 20855 12396 20904 12424
rect 20855 12393 20867 12396
rect 20809 12387 20867 12393
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21174 12384 21180 12436
rect 21232 12384 21238 12436
rect 22465 12427 22523 12433
rect 22465 12393 22477 12427
rect 22511 12424 22523 12427
rect 22830 12424 22836 12436
rect 22511 12396 22836 12424
rect 22511 12393 22523 12396
rect 22465 12387 22523 12393
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 28445 12427 28503 12433
rect 28445 12424 28457 12427
rect 27764 12396 28457 12424
rect 27764 12384 27770 12396
rect 28445 12393 28457 12396
rect 28491 12393 28503 12427
rect 28445 12387 28503 12393
rect 29638 12384 29644 12436
rect 29696 12424 29702 12436
rect 30101 12427 30159 12433
rect 30101 12424 30113 12427
rect 29696 12396 30113 12424
rect 29696 12384 29702 12396
rect 30101 12393 30113 12396
rect 30147 12393 30159 12427
rect 30101 12387 30159 12393
rect 30742 12384 30748 12436
rect 30800 12384 30806 12436
rect 32490 12424 32496 12436
rect 31036 12396 32496 12424
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19392 12328 20208 12356
rect 19392 12316 19398 12328
rect 17926 12260 19380 12288
rect 17405 12251 17463 12257
rect 15611 12192 15700 12220
rect 15841 12223 15899 12229
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15856 12152 15884 12183
rect 15930 12180 15936 12232
rect 15988 12180 15994 12232
rect 16206 12220 16212 12232
rect 16132 12210 16212 12220
rect 16040 12207 16212 12210
rect 16037 12201 16212 12207
rect 16037 12167 16049 12201
rect 16083 12192 16212 12201
rect 16083 12182 16160 12192
rect 16083 12167 16095 12182
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17000 12192 17601 12220
rect 17000 12180 17006 12192
rect 17589 12189 17601 12192
rect 17635 12189 17647 12223
rect 18598 12220 18604 12232
rect 17589 12183 17647 12189
rect 17696 12192 18604 12220
rect 16037 12161 16095 12167
rect 15488 12124 15884 12152
rect 16224 12152 16252 12180
rect 17696 12152 17724 12192
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 16224 12124 17724 12152
rect 19352 12096 19380 12260
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19484 12260 19932 12288
rect 19484 12248 19490 12260
rect 19904 12232 19932 12260
rect 19518 12180 19524 12232
rect 19576 12180 19582 12232
rect 19702 12180 19708 12232
rect 19760 12180 19766 12232
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20180 12229 20208 12328
rect 20622 12316 20628 12368
rect 20680 12316 20686 12368
rect 21637 12359 21695 12365
rect 21637 12325 21649 12359
rect 21683 12325 21695 12359
rect 21637 12319 21695 12325
rect 20441 12291 20499 12297
rect 20441 12257 20453 12291
rect 20487 12288 20499 12291
rect 20640 12288 20668 12316
rect 20487 12260 20668 12288
rect 20487 12257 20499 12260
rect 20441 12251 20499 12257
rect 21358 12248 21364 12300
rect 21416 12248 21422 12300
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 20036 12192 20085 12220
rect 20036 12180 20042 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 20254 12220 20260 12232
rect 20211 12192 20260 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 19536 12152 19564 12180
rect 19797 12155 19855 12161
rect 19797 12152 19809 12155
rect 19536 12124 19809 12152
rect 19797 12121 19809 12124
rect 19843 12121 19855 12155
rect 20088 12152 20116 12183
rect 20254 12180 20260 12192
rect 20312 12180 20318 12232
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20364 12152 20392 12183
rect 20530 12180 20536 12232
rect 20588 12180 20594 12232
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20088 12124 20392 12152
rect 20640 12152 20668 12183
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 21453 12223 21511 12229
rect 21453 12220 21465 12223
rect 20864 12192 21465 12220
rect 20864 12180 20870 12192
rect 21453 12189 21465 12192
rect 21499 12189 21511 12223
rect 21652 12220 21680 12319
rect 21726 12316 21732 12368
rect 21784 12356 21790 12368
rect 22649 12359 22707 12365
rect 22649 12356 22661 12359
rect 21784 12328 22661 12356
rect 21784 12316 21790 12328
rect 22649 12325 22661 12328
rect 22695 12325 22707 12359
rect 22649 12319 22707 12325
rect 23106 12248 23112 12300
rect 23164 12248 23170 12300
rect 23293 12291 23351 12297
rect 23293 12257 23305 12291
rect 23339 12288 23351 12291
rect 23750 12288 23756 12300
rect 23339 12260 23756 12288
rect 23339 12257 23351 12260
rect 23293 12251 23351 12257
rect 23750 12248 23756 12260
rect 23808 12248 23814 12300
rect 30484 12260 30696 12288
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 21652 12192 22385 12220
rect 21453 12183 21511 12189
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 22557 12223 22615 12229
rect 22557 12189 22569 12223
rect 22603 12220 22615 12223
rect 22922 12220 22928 12232
rect 22603 12192 22928 12220
rect 22603 12189 22615 12192
rect 22557 12183 22615 12189
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 28350 12180 28356 12232
rect 28408 12180 28414 12232
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12220 28595 12223
rect 28994 12220 29000 12232
rect 28583 12192 29000 12220
rect 28583 12189 28595 12192
rect 28537 12183 28595 12189
rect 28994 12180 29000 12192
rect 29052 12180 29058 12232
rect 29086 12180 29092 12232
rect 29144 12220 29150 12232
rect 29454 12220 29460 12232
rect 29144 12192 29460 12220
rect 29144 12180 29150 12192
rect 29454 12180 29460 12192
rect 29512 12220 29518 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29512 12192 29745 12220
rect 29512 12180 29518 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 30285 12223 30343 12229
rect 30285 12189 30297 12223
rect 30331 12189 30343 12223
rect 30285 12183 30343 12189
rect 21177 12155 21235 12161
rect 21177 12152 21189 12155
rect 20640 12124 21189 12152
rect 19797 12115 19855 12121
rect 20640 12096 20668 12124
rect 21177 12121 21189 12124
rect 21223 12121 21235 12155
rect 21177 12115 21235 12121
rect 29914 12112 29920 12164
rect 29972 12112 29978 12164
rect 30300 12152 30328 12183
rect 30374 12180 30380 12232
rect 30432 12180 30438 12232
rect 30484 12229 30512 12260
rect 30668 12232 30696 12260
rect 30469 12223 30527 12229
rect 30469 12189 30481 12223
rect 30515 12189 30527 12223
rect 30469 12183 30527 12189
rect 30558 12180 30564 12232
rect 30616 12180 30622 12232
rect 30650 12180 30656 12232
rect 30708 12180 30714 12232
rect 31036 12229 31064 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 36078 12384 36084 12436
rect 36136 12384 36142 12436
rect 32398 12356 32404 12368
rect 31312 12328 32404 12356
rect 30897 12223 30955 12229
rect 30897 12220 30909 12223
rect 30760 12192 30909 12220
rect 30760 12164 30788 12192
rect 30897 12189 30909 12192
rect 30943 12189 30955 12223
rect 30897 12183 30955 12189
rect 31021 12223 31079 12229
rect 31021 12189 31033 12223
rect 31067 12189 31079 12223
rect 31021 12183 31079 12189
rect 31113 12223 31171 12229
rect 31113 12189 31125 12223
rect 31159 12220 31171 12223
rect 31202 12220 31208 12232
rect 31159 12192 31208 12220
rect 31159 12189 31171 12192
rect 31113 12183 31171 12189
rect 31202 12180 31208 12192
rect 31260 12180 31266 12232
rect 31312 12229 31340 12328
rect 32398 12316 32404 12328
rect 32456 12316 32462 12368
rect 34606 12316 34612 12368
rect 34664 12356 34670 12368
rect 34793 12359 34851 12365
rect 34793 12356 34805 12359
rect 34664 12328 34805 12356
rect 34664 12316 34670 12328
rect 34793 12325 34805 12328
rect 34839 12325 34851 12359
rect 34793 12319 34851 12325
rect 31386 12248 31392 12300
rect 31444 12288 31450 12300
rect 35161 12291 35219 12297
rect 31444 12260 32076 12288
rect 31444 12248 31450 12260
rect 31297 12223 31355 12229
rect 31297 12189 31309 12223
rect 31343 12189 31355 12223
rect 31297 12183 31355 12189
rect 31387 12201 31445 12207
rect 31387 12167 31399 12201
rect 31433 12167 31445 12201
rect 31478 12180 31484 12232
rect 31536 12180 31542 12232
rect 31662 12180 31668 12232
rect 31720 12180 31726 12232
rect 31754 12180 31760 12232
rect 31812 12220 31818 12232
rect 32048 12229 32076 12260
rect 35161 12257 35173 12291
rect 35207 12288 35219 12291
rect 37458 12288 37464 12300
rect 35207 12260 37464 12288
rect 35207 12257 35219 12260
rect 35161 12251 35219 12257
rect 37458 12248 37464 12260
rect 37516 12248 37522 12300
rect 37826 12248 37832 12300
rect 37884 12248 37890 12300
rect 31849 12223 31907 12229
rect 31849 12220 31861 12223
rect 31812 12192 31861 12220
rect 31812 12180 31818 12192
rect 31849 12189 31861 12192
rect 31895 12189 31907 12223
rect 31849 12183 31907 12189
rect 31941 12223 31999 12229
rect 31941 12189 31953 12223
rect 31987 12189 31999 12223
rect 31941 12183 31999 12189
rect 32033 12223 32091 12229
rect 32033 12189 32045 12223
rect 32079 12220 32091 12223
rect 32122 12220 32128 12232
rect 32079 12192 32128 12220
rect 32079 12189 32091 12192
rect 32033 12183 32091 12189
rect 31387 12164 31445 12167
rect 30742 12152 30748 12164
rect 30300 12124 30748 12152
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 31386 12112 31392 12164
rect 31444 12112 31450 12164
rect 31496 12152 31524 12180
rect 31956 12152 31984 12183
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 32214 12180 32220 12232
rect 32272 12180 32278 12232
rect 31496 12124 31984 12152
rect 36998 12112 37004 12164
rect 37056 12112 37062 12164
rect 37553 12155 37611 12161
rect 37553 12121 37565 12155
rect 37599 12152 37611 12155
rect 39022 12152 39028 12164
rect 37599 12124 39028 12152
rect 37599 12121 37611 12124
rect 37553 12115 37611 12121
rect 39022 12112 39028 12124
rect 39080 12112 39086 12164
rect 11790 12044 11796 12096
rect 11848 12044 11854 12096
rect 12526 12044 12532 12096
rect 12584 12044 12590 12096
rect 12802 12044 12808 12096
rect 12860 12044 12866 12096
rect 12894 12044 12900 12096
rect 12952 12044 12958 12096
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 13446 12044 13452 12096
rect 13504 12044 13510 12096
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15470 12084 15476 12096
rect 14976 12056 15476 12084
rect 14976 12044 14982 12056
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18506 12084 18512 12096
rect 18288 12056 18512 12084
rect 18288 12044 18294 12056
rect 18506 12044 18512 12056
rect 18564 12084 18570 12096
rect 18966 12084 18972 12096
rect 18564 12056 18972 12084
rect 18564 12044 18570 12056
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19334 12044 19340 12096
rect 19392 12044 19398 12096
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 20162 12084 20168 12096
rect 19567 12056 20168 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20622 12044 20628 12096
rect 20680 12044 20686 12096
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 22796 12056 23029 12084
rect 22796 12044 22802 12056
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 23017 12047 23075 12053
rect 28810 12044 28816 12096
rect 28868 12084 28874 12096
rect 29549 12087 29607 12093
rect 29549 12084 29561 12087
rect 28868 12056 29561 12084
rect 28868 12044 28874 12056
rect 29549 12053 29561 12056
rect 29595 12053 29607 12087
rect 29932 12084 29960 12112
rect 30282 12084 30288 12096
rect 29932 12056 30288 12084
rect 29549 12047 29607 12053
rect 30282 12044 30288 12056
rect 30340 12044 30346 12096
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 31260 12056 31493 12084
rect 31260 12044 31266 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31481 12047 31539 12053
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 34701 12087 34759 12093
rect 34701 12084 34713 12087
rect 34664 12056 34713 12084
rect 34664 12044 34670 12056
rect 34701 12053 34713 12056
rect 34747 12053 34759 12087
rect 34701 12047 34759 12053
rect 1104 11994 45172 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 45172 11994
rect 1104 11920 45172 11942
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11698 11880 11704 11892
rect 11563 11852 11704 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 12710 11880 12716 11892
rect 12575 11852 12716 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13810 11883 13868 11889
rect 13810 11849 13822 11883
rect 13856 11880 13868 11883
rect 13906 11880 13912 11892
rect 13856 11852 13912 11880
rect 13856 11849 13868 11852
rect 13810 11843 13868 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14366 11840 14372 11892
rect 14424 11840 14430 11892
rect 14734 11840 14740 11892
rect 14792 11840 14798 11892
rect 14829 11883 14887 11889
rect 14829 11849 14841 11883
rect 14875 11880 14887 11883
rect 15010 11880 15016 11892
rect 14875 11852 15016 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15105 11883 15163 11889
rect 15105 11849 15117 11883
rect 15151 11849 15163 11883
rect 15105 11843 15163 11849
rect 14384 11812 14412 11840
rect 11808 11784 14412 11812
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11480 11716 11713 11744
rect 11480 11704 11486 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11808 11685 11836 11784
rect 14550 11772 14556 11824
rect 14608 11772 14614 11824
rect 14752 11812 14780 11840
rect 15120 11812 15148 11843
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 18414 11880 18420 11892
rect 15436 11852 18420 11880
rect 15436 11840 15442 11852
rect 18414 11840 18420 11852
rect 18472 11880 18478 11892
rect 18472 11852 18936 11880
rect 18472 11840 18478 11852
rect 14752 11784 15148 11812
rect 18908 11812 18936 11852
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19024 11852 19472 11880
rect 19024 11840 19030 11852
rect 18908 11784 19012 11812
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12303 11716 12357 11744
rect 12345 11713 12357 11716
rect 12391 11744 12403 11747
rect 12802 11744 12808 11756
rect 12391 11716 12808 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11664 11648 11805 11676
rect 11664 11636 11670 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11676 12035 11679
rect 12066 11676 12072 11688
rect 12023 11648 12072 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 11900 11608 11928 11639
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12360 11608 12388 11707
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 13630 11744 13636 11756
rect 12860 11716 13636 11744
rect 12860 11704 12866 11716
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 13814 11744 13820 11756
rect 13771 11716 13820 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 14182 11744 14188 11756
rect 13955 11716 14188 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14458 11704 14464 11756
rect 14516 11704 14522 11756
rect 14568 11744 14596 11772
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14568 11716 14933 11744
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15286 11744 15292 11756
rect 15151 11716 15292 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14056 11648 14565 11676
rect 14056 11636 14062 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 15120 11676 15148 11707
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 18512 11754 18570 11759
rect 18512 11753 18644 11754
rect 18984 11753 19012 11784
rect 19150 11772 19156 11824
rect 19208 11772 19214 11824
rect 18233 11747 18291 11753
rect 18233 11744 18245 11747
rect 17000 11716 18245 11744
rect 17000 11704 17006 11716
rect 18233 11713 18245 11716
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18512 11719 18524 11753
rect 18558 11726 18644 11753
rect 18558 11719 18570 11726
rect 18512 11713 18570 11719
rect 18417 11707 18475 11713
rect 18432 11676 18460 11707
rect 18616 11688 18644 11726
rect 18694 11747 18752 11753
rect 18694 11713 18706 11747
rect 18740 11734 18752 11747
rect 18969 11747 19027 11753
rect 18740 11713 18828 11734
rect 18694 11707 18828 11713
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 19168 11744 19196 11772
rect 19245 11747 19303 11753
rect 19245 11744 19257 11747
rect 19168 11716 19257 11744
rect 18969 11707 19027 11713
rect 19245 11713 19257 11716
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19444 11744 19472 11852
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19889 11883 19947 11889
rect 19576 11852 19656 11880
rect 19576 11840 19582 11852
rect 19628 11821 19656 11852
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20070 11880 20076 11892
rect 19935 11852 20076 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20162 11840 20168 11892
rect 20220 11840 20226 11892
rect 20438 11840 20444 11892
rect 20496 11840 20502 11892
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 23934 11880 23940 11892
rect 23624 11852 23940 11880
rect 23624 11840 23630 11852
rect 23934 11840 23940 11852
rect 23992 11880 23998 11892
rect 24765 11883 24823 11889
rect 24765 11880 24777 11883
rect 23992 11852 24777 11880
rect 23992 11840 23998 11852
rect 24765 11849 24777 11852
rect 24811 11849 24823 11883
rect 24765 11843 24823 11849
rect 25222 11840 25228 11892
rect 25280 11840 25286 11892
rect 27062 11840 27068 11892
rect 27120 11840 27126 11892
rect 29822 11840 29828 11892
rect 29880 11880 29886 11892
rect 29917 11883 29975 11889
rect 29917 11880 29929 11883
rect 29880 11852 29929 11880
rect 29880 11840 29886 11852
rect 29917 11849 29929 11852
rect 29963 11849 29975 11883
rect 29917 11843 29975 11849
rect 30558 11840 30564 11892
rect 30616 11880 30622 11892
rect 31113 11883 31171 11889
rect 31113 11880 31125 11883
rect 30616 11852 31125 11880
rect 30616 11840 30622 11852
rect 31113 11849 31125 11852
rect 31159 11849 31171 11883
rect 31113 11843 31171 11849
rect 19613 11815 19671 11821
rect 19613 11781 19625 11815
rect 19659 11781 19671 11815
rect 20180 11812 20208 11840
rect 19613 11775 19671 11781
rect 19812 11784 20116 11812
rect 20180 11784 20300 11812
rect 19521 11747 19579 11753
rect 19521 11744 19533 11747
rect 19444 11716 19533 11744
rect 18708 11706 18828 11707
rect 14553 11639 14611 11645
rect 14660 11648 15148 11676
rect 17972 11648 18460 11676
rect 11716 11580 12388 11608
rect 11716 11552 11744 11580
rect 13078 11568 13084 11620
rect 13136 11608 13142 11620
rect 14660 11608 14688 11648
rect 13136 11580 14688 11608
rect 13136 11568 13142 11580
rect 17972 11552 18000 11648
rect 18432 11608 18460 11648
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 18800 11676 18828 11706
rect 18708 11648 18828 11676
rect 18877 11679 18935 11685
rect 18708 11608 18736 11648
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 19153 11679 19211 11685
rect 18923 11648 19012 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 18984 11620 19012 11648
rect 19153 11645 19165 11679
rect 19199 11676 19211 11679
rect 19352 11676 19380 11707
rect 19199 11648 19380 11676
rect 19444 11676 19472 11716
rect 19521 11713 19533 11716
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 19702 11704 19708 11756
rect 19760 11704 19766 11756
rect 19812 11676 19840 11784
rect 20088 11753 20116 11784
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20162 11744 20168 11756
rect 20119 11716 20168 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 19444 11648 19840 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 18432 11580 18736 11608
rect 18785 11611 18843 11617
rect 18785 11577 18797 11611
rect 18831 11577 18843 11611
rect 18785 11571 18843 11577
rect 11698 11500 11704 11552
rect 11756 11500 11762 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 13872 11512 14657 11540
rect 13872 11500 13878 11512
rect 14645 11509 14657 11512
rect 14691 11540 14703 11543
rect 16114 11540 16120 11552
rect 14691 11512 16120 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 17954 11500 17960 11552
rect 18012 11500 18018 11552
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11540 18107 11543
rect 18322 11540 18328 11552
rect 18095 11512 18328 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18800 11540 18828 11571
rect 18966 11568 18972 11620
rect 19024 11568 19030 11620
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19996 11608 20024 11707
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 20272 11753 20300 11784
rect 20622 11772 20628 11824
rect 20680 11772 20686 11824
rect 27522 11772 27528 11824
rect 27580 11812 27586 11824
rect 28353 11815 28411 11821
rect 28353 11812 28365 11815
rect 27580 11784 28365 11812
rect 27580 11772 27586 11784
rect 28353 11781 28365 11784
rect 28399 11781 28411 11815
rect 28353 11775 28411 11781
rect 30285 11815 30343 11821
rect 30285 11781 30297 11815
rect 30331 11812 30343 11815
rect 30374 11812 30380 11824
rect 30331 11784 30380 11812
rect 30331 11781 30343 11784
rect 30285 11775 30343 11781
rect 30374 11772 30380 11784
rect 30432 11812 30438 11824
rect 35161 11815 35219 11821
rect 30432 11784 30696 11812
rect 30432 11772 30438 11784
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 20496 11716 20545 11744
rect 20496 11704 20502 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20714 11704 20720 11756
rect 20772 11704 20778 11756
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 25958 11704 25964 11756
rect 26016 11704 26022 11756
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11744 27491 11747
rect 27982 11744 27988 11756
rect 27479 11716 27988 11744
rect 27479 11713 27491 11716
rect 27433 11707 27491 11713
rect 27982 11704 27988 11716
rect 28040 11704 28046 11756
rect 28629 11747 28687 11753
rect 28629 11713 28641 11747
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 20180 11676 20208 11704
rect 21174 11676 21180 11688
rect 20180 11648 21180 11676
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 25406 11636 25412 11688
rect 25464 11636 25470 11688
rect 26050 11636 26056 11688
rect 26108 11636 26114 11688
rect 26142 11636 26148 11688
rect 26200 11636 26206 11688
rect 27062 11636 27068 11688
rect 27120 11676 27126 11688
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 27120 11648 27629 11676
rect 27120 11636 27126 11648
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 28353 11679 28411 11685
rect 28353 11645 28365 11679
rect 28399 11645 28411 11679
rect 28644 11676 28672 11707
rect 28994 11704 29000 11756
rect 29052 11704 29058 11756
rect 29181 11747 29239 11753
rect 29181 11713 29193 11747
rect 29227 11713 29239 11747
rect 29181 11707 29239 11713
rect 30101 11747 30159 11753
rect 30101 11713 30113 11747
rect 30147 11744 30159 11747
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 30147 11716 30481 11744
rect 30147 11713 30159 11716
rect 30101 11707 30159 11713
rect 30469 11713 30481 11716
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 29089 11679 29147 11685
rect 29089 11676 29101 11679
rect 28644 11648 29101 11676
rect 28353 11639 28411 11645
rect 29089 11645 29101 11648
rect 29135 11645 29147 11679
rect 29196 11676 29224 11707
rect 30006 11676 30012 11688
rect 29196 11648 30012 11676
rect 29089 11639 29147 11645
rect 19392 11580 20024 11608
rect 24780 11608 24808 11636
rect 25593 11611 25651 11617
rect 25593 11608 25605 11611
rect 24780 11580 25605 11608
rect 19392 11568 19398 11580
rect 25593 11577 25605 11580
rect 25639 11577 25651 11611
rect 28368 11608 28396 11639
rect 30006 11636 30012 11648
rect 30064 11636 30070 11688
rect 28810 11608 28816 11620
rect 28368 11580 28816 11608
rect 25593 11571 25651 11577
rect 28810 11568 28816 11580
rect 28868 11608 28874 11620
rect 30116 11608 30144 11707
rect 30558 11704 30564 11756
rect 30616 11704 30622 11756
rect 30668 11753 30696 11784
rect 31312 11784 32352 11812
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11744 30711 11747
rect 31018 11744 31024 11756
rect 30699 11716 31024 11744
rect 30699 11713 30711 11716
rect 30653 11707 30711 11713
rect 31018 11704 31024 11716
rect 31076 11704 31082 11756
rect 31312 11753 31340 11784
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 31312 11676 31340 11707
rect 31478 11704 31484 11756
rect 31536 11704 31542 11756
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11744 31631 11747
rect 31619 11716 31800 11744
rect 31619 11713 31631 11716
rect 31573 11707 31631 11713
rect 31772 11688 31800 11716
rect 31846 11704 31852 11756
rect 31904 11744 31910 11756
rect 32122 11744 32128 11756
rect 31904 11716 32128 11744
rect 31904 11704 31910 11716
rect 32122 11704 32128 11716
rect 32180 11744 32186 11756
rect 32217 11747 32275 11753
rect 32217 11744 32229 11747
rect 32180 11716 32229 11744
rect 32180 11704 32186 11716
rect 32217 11713 32229 11716
rect 32263 11713 32275 11747
rect 32217 11707 32275 11713
rect 28868 11580 30144 11608
rect 30576 11648 31340 11676
rect 28868 11568 28874 11580
rect 19978 11540 19984 11552
rect 18800 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 26970 11500 26976 11552
rect 27028 11540 27034 11552
rect 27246 11540 27252 11552
rect 27028 11512 27252 11540
rect 27028 11500 27034 11512
rect 27246 11500 27252 11512
rect 27304 11500 27310 11552
rect 28534 11500 28540 11552
rect 28592 11500 28598 11552
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 30576 11540 30604 11648
rect 31754 11636 31760 11688
rect 31812 11636 31818 11688
rect 30156 11512 30604 11540
rect 30156 11500 30162 11512
rect 32214 11500 32220 11552
rect 32272 11540 32278 11552
rect 32324 11540 32352 11784
rect 35161 11781 35173 11815
rect 35207 11812 35219 11815
rect 35342 11812 35348 11824
rect 35207 11784 35348 11812
rect 35207 11781 35219 11784
rect 35161 11775 35219 11781
rect 35342 11772 35348 11784
rect 35400 11772 35406 11824
rect 32490 11704 32496 11756
rect 32548 11704 32554 11756
rect 37458 11704 37464 11756
rect 37516 11744 37522 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 37516 11716 37841 11744
rect 37516 11704 37522 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 34422 11568 34428 11620
rect 34480 11608 34486 11620
rect 34977 11611 35035 11617
rect 34977 11608 34989 11611
rect 34480 11580 34989 11608
rect 34480 11568 34486 11580
rect 34977 11577 34989 11580
rect 35023 11608 35035 11611
rect 36998 11608 37004 11620
rect 35023 11580 37004 11608
rect 35023 11577 35035 11580
rect 34977 11571 35035 11577
rect 36998 11568 37004 11580
rect 37056 11568 37062 11620
rect 32401 11543 32459 11549
rect 32401 11540 32413 11543
rect 32272 11512 32413 11540
rect 32272 11500 32278 11512
rect 32401 11509 32413 11512
rect 32447 11509 32459 11543
rect 32401 11503 32459 11509
rect 34698 11500 34704 11552
rect 34756 11540 34762 11552
rect 35618 11540 35624 11552
rect 34756 11512 35624 11540
rect 34756 11500 34762 11512
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 36446 11500 36452 11552
rect 36504 11540 36510 11552
rect 36722 11540 36728 11552
rect 36504 11512 36728 11540
rect 36504 11500 36510 11512
rect 36722 11500 36728 11512
rect 36780 11540 36786 11552
rect 37277 11543 37335 11549
rect 37277 11540 37289 11543
rect 36780 11512 37289 11540
rect 36780 11500 36786 11512
rect 37277 11509 37289 11512
rect 37323 11509 37335 11543
rect 37277 11503 37335 11509
rect 1104 11450 45172 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 45172 11450
rect 1104 11376 45172 11398
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 14642 11336 14648 11348
rect 12216 11308 14648 11336
rect 12216 11296 12222 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 16206 11296 16212 11348
rect 16264 11296 16270 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18969 11339 19027 11345
rect 18969 11336 18981 11339
rect 18012 11308 18981 11336
rect 18012 11296 18018 11308
rect 18969 11305 18981 11308
rect 19015 11305 19027 11339
rect 18969 11299 19027 11305
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 19116 11308 19257 11336
rect 19116 11296 19122 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 22189 11339 22247 11345
rect 19245 11299 19303 11305
rect 19352 11308 19748 11336
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 15930 11268 15936 11280
rect 14516 11240 15936 11268
rect 14516 11228 14522 11240
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 16224 11268 16252 11296
rect 17773 11271 17831 11277
rect 16224 11240 16712 11268
rect 14550 11160 14556 11212
rect 14608 11160 14614 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 15059 11172 16129 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16684 11200 16712 11240
rect 17773 11237 17785 11271
rect 17819 11268 17831 11271
rect 19352 11268 19380 11308
rect 17819 11240 19380 11268
rect 19720 11268 19748 11308
rect 22189 11305 22201 11339
rect 22235 11336 22247 11339
rect 23198 11336 23204 11348
rect 22235 11308 23204 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 24854 11296 24860 11348
rect 24912 11296 24918 11348
rect 25130 11296 25136 11348
rect 25188 11336 25194 11348
rect 26973 11339 27031 11345
rect 26973 11336 26985 11339
rect 25188 11308 26985 11336
rect 25188 11296 25194 11308
rect 26973 11305 26985 11308
rect 27019 11305 27031 11339
rect 26973 11299 27031 11305
rect 27522 11296 27528 11348
rect 27580 11296 27586 11348
rect 28534 11296 28540 11348
rect 28592 11336 28598 11348
rect 28629 11339 28687 11345
rect 28629 11336 28641 11339
rect 28592 11308 28641 11336
rect 28592 11296 28598 11308
rect 28629 11305 28641 11308
rect 28675 11305 28687 11339
rect 28629 11299 28687 11305
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 30098 11336 30104 11348
rect 29052 11308 30104 11336
rect 29052 11296 29058 11308
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 30558 11296 30564 11348
rect 30616 11336 30622 11348
rect 31386 11336 31392 11348
rect 30616 11308 31392 11336
rect 30616 11296 30622 11308
rect 31386 11296 31392 11308
rect 31444 11296 31450 11348
rect 32214 11296 32220 11348
rect 32272 11296 32278 11348
rect 37366 11336 37372 11348
rect 35636 11308 37372 11336
rect 22649 11271 22707 11277
rect 22649 11268 22661 11271
rect 19720 11240 22661 11268
rect 17819 11237 17831 11240
rect 17773 11231 17831 11237
rect 22649 11237 22661 11240
rect 22695 11237 22707 11271
rect 26142 11268 26148 11280
rect 22649 11231 22707 11237
rect 25148 11240 26148 11268
rect 16970 11203 17028 11209
rect 16970 11200 16982 11203
rect 16684 11172 16982 11200
rect 16970 11169 16982 11172
rect 17016 11169 17028 11203
rect 16970 11163 17028 11169
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17310 11200 17316 11212
rect 17175 11172 17316 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 17552 11172 17724 11200
rect 17552 11160 17558 11172
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13412 11104 14473 11132
rect 13412 11092 13418 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 14090 11064 14096 11076
rect 11480 11036 14096 11064
rect 11480 11024 11486 11036
rect 14090 11024 14096 11036
rect 14148 11024 14154 11076
rect 14476 11064 14504 11095
rect 14734 11092 14740 11144
rect 14792 11092 14798 11144
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 15930 11092 15936 11144
rect 15988 11092 15994 11144
rect 16850 11092 16856 11144
rect 16908 11092 16914 11144
rect 17696 11132 17724 11172
rect 18230 11160 18236 11212
rect 18288 11160 18294 11212
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 18555 11172 19717 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 23198 11160 23204 11212
rect 23256 11200 23262 11212
rect 24670 11200 24676 11212
rect 23256 11172 24676 11200
rect 23256 11160 23262 11172
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17696 11104 17877 11132
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18012 11104 18337 11132
rect 18012 11092 18018 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18325 11095 18383 11101
rect 18432 11104 18889 11132
rect 15672 11064 15700 11092
rect 16114 11064 16120 11076
rect 14476 11036 16120 11064
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 17604 11036 18092 11064
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12986 10996 12992 11008
rect 12584 10968 12992 10996
rect 12584 10956 12590 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17218 10996 17224 11008
rect 16632 10968 17224 10996
rect 16632 10956 16638 10968
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17402 10956 17408 11008
rect 17460 10996 17466 11008
rect 17604 10996 17632 11036
rect 17460 10968 17632 10996
rect 17460 10956 17466 10968
rect 17954 10956 17960 11008
rect 18012 10956 18018 11008
rect 18064 11005 18092 11036
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 18432 11064 18460 11104
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19061 11135 19119 11141
rect 19061 11101 19073 11135
rect 19107 11101 19119 11135
rect 19061 11095 19119 11101
rect 18196 11036 18460 11064
rect 18196 11024 18202 11036
rect 18598 11024 18604 11076
rect 18656 11064 18662 11076
rect 19076 11064 19104 11095
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 19392 11104 19441 11132
rect 19392 11092 19398 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19518 11092 19524 11144
rect 19576 11092 19582 11144
rect 19610 11092 19616 11144
rect 19668 11092 19674 11144
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 22646 11132 22652 11144
rect 22511 11104 22652 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 22646 11092 22652 11104
rect 22704 11092 22710 11144
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11132 22799 11135
rect 24486 11132 24492 11144
rect 22787 11104 24492 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 25148 11141 25176 11240
rect 26142 11228 26148 11240
rect 26200 11228 26206 11280
rect 27540 11268 27568 11296
rect 27448 11240 27568 11268
rect 25240 11172 26096 11200
rect 25240 11141 25268 11172
rect 26068 11144 26096 11172
rect 27246 11160 27252 11212
rect 27304 11160 27310 11212
rect 27448 11209 27476 11240
rect 31294 11228 31300 11280
rect 31352 11228 31358 11280
rect 31662 11228 31668 11280
rect 31720 11268 31726 11280
rect 31720 11240 31800 11268
rect 31720 11228 31726 11240
rect 27433 11203 27491 11209
rect 27433 11169 27445 11203
rect 27479 11169 27491 11203
rect 27433 11163 27491 11169
rect 27525 11203 27583 11209
rect 27525 11169 27537 11203
rect 27571 11169 27583 11203
rect 27525 11163 27583 11169
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 25133 11095 25191 11101
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11101 25283 11135
rect 25225 11095 25283 11101
rect 25314 11092 25320 11144
rect 25372 11092 25378 11144
rect 25501 11135 25559 11141
rect 25501 11101 25513 11135
rect 25547 11101 25559 11135
rect 25501 11095 25559 11101
rect 18656 11036 19104 11064
rect 18656 11024 18662 11036
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 19352 11064 19380 11092
rect 19208 11036 19380 11064
rect 19208 11024 19214 11036
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10965 18107 10999
rect 18049 10959 18107 10965
rect 19058 10956 19064 11008
rect 19116 10996 19122 11008
rect 19628 10996 19656 11092
rect 23382 11024 23388 11076
rect 23440 11024 23446 11076
rect 19116 10968 19656 10996
rect 23400 10996 23428 11024
rect 25516 10996 25544 11095
rect 26050 11092 26056 11144
rect 26108 11092 26114 11144
rect 27264 11132 27292 11160
rect 27540 11132 27568 11163
rect 28442 11160 28448 11212
rect 28500 11160 28506 11212
rect 29089 11203 29147 11209
rect 29089 11169 29101 11203
rect 29135 11200 29147 11203
rect 31312 11200 31340 11228
rect 31772 11209 31800 11240
rect 29135 11172 29960 11200
rect 29135 11169 29147 11172
rect 29089 11163 29147 11169
rect 27264 11104 27568 11132
rect 28353 11135 28411 11141
rect 28353 11101 28365 11135
rect 28399 11132 28411 11135
rect 28460 11132 28488 11160
rect 29932 11144 29960 11172
rect 31128 11172 31340 11200
rect 31757 11203 31815 11209
rect 28399 11104 28488 11132
rect 28813 11135 28871 11141
rect 28399 11101 28411 11104
rect 28353 11095 28411 11101
rect 28813 11101 28825 11135
rect 28859 11132 28871 11135
rect 28902 11132 28908 11144
rect 28859 11104 28908 11132
rect 28859 11101 28871 11104
rect 28813 11095 28871 11101
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 29914 11092 29920 11144
rect 29972 11092 29978 11144
rect 30742 11092 30748 11144
rect 30800 11132 30806 11144
rect 31128 11141 31156 11172
rect 31757 11169 31769 11203
rect 31803 11169 31815 11203
rect 31757 11163 31815 11169
rect 31846 11160 31852 11212
rect 31904 11160 31910 11212
rect 32232 11200 32260 11296
rect 35636 11277 35664 11308
rect 37366 11296 37372 11308
rect 37424 11296 37430 11348
rect 35621 11271 35679 11277
rect 35621 11237 35633 11271
rect 35667 11237 35679 11271
rect 35621 11231 35679 11237
rect 38105 11271 38163 11277
rect 38105 11237 38117 11271
rect 38151 11268 38163 11271
rect 38562 11268 38568 11280
rect 38151 11240 38568 11268
rect 38151 11237 38163 11240
rect 38105 11231 38163 11237
rect 38562 11228 38568 11240
rect 38620 11268 38626 11280
rect 38620 11240 38792 11268
rect 38620 11228 38626 11240
rect 32232 11172 32352 11200
rect 30929 11135 30987 11141
rect 30929 11132 30941 11135
rect 30800 11104 30941 11132
rect 30800 11092 30806 11104
rect 30929 11101 30941 11104
rect 30975 11101 30987 11135
rect 30929 11095 30987 11101
rect 31113 11135 31171 11141
rect 31113 11101 31125 11135
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 31294 11092 31300 11144
rect 31352 11092 31358 11144
rect 31386 11092 31392 11144
rect 31444 11092 31450 11144
rect 31666 11135 31724 11141
rect 31666 11110 31678 11135
rect 31588 11101 31678 11110
rect 31712 11101 31724 11135
rect 31588 11095 31724 11101
rect 31941 11135 31999 11141
rect 31941 11101 31953 11135
rect 31987 11101 31999 11135
rect 31941 11095 31999 11101
rect 31588 11082 31708 11095
rect 27341 11067 27399 11073
rect 27341 11033 27353 11067
rect 27387 11064 27399 11067
rect 28258 11064 28264 11076
rect 27387 11036 28264 11064
rect 27387 11033 27399 11036
rect 27341 11027 27399 11033
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 31021 11067 31079 11073
rect 31021 11033 31033 11067
rect 31067 11064 31079 11067
rect 31588 11064 31616 11082
rect 31067 11036 31616 11064
rect 31956 11064 31984 11095
rect 32122 11092 32128 11144
rect 32180 11092 32186 11144
rect 32214 11092 32220 11144
rect 32272 11092 32278 11144
rect 32324 11141 32352 11172
rect 37182 11160 37188 11212
rect 37240 11200 37246 11212
rect 38764 11209 38792 11240
rect 38197 11203 38255 11209
rect 38197 11200 38209 11203
rect 37240 11172 38209 11200
rect 37240 11160 37246 11172
rect 38197 11169 38209 11172
rect 38243 11169 38255 11203
rect 38197 11163 38255 11169
rect 38749 11203 38807 11209
rect 38749 11169 38761 11203
rect 38795 11169 38807 11203
rect 38749 11163 38807 11169
rect 32309 11135 32367 11141
rect 32309 11101 32321 11135
rect 32355 11101 32367 11135
rect 32309 11095 32367 11101
rect 32398 11092 32404 11144
rect 32456 11092 32462 11144
rect 34698 11092 34704 11144
rect 34756 11092 34762 11144
rect 36354 11092 36360 11144
rect 36412 11092 36418 11144
rect 38930 11092 38936 11144
rect 38988 11092 38994 11144
rect 32416 11064 32444 11092
rect 31956 11036 32444 11064
rect 31067 11033 31079 11036
rect 31021 11027 31079 11033
rect 23400 10968 25544 10996
rect 19116 10956 19122 10968
rect 30742 10956 30748 11008
rect 30800 10956 30806 11008
rect 30834 10956 30840 11008
rect 30892 10996 30898 11008
rect 31481 10999 31539 11005
rect 31481 10996 31493 10999
rect 30892 10968 31493 10996
rect 30892 10956 30898 10968
rect 31481 10965 31493 10968
rect 31527 10965 31539 10999
rect 31588 10996 31616 11036
rect 32490 11024 32496 11076
rect 32548 11024 32554 11076
rect 35345 11067 35403 11073
rect 35345 11033 35357 11067
rect 35391 11064 35403 11067
rect 35897 11067 35955 11073
rect 35897 11064 35909 11067
rect 35391 11036 35909 11064
rect 35391 11033 35403 11036
rect 35345 11027 35403 11033
rect 35897 11033 35909 11036
rect 35943 11033 35955 11067
rect 35897 11027 35955 11033
rect 36630 11024 36636 11076
rect 36688 11024 36694 11076
rect 38838 11064 38844 11076
rect 37858 11036 38844 11064
rect 32122 10996 32128 11008
rect 31588 10968 32128 10996
rect 31481 10959 31539 10965
rect 32122 10956 32128 10968
rect 32180 10996 32186 11008
rect 32508 10996 32536 11024
rect 32180 10968 32536 10996
rect 32180 10956 32186 10968
rect 35434 10956 35440 11008
rect 35492 10956 35498 11008
rect 36998 10956 37004 11008
rect 37056 10996 37062 11008
rect 37936 10996 37964 11036
rect 38838 11024 38844 11036
rect 38896 11024 38902 11076
rect 37056 10968 37964 10996
rect 37056 10956 37062 10968
rect 39114 10956 39120 11008
rect 39172 10956 39178 11008
rect 1104 10906 45172 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 45172 10906
rect 1104 10832 45172 10854
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 12710 10752 12716 10804
rect 12768 10752 12774 10804
rect 12820 10764 14872 10792
rect 12544 10724 12572 10752
rect 11624 10696 12020 10724
rect 11624 10668 11652 10696
rect 11606 10616 11612 10668
rect 11664 10616 11670 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11992 10665 12020 10696
rect 12452 10696 12572 10724
rect 12452 10665 12480 10696
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12728 10656 12756 10752
rect 12575 10628 12756 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12342 10588 12348 10600
rect 11756 10560 12348 10588
rect 11756 10548 11762 10560
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 12820 10588 12848 10764
rect 14844 10736 14872 10764
rect 15930 10752 15936 10804
rect 15988 10792 15994 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 15988 10764 16957 10792
rect 15988 10752 15994 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 16945 10755 17003 10761
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 18690 10792 18696 10804
rect 17276 10764 18696 10792
rect 17276 10752 17282 10764
rect 18690 10752 18696 10764
rect 18748 10792 18754 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 18748 10764 19073 10792
rect 18748 10752 18754 10764
rect 19061 10761 19073 10764
rect 19107 10792 19119 10795
rect 19150 10792 19156 10804
rect 19107 10764 19156 10792
rect 19107 10761 19119 10764
rect 19061 10755 19119 10761
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 20530 10792 20536 10804
rect 19392 10764 20536 10792
rect 19392 10752 19398 10764
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 22554 10752 22560 10804
rect 22612 10752 22618 10804
rect 22646 10752 22652 10804
rect 22704 10752 22710 10804
rect 23569 10795 23627 10801
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 24026 10792 24032 10804
rect 23615 10764 24032 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 25314 10752 25320 10804
rect 25372 10752 25378 10804
rect 25593 10795 25651 10801
rect 25593 10761 25605 10795
rect 25639 10792 25651 10795
rect 26050 10792 26056 10804
rect 25639 10764 26056 10792
rect 25639 10761 25651 10764
rect 25593 10755 25651 10761
rect 26050 10752 26056 10764
rect 26108 10752 26114 10804
rect 28905 10795 28963 10801
rect 28905 10792 28917 10795
rect 27172 10764 28917 10792
rect 13280 10696 13584 10724
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12759 10560 12848 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 12912 10520 12940 10619
rect 13078 10548 13084 10600
rect 13136 10588 13142 10600
rect 13280 10588 13308 10696
rect 13354 10616 13360 10668
rect 13412 10616 13418 10668
rect 13556 10665 13584 10696
rect 13630 10684 13636 10736
rect 13688 10724 13694 10736
rect 13688 10696 14044 10724
rect 13688 10684 13694 10696
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 13771 10628 13952 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 13136 10560 13308 10588
rect 13372 10588 13400 10616
rect 13924 10600 13952 10628
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13372 10560 13829 10588
rect 13136 10548 13142 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14016 10597 14044 10696
rect 14826 10684 14832 10736
rect 14884 10684 14890 10736
rect 15470 10684 15476 10736
rect 15528 10724 15534 10736
rect 15746 10724 15752 10736
rect 15528 10696 15752 10724
rect 15528 10684 15534 10696
rect 15746 10684 15752 10696
rect 15804 10724 15810 10736
rect 15804 10696 16620 10724
rect 15804 10684 15810 10696
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 14976 10628 16221 10656
rect 14976 10616 14982 10628
rect 16209 10625 16221 10628
rect 16255 10656 16267 10659
rect 16298 10656 16304 10668
rect 16255 10628 16304 10656
rect 16255 10625 16267 10628
rect 16209 10619 16267 10625
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 16485 10662 16543 10665
rect 16592 10662 16620 10696
rect 17034 10684 17040 10736
rect 17092 10724 17098 10736
rect 22189 10727 22247 10733
rect 22189 10724 22201 10727
rect 17092 10696 22201 10724
rect 17092 10684 17098 10696
rect 22189 10693 22201 10696
rect 22235 10693 22247 10727
rect 22189 10687 22247 10693
rect 23014 10684 23020 10736
rect 23072 10724 23078 10736
rect 23201 10727 23259 10733
rect 23201 10724 23213 10727
rect 23072 10696 23213 10724
rect 23072 10684 23078 10696
rect 23201 10693 23213 10696
rect 23247 10724 23259 10727
rect 23290 10724 23296 10736
rect 23247 10696 23296 10724
rect 23247 10693 23259 10696
rect 23201 10687 23259 10693
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 23750 10684 23756 10736
rect 23808 10724 23814 10736
rect 23845 10727 23903 10733
rect 23845 10724 23857 10727
rect 23808 10696 23857 10724
rect 23808 10684 23814 10696
rect 23845 10693 23857 10696
rect 23891 10693 23903 10727
rect 23845 10687 23903 10693
rect 23934 10687 23940 10736
rect 23933 10684 23940 10687
rect 23992 10684 23998 10736
rect 25332 10724 25360 10752
rect 26973 10727 27031 10733
rect 26973 10724 26985 10727
rect 25332 10696 26985 10724
rect 26973 10693 26985 10696
rect 27019 10693 27031 10727
rect 26973 10687 27031 10693
rect 16485 10659 16620 10662
rect 16485 10625 16497 10659
rect 16531 10634 16620 10659
rect 17129 10659 17187 10665
rect 16531 10625 16543 10634
rect 16485 10619 16543 10625
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10656 17463 10659
rect 17494 10656 17500 10668
rect 17451 10628 17500 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 15194 10588 15200 10600
rect 14047 10560 15200 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16408 10588 16436 10619
rect 15896 10560 16436 10588
rect 15896 10548 15902 10560
rect 13722 10520 13728 10532
rect 12912 10492 13728 10520
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11790 10452 11796 10464
rect 11296 10424 11796 10452
rect 11296 10412 11302 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 12250 10412 12256 10464
rect 12308 10412 12314 10464
rect 13357 10455 13415 10461
rect 13357 10421 13369 10455
rect 13403 10452 13415 10455
rect 13538 10452 13544 10464
rect 13403 10424 13544 10452
rect 13403 10421 13415 10424
rect 13357 10415 13415 10421
rect 13538 10412 13544 10424
rect 13596 10452 13602 10464
rect 13814 10452 13820 10464
rect 13596 10424 13820 10452
rect 13596 10412 13602 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 13909 10455 13967 10461
rect 13909 10421 13921 10455
rect 13955 10452 13967 10455
rect 14550 10452 14556 10464
rect 13955 10424 14556 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 14642 10412 14648 10464
rect 14700 10452 14706 10464
rect 15378 10452 15384 10464
rect 14700 10424 15384 10452
rect 14700 10412 14706 10424
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 16114 10412 16120 10464
rect 16172 10452 16178 10464
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 16172 10424 16221 10452
rect 16172 10412 16178 10424
rect 16209 10421 16221 10424
rect 16255 10421 16267 10455
rect 16209 10415 16267 10421
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16408 10452 16436 10560
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17144 10588 17172 10619
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 19337 10659 19395 10665
rect 19337 10656 19349 10659
rect 19024 10628 19349 10656
rect 19024 10616 19030 10628
rect 19337 10625 19349 10628
rect 19383 10625 19395 10659
rect 19337 10619 19395 10625
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 22462 10656 22468 10668
rect 19613 10619 19671 10625
rect 22020 10628 22468 10656
rect 16632 10560 17172 10588
rect 18892 10588 18920 10616
rect 19628 10588 19656 10619
rect 22020 10597 22048 10628
rect 22462 10616 22468 10628
rect 22520 10656 22526 10668
rect 22925 10659 22983 10665
rect 22520 10628 22692 10656
rect 22520 10616 22526 10628
rect 22664 10597 22692 10628
rect 22925 10625 22937 10659
rect 22971 10625 22983 10659
rect 22925 10619 22983 10625
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10656 23443 10659
rect 23566 10656 23572 10668
rect 23431 10628 23572 10656
rect 23431 10625 23443 10628
rect 23385 10619 23443 10625
rect 18892 10560 19656 10588
rect 22005 10591 22063 10597
rect 16632 10548 16638 10560
rect 19352 10532 19380 10560
rect 22005 10557 22017 10591
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10557 22155 10591
rect 22097 10551 22155 10557
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10557 22707 10591
rect 22940 10588 22968 10619
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 23658 10616 23664 10668
rect 23716 10616 23722 10668
rect 23474 10588 23480 10600
rect 22940 10560 23480 10588
rect 22649 10551 22707 10557
rect 17218 10480 17224 10532
rect 17276 10480 17282 10532
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 18506 10520 18512 10532
rect 17359 10492 18512 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 18506 10480 18512 10492
rect 18564 10520 18570 10532
rect 18874 10520 18880 10532
rect 18564 10492 18880 10520
rect 18564 10480 18570 10492
rect 18874 10480 18880 10492
rect 18932 10480 18938 10532
rect 19334 10480 19340 10532
rect 19392 10480 19398 10532
rect 17954 10452 17960 10464
rect 16356 10424 17960 10452
rect 16356 10412 16362 10424
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19705 10455 19763 10461
rect 19705 10452 19717 10455
rect 19116 10424 19717 10452
rect 19116 10412 19122 10424
rect 19705 10421 19717 10424
rect 19751 10421 19763 10455
rect 22020 10452 22048 10551
rect 22112 10520 22140 10551
rect 23474 10548 23480 10560
rect 23532 10588 23538 10600
rect 23768 10588 23796 10684
rect 23933 10681 23991 10684
rect 23933 10647 23945 10681
rect 23979 10647 23991 10681
rect 27172 10668 27200 10764
rect 28905 10761 28917 10764
rect 28951 10761 28963 10795
rect 28905 10755 28963 10761
rect 29638 10752 29644 10804
rect 29696 10792 29702 10804
rect 29822 10792 29828 10804
rect 29696 10764 29828 10792
rect 29696 10752 29702 10764
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 31018 10752 31024 10804
rect 31076 10752 31082 10804
rect 32493 10795 32551 10801
rect 32493 10792 32505 10795
rect 31128 10764 32505 10792
rect 31128 10724 31156 10764
rect 32493 10761 32505 10764
rect 32539 10761 32551 10795
rect 32493 10755 32551 10761
rect 33597 10795 33655 10801
rect 33597 10761 33609 10795
rect 33643 10792 33655 10795
rect 34698 10792 34704 10804
rect 33643 10764 34704 10792
rect 33643 10761 33655 10764
rect 33597 10755 33655 10761
rect 34698 10752 34704 10764
rect 34756 10752 34762 10804
rect 36630 10752 36636 10804
rect 36688 10792 36694 10804
rect 37001 10795 37059 10801
rect 37001 10792 37013 10795
rect 36688 10764 37013 10792
rect 36688 10752 36694 10764
rect 37001 10761 37013 10764
rect 37047 10761 37059 10795
rect 37001 10755 37059 10761
rect 39114 10752 39120 10804
rect 39172 10792 39178 10804
rect 39172 10764 39896 10792
rect 39172 10752 39178 10764
rect 31570 10724 31576 10736
rect 28184 10696 31156 10724
rect 31220 10696 31576 10724
rect 23933 10641 23991 10647
rect 25961 10659 26019 10665
rect 25961 10625 25973 10659
rect 26007 10656 26019 10659
rect 26786 10656 26792 10668
rect 26007 10628 26792 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 26786 10616 26792 10628
rect 26844 10616 26850 10668
rect 27062 10616 27068 10668
rect 27120 10616 27126 10668
rect 27154 10616 27160 10668
rect 27212 10616 27218 10668
rect 27522 10665 27528 10668
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10625 27307 10659
rect 27249 10619 27307 10625
rect 27418 10659 27476 10665
rect 27418 10625 27430 10659
rect 27464 10625 27476 10659
rect 27418 10619 27476 10625
rect 27515 10659 27528 10665
rect 27515 10625 27527 10659
rect 27580 10656 27586 10668
rect 27580 10628 27615 10656
rect 27515 10619 27528 10625
rect 23532 10560 23796 10588
rect 26053 10591 26111 10597
rect 23532 10548 23538 10560
rect 26053 10557 26065 10591
rect 26099 10557 26111 10591
rect 26053 10551 26111 10557
rect 23661 10523 23719 10529
rect 23661 10520 23673 10523
rect 22112 10492 23673 10520
rect 23661 10489 23673 10492
rect 23707 10489 23719 10523
rect 23661 10483 23719 10489
rect 25406 10480 25412 10532
rect 25464 10480 25470 10532
rect 26068 10520 26096 10551
rect 26234 10548 26240 10600
rect 26292 10548 26298 10600
rect 27080 10588 27108 10616
rect 27264 10588 27292 10619
rect 27080 10560 27292 10588
rect 27448 10588 27476 10619
rect 27522 10616 27528 10619
rect 27580 10616 27586 10628
rect 28074 10588 28080 10600
rect 27448 10560 28080 10588
rect 28074 10548 28080 10560
rect 28132 10548 28138 10600
rect 26510 10520 26516 10532
rect 26068 10492 26516 10520
rect 26510 10480 26516 10492
rect 26568 10520 26574 10532
rect 28184 10520 28212 10696
rect 28258 10616 28264 10668
rect 28316 10656 28322 10668
rect 28353 10659 28411 10665
rect 28353 10656 28365 10659
rect 28316 10628 28365 10656
rect 28316 10616 28322 10628
rect 28353 10625 28365 10628
rect 28399 10625 28411 10659
rect 28353 10619 28411 10625
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 29086 10616 29092 10668
rect 29144 10656 29150 10668
rect 29457 10659 29515 10665
rect 29457 10656 29469 10659
rect 29144 10628 29469 10656
rect 29144 10616 29150 10628
rect 29457 10625 29469 10628
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 29549 10659 29607 10665
rect 29549 10625 29561 10659
rect 29595 10656 29607 10659
rect 29638 10656 29644 10668
rect 29595 10628 29644 10656
rect 29595 10625 29607 10628
rect 29549 10619 29607 10625
rect 29638 10616 29644 10628
rect 29696 10616 29702 10668
rect 29733 10659 29791 10665
rect 29733 10625 29745 10659
rect 29779 10656 29791 10659
rect 29914 10656 29920 10668
rect 29779 10628 29920 10656
rect 29779 10625 29791 10628
rect 29733 10619 29791 10625
rect 29914 10616 29920 10628
rect 29972 10616 29978 10668
rect 30006 10616 30012 10668
rect 30064 10616 30070 10668
rect 30098 10616 30104 10668
rect 30156 10656 30162 10668
rect 31220 10665 31248 10696
rect 31570 10684 31576 10696
rect 31628 10684 31634 10736
rect 31662 10684 31668 10736
rect 31720 10684 31726 10736
rect 31846 10684 31852 10736
rect 31904 10724 31910 10736
rect 31904 10696 32260 10724
rect 31904 10684 31910 10696
rect 30193 10659 30251 10665
rect 30193 10656 30205 10659
rect 30156 10628 30205 10656
rect 30156 10616 30162 10628
rect 30193 10625 30205 10628
rect 30239 10625 30251 10659
rect 30193 10619 30251 10625
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10625 31079 10659
rect 31021 10619 31079 10625
rect 31205 10659 31263 10665
rect 31205 10625 31217 10659
rect 31251 10625 31263 10659
rect 31205 10619 31263 10625
rect 28537 10591 28595 10597
rect 28537 10557 28549 10591
rect 28583 10557 28595 10591
rect 28537 10551 28595 10557
rect 26568 10492 28212 10520
rect 28552 10520 28580 10551
rect 29178 10548 29184 10600
rect 29236 10548 29242 10600
rect 28994 10520 29000 10532
rect 28552 10492 29000 10520
rect 26568 10480 26574 10492
rect 28994 10480 29000 10492
rect 29052 10520 29058 10532
rect 29549 10523 29607 10529
rect 29549 10520 29561 10523
rect 29052 10492 29561 10520
rect 29052 10480 29058 10492
rect 29549 10489 29561 10492
rect 29595 10489 29607 10523
rect 29549 10483 29607 10489
rect 29748 10492 30880 10520
rect 22094 10452 22100 10464
rect 22020 10424 22100 10452
rect 19705 10415 19763 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22830 10412 22836 10464
rect 22888 10412 22894 10464
rect 25424 10452 25452 10480
rect 27522 10452 27528 10464
rect 25424 10424 27528 10452
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 28166 10412 28172 10464
rect 28224 10412 28230 10464
rect 28721 10455 28779 10461
rect 28721 10421 28733 10455
rect 28767 10452 28779 10455
rect 29270 10452 29276 10464
rect 28767 10424 29276 10452
rect 28767 10421 28779 10424
rect 28721 10415 28779 10421
rect 29270 10412 29276 10424
rect 29328 10412 29334 10464
rect 29365 10455 29423 10461
rect 29365 10421 29377 10455
rect 29411 10452 29423 10455
rect 29748 10452 29776 10492
rect 30852 10464 30880 10492
rect 29411 10424 29776 10452
rect 29411 10421 29423 10424
rect 29365 10415 29423 10421
rect 29822 10412 29828 10464
rect 29880 10452 29886 10464
rect 29917 10455 29975 10461
rect 29917 10452 29929 10455
rect 29880 10424 29929 10452
rect 29880 10412 29886 10424
rect 29917 10421 29929 10424
rect 29963 10421 29975 10455
rect 29917 10415 29975 10421
rect 30834 10412 30840 10464
rect 30892 10412 30898 10464
rect 31036 10452 31064 10619
rect 31386 10616 31392 10668
rect 31444 10656 31450 10668
rect 31481 10659 31539 10665
rect 31481 10656 31493 10659
rect 31444 10628 31493 10656
rect 31444 10616 31450 10628
rect 31481 10625 31493 10628
rect 31527 10656 31539 10659
rect 31680 10656 31708 10684
rect 31527 10628 31708 10656
rect 31527 10625 31539 10628
rect 31481 10619 31539 10625
rect 32030 10616 32036 10668
rect 32088 10616 32094 10668
rect 32232 10665 32260 10696
rect 34422 10684 34428 10736
rect 34480 10684 34486 10736
rect 35069 10727 35127 10733
rect 35069 10693 35081 10727
rect 35115 10724 35127 10727
rect 36446 10724 36452 10736
rect 35115 10696 36452 10724
rect 35115 10693 35127 10696
rect 35069 10687 35127 10693
rect 36446 10684 36452 10696
rect 36504 10684 36510 10736
rect 39868 10733 39896 10764
rect 39853 10727 39911 10733
rect 39853 10693 39865 10727
rect 39899 10693 39911 10727
rect 39853 10687 39911 10693
rect 32125 10659 32183 10665
rect 32125 10625 32137 10659
rect 32171 10625 32183 10659
rect 32125 10619 32183 10625
rect 32217 10659 32275 10665
rect 32217 10625 32229 10659
rect 32263 10625 32275 10659
rect 32217 10619 32275 10625
rect 36909 10659 36967 10665
rect 36909 10625 36921 10659
rect 36955 10625 36967 10659
rect 36909 10619 36967 10625
rect 37093 10659 37151 10665
rect 37093 10625 37105 10659
rect 37139 10656 37151 10659
rect 37366 10656 37372 10668
rect 37139 10628 37372 10656
rect 37139 10625 37151 10628
rect 37093 10619 37151 10625
rect 31941 10591 31999 10597
rect 31941 10557 31953 10591
rect 31987 10588 31999 10591
rect 32048 10588 32076 10616
rect 31987 10560 32076 10588
rect 31987 10557 31999 10560
rect 31941 10551 31999 10557
rect 31478 10480 31484 10532
rect 31536 10520 31542 10532
rect 32140 10520 32168 10619
rect 35345 10591 35403 10597
rect 35345 10557 35357 10591
rect 35391 10557 35403 10591
rect 36924 10588 36952 10619
rect 37366 10616 37372 10628
rect 37424 10616 37430 10668
rect 38838 10656 38844 10668
rect 38778 10628 38844 10656
rect 38838 10616 38844 10628
rect 38896 10616 38902 10668
rect 40129 10659 40187 10665
rect 40129 10625 40141 10659
rect 40175 10656 40187 10659
rect 40678 10656 40684 10668
rect 40175 10628 40684 10656
rect 40175 10625 40187 10628
rect 40129 10619 40187 10625
rect 40678 10616 40684 10628
rect 40736 10616 40742 10668
rect 37277 10591 37335 10597
rect 37277 10588 37289 10591
rect 36924 10560 37289 10588
rect 35345 10551 35403 10557
rect 37277 10557 37289 10560
rect 37323 10557 37335 10591
rect 37277 10551 37335 10557
rect 31536 10492 32168 10520
rect 31536 10480 31542 10492
rect 35360 10464 35388 10551
rect 37826 10548 37832 10600
rect 37884 10548 37890 10600
rect 40218 10548 40224 10600
rect 40276 10588 40282 10600
rect 40497 10591 40555 10597
rect 40497 10588 40509 10591
rect 40276 10560 40509 10588
rect 40276 10548 40282 10560
rect 40497 10557 40509 10560
rect 40543 10557 40555 10591
rect 40497 10551 40555 10557
rect 31662 10452 31668 10464
rect 31036 10424 31668 10452
rect 31662 10412 31668 10424
rect 31720 10412 31726 10464
rect 32214 10412 32220 10464
rect 32272 10412 32278 10464
rect 34698 10412 34704 10464
rect 34756 10452 34762 10464
rect 35342 10452 35348 10464
rect 34756 10424 35348 10452
rect 34756 10412 34762 10424
rect 35342 10412 35348 10424
rect 35400 10412 35406 10464
rect 38378 10412 38384 10464
rect 38436 10412 38442 10464
rect 41141 10455 41199 10461
rect 41141 10421 41153 10455
rect 41187 10452 41199 10455
rect 41230 10452 41236 10464
rect 41187 10424 41236 10452
rect 41187 10421 41199 10424
rect 41141 10415 41199 10421
rect 41230 10412 41236 10424
rect 41288 10412 41294 10464
rect 1104 10362 45172 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 45172 10362
rect 1104 10288 45172 10310
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 12250 10208 12256 10260
rect 12308 10208 12314 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12400 10220 12572 10248
rect 12400 10208 12406 10220
rect 12158 10140 12164 10192
rect 12216 10140 12222 10192
rect 12268 10180 12296 10208
rect 12544 10180 12572 10220
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 12676 10220 13553 10248
rect 12676 10208 12682 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 14921 10251 14979 10257
rect 13955 10220 14872 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 14553 10183 14611 10189
rect 14553 10180 14565 10183
rect 12268 10152 12434 10180
rect 12544 10152 14565 10180
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11572 10084 11713 10112
rect 11572 10072 11578 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 12176 10112 12204 10140
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 12176 10084 12265 10112
rect 11701 10075 11759 10081
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12406 10112 12434 10152
rect 14553 10149 14565 10152
rect 14599 10149 14611 10183
rect 14844 10180 14872 10220
rect 14921 10217 14933 10251
rect 14967 10248 14979 10251
rect 15562 10248 15568 10260
rect 14967 10220 15568 10248
rect 14967 10217 14979 10220
rect 14921 10211 14979 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16850 10248 16856 10260
rect 16531 10220 16856 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19116 10220 19656 10248
rect 19116 10208 19122 10220
rect 19426 10180 19432 10192
rect 14844 10152 19432 10180
rect 14553 10143 14611 10149
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12406 10084 12725 10112
rect 12253 10075 12311 10081
rect 12713 10081 12725 10084
rect 12759 10081 12771 10115
rect 12713 10075 12771 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 14182 10112 14188 10124
rect 13136 10084 14188 10112
rect 13136 10072 13142 10084
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14240 10084 14473 10112
rect 14240 10072 14246 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14568 10112 14596 10143
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 14568 10084 15976 10112
rect 14461 10075 14519 10081
rect 11882 10053 11888 10056
rect 11860 10047 11888 10053
rect 11860 10013 11872 10047
rect 11860 10007 11888 10013
rect 11882 10004 11888 10007
rect 11940 10004 11946 10056
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 12894 10004 12900 10056
rect 12952 10004 12958 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14274 10044 14280 10056
rect 13771 10016 14280 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 13556 9976 13584 10007
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14476 10044 14504 10075
rect 14642 10044 14648 10056
rect 14476 10016 14648 10044
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 14752 9976 14780 10007
rect 12820 9948 13584 9976
rect 14568 9948 14780 9976
rect 15948 9976 15976 10084
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 16666 10112 16672 10124
rect 16172 10084 16528 10112
rect 16172 10072 16178 10084
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 16500 10053 16528 10084
rect 16592 10084 16672 10112
rect 16592 10053 16620 10084
rect 16666 10072 16672 10084
rect 16724 10112 16730 10124
rect 16850 10112 16856 10124
rect 16724 10084 16856 10112
rect 16724 10072 16730 10084
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 19628 10112 19656 10220
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20128 10220 20668 10248
rect 20128 10208 20134 10220
rect 19978 10140 19984 10192
rect 20036 10140 20042 10192
rect 19996 10112 20024 10140
rect 20088 10121 20116 10208
rect 20346 10180 20352 10192
rect 20272 10152 20352 10180
rect 17920 10084 19564 10112
rect 17920 10072 17926 10084
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 16942 10044 16948 10056
rect 16807 10016 16948 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 16776 9976 16804 10007
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 19536 10053 19564 10084
rect 19628 10084 20024 10112
rect 20073 10115 20131 10121
rect 19628 10053 19656 10084
rect 20073 10081 20085 10115
rect 20119 10081 20131 10115
rect 20073 10075 20131 10081
rect 20272 10053 20300 10152
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 20640 10112 20668 10220
rect 22738 10208 22744 10260
rect 22796 10208 22802 10260
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 22888 10220 25697 10248
rect 22888 10208 22894 10220
rect 25685 10217 25697 10220
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 26786 10208 26792 10260
rect 26844 10248 26850 10260
rect 26844 10220 27568 10248
rect 26844 10208 26850 10220
rect 22756 10180 22784 10208
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 22756 10152 24501 10180
rect 24489 10149 24501 10152
rect 24535 10149 24547 10183
rect 25406 10180 25412 10192
rect 24489 10143 24547 10149
rect 25056 10152 25412 10180
rect 20579 10084 20668 10112
rect 20993 10115 21051 10121
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 20993 10081 21005 10115
rect 21039 10112 21051 10115
rect 23842 10112 23848 10124
rect 21039 10084 23848 10112
rect 21039 10081 21051 10084
rect 20993 10075 21051 10081
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 25056 10121 25084 10152
rect 25406 10140 25412 10152
rect 25464 10180 25470 10192
rect 27154 10180 27160 10192
rect 25464 10152 25820 10180
rect 25464 10140 25470 10152
rect 25792 10124 25820 10152
rect 26804 10152 27160 10180
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10081 25099 10115
rect 25041 10075 25099 10081
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 25774 10072 25780 10124
rect 25832 10072 25838 10124
rect 26142 10072 26148 10124
rect 26200 10112 26206 10124
rect 26510 10121 26516 10124
rect 26329 10115 26387 10121
rect 26329 10112 26341 10115
rect 26200 10084 26341 10112
rect 26200 10072 26206 10084
rect 26329 10081 26341 10084
rect 26375 10081 26387 10115
rect 26329 10075 26387 10081
rect 26488 10115 26516 10121
rect 26488 10081 26500 10115
rect 26488 10075 26516 10081
rect 26510 10072 26516 10075
rect 26568 10072 26574 10124
rect 26605 10115 26663 10121
rect 26605 10081 26617 10115
rect 26651 10112 26663 10115
rect 26804 10112 26832 10152
rect 27154 10140 27160 10152
rect 27212 10140 27218 10192
rect 27540 10180 27568 10220
rect 27982 10208 27988 10260
rect 28040 10248 28046 10260
rect 28629 10251 28687 10257
rect 28629 10248 28641 10251
rect 28040 10220 28641 10248
rect 28040 10208 28046 10220
rect 28629 10217 28641 10220
rect 28675 10217 28687 10251
rect 28629 10211 28687 10217
rect 28994 10208 29000 10260
rect 29052 10208 29058 10260
rect 29178 10208 29184 10260
rect 29236 10208 29242 10260
rect 29270 10208 29276 10260
rect 29328 10248 29334 10260
rect 31113 10251 31171 10257
rect 31113 10248 31125 10251
rect 29328 10220 31125 10248
rect 29328 10208 29334 10220
rect 31113 10217 31125 10220
rect 31159 10248 31171 10251
rect 31294 10248 31300 10260
rect 31159 10220 31300 10248
rect 31159 10217 31171 10220
rect 31113 10211 31171 10217
rect 31294 10208 31300 10220
rect 31352 10208 31358 10260
rect 31386 10208 31392 10260
rect 31444 10208 31450 10260
rect 31570 10208 31576 10260
rect 31628 10208 31634 10260
rect 35342 10208 35348 10260
rect 35400 10248 35406 10260
rect 36354 10248 36360 10260
rect 35400 10220 36360 10248
rect 35400 10208 35406 10220
rect 36354 10208 36360 10220
rect 36412 10248 36418 10260
rect 36725 10251 36783 10257
rect 36725 10248 36737 10251
rect 36412 10220 36737 10248
rect 36412 10208 36418 10220
rect 36725 10217 36737 10220
rect 36771 10217 36783 10251
rect 36725 10211 36783 10217
rect 39577 10251 39635 10257
rect 39577 10217 39589 10251
rect 39623 10248 39635 10251
rect 40218 10248 40224 10260
rect 39623 10220 40224 10248
rect 39623 10217 39635 10220
rect 39577 10211 39635 10217
rect 30742 10180 30748 10192
rect 27540 10152 30748 10180
rect 26651 10084 26832 10112
rect 26881 10115 26939 10121
rect 26651 10081 26663 10084
rect 26605 10075 26663 10081
rect 26881 10081 26893 10115
rect 26927 10112 26939 10115
rect 27246 10112 27252 10124
rect 26927 10084 27252 10112
rect 26927 10081 26939 10084
rect 26881 10075 26939 10081
rect 27246 10072 27252 10084
rect 27304 10072 27310 10124
rect 27540 10121 27568 10152
rect 30742 10140 30748 10152
rect 30800 10140 30806 10192
rect 31202 10140 31208 10192
rect 31260 10140 31266 10192
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10081 27583 10115
rect 31220 10112 31248 10140
rect 27525 10075 27583 10081
rect 29196 10084 31248 10112
rect 31404 10112 31432 10208
rect 35434 10180 35440 10192
rect 34164 10152 35440 10180
rect 31404 10084 31616 10112
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 18104 10016 19257 10044
rect 18104 10004 18110 10016
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10013 19671 10047
rect 19987 10047 20045 10053
rect 19987 10046 19999 10047
rect 19613 10007 19671 10013
rect 19904 10018 19999 10046
rect 19444 9976 19472 10007
rect 19904 9976 19932 10018
rect 19987 10013 19999 10018
rect 20033 10013 20045 10047
rect 20165 10047 20223 10053
rect 20165 10042 20177 10047
rect 19987 10007 20045 10013
rect 20088 10014 20177 10042
rect 15948 9948 16804 9976
rect 18984 9948 19472 9976
rect 19628 9948 19932 9976
rect 12820 9920 12848 9948
rect 14568 9920 14596 9948
rect 18984 9920 19012 9948
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12526 9908 12532 9920
rect 12308 9880 12532 9908
rect 12308 9868 12314 9880
rect 12526 9868 12532 9880
rect 12584 9908 12590 9920
rect 12710 9908 12716 9920
rect 12584 9880 12716 9908
rect 12584 9868 12590 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12802 9868 12808 9920
rect 12860 9868 12866 9920
rect 14550 9868 14556 9920
rect 14608 9868 14614 9920
rect 16301 9911 16359 9917
rect 16301 9877 16313 9911
rect 16347 9908 16359 9911
rect 16666 9908 16672 9920
rect 16347 9880 16672 9908
rect 16347 9877 16359 9880
rect 16301 9871 16359 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 18966 9868 18972 9920
rect 19024 9868 19030 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19628 9908 19656 9948
rect 19208 9880 19656 9908
rect 19889 9911 19947 9917
rect 19208 9868 19214 9880
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 19978 9908 19984 9920
rect 19935 9880 19984 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20088 9908 20116 10014
rect 20165 10013 20177 10014
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10041 20315 10047
rect 20346 10041 20352 10056
rect 20303 10013 20352 10041
rect 20257 10007 20315 10013
rect 20346 10004 20352 10013
rect 20404 10004 20410 10056
rect 20438 10006 20444 10058
rect 20496 10006 20502 10058
rect 20625 10047 20683 10053
rect 20625 10013 20637 10047
rect 20671 10044 20683 10047
rect 20714 10044 20720 10056
rect 20671 10016 20720 10044
rect 20671 10013 20683 10016
rect 20625 10007 20683 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 20806 10004 20812 10056
rect 20864 10004 20870 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25148 10044 25176 10072
rect 24995 10016 25176 10044
rect 27341 10047 27399 10053
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 27341 10013 27353 10047
rect 27387 10044 27399 10047
rect 27430 10044 27436 10056
rect 27387 10016 27436 10044
rect 27387 10013 27399 10016
rect 27341 10007 27399 10013
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10013 28871 10047
rect 28813 10007 28871 10013
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10044 29055 10047
rect 29196 10044 29224 10084
rect 29043 10016 29224 10044
rect 29273 10047 29331 10053
rect 29043 10013 29055 10016
rect 28997 10007 29055 10013
rect 29273 10013 29285 10047
rect 29319 10044 29331 10047
rect 29319 10016 29684 10044
rect 29319 10013 29331 10016
rect 29273 10007 29331 10013
rect 22554 9936 22560 9988
rect 22612 9976 22618 9988
rect 28828 9976 28856 10007
rect 29178 9976 29184 9988
rect 22612 9948 25728 9976
rect 28828 9948 29184 9976
rect 22612 9936 22618 9948
rect 20530 9908 20536 9920
rect 20088 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9908 20594 9920
rect 20990 9908 20996 9920
rect 20588 9880 20996 9908
rect 20588 9868 20594 9880
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 22244 9880 22293 9908
rect 22244 9868 22250 9880
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 22281 9871 22339 9877
rect 24857 9911 24915 9917
rect 24857 9877 24869 9911
rect 24903 9908 24915 9911
rect 25590 9908 25596 9920
rect 24903 9880 25596 9908
rect 24903 9877 24915 9880
rect 24857 9871 24915 9877
rect 25590 9868 25596 9880
rect 25648 9868 25654 9920
rect 25700 9908 25728 9948
rect 29178 9936 29184 9948
rect 29236 9936 29242 9988
rect 29454 9936 29460 9988
rect 29512 9936 29518 9988
rect 29472 9908 29500 9936
rect 29656 9920 29684 10016
rect 30006 10004 30012 10056
rect 30064 10044 30070 10056
rect 30929 10047 30987 10053
rect 30929 10044 30941 10047
rect 30064 10016 30941 10044
rect 30064 10004 30070 10016
rect 30929 10013 30941 10016
rect 30975 10013 30987 10047
rect 30929 10007 30987 10013
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10044 31171 10047
rect 31294 10044 31300 10056
rect 31159 10016 31300 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 30944 9976 30972 10007
rect 31294 10004 31300 10016
rect 31352 10004 31358 10056
rect 31404 9976 31432 10084
rect 31481 10047 31539 10053
rect 31481 10013 31493 10047
rect 31527 10013 31539 10047
rect 31588 10044 31616 10084
rect 31656 10047 31714 10053
rect 31656 10044 31668 10047
rect 31588 10016 31668 10044
rect 31481 10007 31539 10013
rect 31656 10013 31668 10016
rect 31702 10013 31714 10047
rect 31656 10007 31714 10013
rect 30944 9948 31432 9976
rect 31496 9976 31524 10007
rect 31754 10004 31760 10056
rect 31812 10004 31818 10056
rect 31941 10047 31999 10053
rect 31941 10013 31953 10047
rect 31987 10044 31999 10047
rect 32122 10044 32128 10056
rect 31987 10016 32128 10044
rect 31987 10013 31999 10016
rect 31941 10007 31999 10013
rect 31956 9976 31984 10007
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 34164 10053 34192 10152
rect 35434 10140 35440 10152
rect 35492 10140 35498 10192
rect 34606 10072 34612 10124
rect 34664 10072 34670 10124
rect 36740 10112 36768 10211
rect 40218 10208 40224 10220
rect 40276 10208 40282 10260
rect 37277 10115 37335 10121
rect 37277 10112 37289 10115
rect 36740 10084 37289 10112
rect 37277 10081 37289 10084
rect 37323 10081 37335 10115
rect 37277 10075 37335 10081
rect 39206 10072 39212 10124
rect 39264 10072 39270 10124
rect 41230 10072 41236 10124
rect 41288 10112 41294 10124
rect 41325 10115 41383 10121
rect 41325 10112 41337 10115
rect 41288 10084 41337 10112
rect 41288 10072 41294 10084
rect 41325 10081 41337 10084
rect 41371 10081 41383 10115
rect 41325 10075 41383 10081
rect 41601 10115 41659 10121
rect 41601 10081 41613 10115
rect 41647 10112 41659 10115
rect 43441 10115 43499 10121
rect 43441 10112 43453 10115
rect 41647 10084 43453 10112
rect 41647 10081 41659 10084
rect 41601 10075 41659 10081
rect 43441 10081 43453 10084
rect 43487 10112 43499 10115
rect 43622 10112 43628 10124
rect 43487 10084 43628 10112
rect 43487 10081 43499 10084
rect 43441 10075 43499 10081
rect 43622 10072 43628 10084
rect 43680 10072 43686 10124
rect 34149 10047 34207 10053
rect 34149 10013 34161 10047
rect 34195 10013 34207 10047
rect 34149 10007 34207 10013
rect 34425 10047 34483 10053
rect 34425 10013 34437 10047
rect 34471 10044 34483 10047
rect 34624 10044 34652 10072
rect 34471 10016 34652 10044
rect 34471 10013 34483 10016
rect 34425 10007 34483 10013
rect 39298 10004 39304 10056
rect 39356 10004 39362 10056
rect 31496 9948 31984 9976
rect 35437 9979 35495 9985
rect 35437 9945 35449 9979
rect 35483 9976 35495 9979
rect 37274 9976 37280 9988
rect 35483 9948 37280 9976
rect 35483 9945 35495 9948
rect 35437 9939 35495 9945
rect 37274 9936 37280 9948
rect 37332 9936 37338 9988
rect 37550 9936 37556 9988
rect 37608 9936 37614 9988
rect 38838 9976 38844 9988
rect 38778 9948 38844 9976
rect 38838 9936 38844 9948
rect 38896 9976 38902 9988
rect 38896 9948 39988 9976
rect 38896 9936 38902 9948
rect 25700 9880 29500 9908
rect 29638 9868 29644 9920
rect 29696 9868 29702 9920
rect 31294 9868 31300 9920
rect 31352 9908 31358 9920
rect 31662 9908 31668 9920
rect 31352 9880 31668 9908
rect 31352 9868 31358 9880
rect 31662 9868 31668 9880
rect 31720 9908 31726 9920
rect 31757 9911 31815 9917
rect 31757 9908 31769 9911
rect 31720 9880 31769 9908
rect 31720 9868 31726 9880
rect 31757 9877 31769 9880
rect 31803 9877 31815 9911
rect 31757 9871 31815 9877
rect 33962 9868 33968 9920
rect 34020 9868 34026 9920
rect 34238 9868 34244 9920
rect 34296 9868 34302 9920
rect 39022 9868 39028 9920
rect 39080 9868 39086 9920
rect 39850 9868 39856 9920
rect 39908 9868 39914 9920
rect 39960 9908 39988 9948
rect 40862 9936 40868 9988
rect 40920 9976 40926 9988
rect 40920 9948 41998 9976
rect 40920 9936 40926 9948
rect 40972 9908 41000 9948
rect 43162 9936 43168 9988
rect 43220 9936 43226 9988
rect 39960 9880 41000 9908
rect 41690 9868 41696 9920
rect 41748 9908 41754 9920
rect 42150 9908 42156 9920
rect 41748 9880 42156 9908
rect 41748 9868 41754 9880
rect 42150 9868 42156 9880
rect 42208 9868 42214 9920
rect 1104 9818 45172 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 45172 9818
rect 1104 9744 45172 9766
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12032 9676 12204 9704
rect 12032 9664 12038 9676
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 11164 9500 11192 9531
rect 11238 9500 11244 9512
rect 11164 9472 11244 9500
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11348 9500 11376 9531
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12176 9577 12204 9676
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 16206 9704 16212 9716
rect 16080 9676 16212 9704
rect 16080 9664 16086 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 19610 9704 19616 9716
rect 16356 9676 16896 9704
rect 16356 9664 16362 9676
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9605 12311 9639
rect 12253 9599 12311 9605
rect 12529 9639 12587 9645
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 14642 9636 14648 9648
rect 12575 9608 13032 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12268 9568 12296 9599
rect 13004 9580 13032 9608
rect 13096 9608 14648 9636
rect 12342 9568 12348 9580
rect 12268 9540 12348 9568
rect 12161 9531 12219 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12657 9571 12715 9577
rect 12657 9537 12669 9571
rect 12703 9568 12715 9571
rect 12802 9568 12808 9580
rect 12703 9540 12808 9568
rect 12703 9537 12715 9540
rect 12657 9531 12715 9537
rect 12452 9500 12480 9531
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12986 9528 12992 9580
rect 13044 9528 13050 9580
rect 13096 9577 13124 9608
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 15286 9636 15292 9648
rect 14844 9608 15292 9636
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 11348 9472 11468 9500
rect 11440 9444 11468 9472
rect 11716 9472 12480 9500
rect 12529 9503 12587 9509
rect 11422 9392 11428 9444
rect 11480 9392 11486 9444
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9364 11299 9367
rect 11716 9364 11744 9472
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12894 9500 12900 9512
rect 12575 9472 12900 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 13096 9432 13124 9531
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13538 9568 13544 9580
rect 13495 9540 13544 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13832 9540 14289 9568
rect 13832 9512 13860 9540
rect 14277 9537 14289 9540
rect 14323 9568 14335 9571
rect 14550 9568 14556 9580
rect 14323 9540 14556 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14844 9577 14872 9608
rect 15286 9596 15292 9608
rect 15344 9636 15350 9648
rect 15344 9608 16160 9636
rect 15344 9596 15350 9608
rect 16132 9577 16160 9608
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 14829 9531 14887 9537
rect 15396 9540 15945 9568
rect 13814 9460 13820 9512
rect 13872 9460 13878 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14366 9500 14372 9512
rect 13964 9472 14372 9500
rect 13964 9460 13970 9472
rect 14366 9460 14372 9472
rect 14424 9500 14430 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14424 9472 14473 9500
rect 14424 9460 14430 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 15396 9432 15424 9540
rect 15933 9537 15945 9540
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16206 9568 16212 9580
rect 16163 9540 16212 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 15948 9500 15976 9531
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16666 9528 16672 9580
rect 16724 9528 16730 9580
rect 16868 9577 16896 9676
rect 19536 9676 19616 9704
rect 18966 9636 18972 9648
rect 17144 9608 17632 9636
rect 17144 9577 17172 9608
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17218 9528 17224 9580
rect 17276 9528 17282 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17359 9540 17540 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 16574 9500 16580 9512
rect 15948 9472 16580 9500
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16684 9500 16712 9528
rect 16684 9472 17448 9500
rect 17420 9444 17448 9472
rect 11848 9404 13124 9432
rect 14016 9404 15424 9432
rect 11848 9392 11854 9404
rect 14016 9376 14044 9404
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 16448 9404 17359 9432
rect 16448 9392 16454 9404
rect 11287 9336 11744 9364
rect 11287 9333 11299 9336
rect 11241 9327 11299 9333
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 13998 9364 14004 9376
rect 12032 9336 14004 9364
rect 12032 9324 12038 9336
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14090 9324 14096 9376
rect 14148 9324 14154 9376
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 14826 9364 14832 9376
rect 14691 9336 14832 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 14826 9324 14832 9336
rect 14884 9364 14890 9376
rect 16574 9364 16580 9376
rect 14884 9336 16580 9364
rect 14884 9324 14890 9336
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16761 9367 16819 9373
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 16850 9364 16856 9376
rect 16807 9336 16856 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17331 9364 17359 9404
rect 17402 9392 17408 9444
rect 17460 9392 17466 9444
rect 17512 9364 17540 9540
rect 17604 9376 17632 9608
rect 18524 9608 18972 9636
rect 18524 9580 18552 9608
rect 18966 9596 18972 9608
rect 19024 9596 19030 9648
rect 19429 9639 19487 9645
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 19536 9636 19564 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 20530 9704 20536 9716
rect 19852 9676 20536 9704
rect 19852 9664 19858 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 22649 9707 22707 9713
rect 22649 9673 22661 9707
rect 22695 9704 22707 9707
rect 23474 9704 23480 9716
rect 22695 9676 23480 9704
rect 22695 9673 22707 9676
rect 22649 9667 22707 9673
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23716 9676 23857 9704
rect 23716 9664 23722 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 26145 9707 26203 9713
rect 26145 9673 26157 9707
rect 26191 9704 26203 9707
rect 26786 9704 26792 9716
rect 26191 9676 26792 9704
rect 26191 9673 26203 9676
rect 26145 9667 26203 9673
rect 26786 9664 26792 9676
rect 26844 9664 26850 9716
rect 27062 9664 27068 9716
rect 27120 9704 27126 9716
rect 27338 9704 27344 9716
rect 27120 9676 27344 9704
rect 27120 9664 27126 9676
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 28902 9664 28908 9716
rect 28960 9704 28966 9716
rect 30929 9707 30987 9713
rect 28960 9676 30420 9704
rect 28960 9664 28966 9676
rect 30392 9674 30420 9676
rect 19475 9608 19564 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 22925 9639 22983 9645
rect 22925 9636 22937 9639
rect 22428 9608 22937 9636
rect 22428 9596 22434 9608
rect 22925 9605 22937 9608
rect 22971 9605 22983 9639
rect 23566 9636 23572 9648
rect 22925 9599 22983 9605
rect 23492 9608 23572 9636
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18506 9528 18512 9580
rect 18564 9528 18570 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9537 18843 9571
rect 18785 9531 18843 9537
rect 19153 9571 19211 9577
rect 19153 9537 19165 9571
rect 19199 9537 19211 9571
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 19153 9531 19211 9537
rect 19352 9540 19809 9568
rect 18064 9500 18092 9528
rect 18708 9500 18736 9531
rect 18064 9472 18736 9500
rect 18230 9392 18236 9444
rect 18288 9432 18294 9444
rect 18690 9432 18696 9444
rect 18288 9404 18696 9432
rect 18288 9392 18294 9404
rect 18690 9392 18696 9404
rect 18748 9432 18754 9444
rect 18800 9432 18828 9531
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19168 9500 19196 9531
rect 19352 9512 19380 9540
rect 19797 9537 19809 9540
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 19978 9528 19984 9580
rect 20036 9528 20042 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 20180 9540 20361 9568
rect 18932 9472 19196 9500
rect 18932 9460 18938 9472
rect 19334 9460 19340 9512
rect 19392 9460 19398 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19475 9472 19533 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 19996 9500 20024 9528
rect 19659 9472 20024 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 18748 9404 18828 9432
rect 18969 9435 19027 9441
rect 18748 9392 18754 9404
rect 18969 9401 18981 9435
rect 19015 9432 19027 9435
rect 19444 9432 19472 9463
rect 20070 9460 20076 9512
rect 20128 9460 20134 9512
rect 20180 9432 20208 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22244 9540 22477 9568
rect 22244 9528 22250 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 22738 9528 22744 9580
rect 22796 9528 22802 9580
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 23017 9571 23075 9577
rect 23017 9537 23029 9571
rect 23063 9568 23075 9571
rect 23382 9568 23388 9580
rect 23063 9540 23388 9568
rect 23063 9537 23075 9540
rect 23017 9531 23075 9537
rect 22848 9500 22876 9531
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23492 9577 23520 9608
rect 23566 9596 23572 9608
rect 23624 9636 23630 9648
rect 27356 9636 27384 9664
rect 23624 9608 23980 9636
rect 27356 9608 27568 9636
rect 23624 9596 23630 9608
rect 23952 9580 23980 9608
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 23661 9571 23719 9577
rect 23661 9537 23673 9571
rect 23707 9568 23719 9571
rect 23750 9568 23756 9580
rect 23707 9540 23756 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23992 9540 24041 9568
rect 23992 9528 23998 9540
rect 24029 9537 24041 9540
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9568 26111 9571
rect 27341 9571 27399 9577
rect 27341 9568 27353 9571
rect 26099 9540 27353 9568
rect 26099 9537 26111 9540
rect 26053 9531 26111 9537
rect 27341 9537 27353 9540
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 23400 9500 23428 9528
rect 24305 9503 24363 9509
rect 24305 9500 24317 9503
rect 22848 9472 23060 9500
rect 23400 9472 24317 9500
rect 19015 9404 20208 9432
rect 19015 9401 19027 9404
rect 18969 9395 19027 9401
rect 23032 9376 23060 9472
rect 24305 9469 24317 9472
rect 24351 9469 24363 9503
rect 24305 9463 24363 9469
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 26329 9503 26387 9509
rect 26329 9500 26341 9503
rect 26292 9472 26341 9500
rect 26292 9460 26298 9472
rect 26329 9469 26341 9472
rect 26375 9500 26387 9503
rect 27246 9500 27252 9512
rect 26375 9472 27252 9500
rect 26375 9469 26387 9472
rect 26329 9463 26387 9469
rect 27246 9460 27252 9472
rect 27304 9460 27310 9512
rect 25958 9392 25964 9444
rect 26016 9432 26022 9444
rect 26973 9435 27031 9441
rect 26973 9432 26985 9435
rect 26016 9404 26985 9432
rect 26016 9392 26022 9404
rect 26973 9401 26985 9404
rect 27019 9401 27031 9435
rect 26973 9395 27031 9401
rect 17331 9336 17540 9364
rect 17586 9324 17592 9376
rect 17644 9324 17650 9376
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 19150 9364 19156 9376
rect 18196 9336 19156 9364
rect 18196 9324 18202 9336
rect 19150 9324 19156 9336
rect 19208 9364 19214 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19208 9336 19257 9364
rect 19208 9324 19214 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19392 9336 19993 9364
rect 19392 9324 19398 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 19981 9327 20039 9333
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 20128 9336 20177 9364
rect 20128 9324 20134 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 20530 9324 20536 9376
rect 20588 9324 20594 9376
rect 22462 9324 22468 9376
rect 22520 9324 22526 9376
rect 23014 9324 23020 9376
rect 23072 9324 23078 9376
rect 25682 9324 25688 9376
rect 25740 9324 25746 9376
rect 27356 9364 27384 9531
rect 27540 9509 27568 9608
rect 28350 9596 28356 9648
rect 28408 9636 28414 9648
rect 30190 9636 30196 9648
rect 28408 9608 30196 9636
rect 28408 9596 28414 9608
rect 30190 9596 30196 9608
rect 30248 9596 30254 9648
rect 30392 9646 30480 9674
rect 30929 9673 30941 9707
rect 30975 9673 30987 9707
rect 30929 9667 30987 9673
rect 30452 9636 30480 9646
rect 30944 9636 30972 9667
rect 31018 9664 31024 9716
rect 31076 9704 31082 9716
rect 31478 9704 31484 9716
rect 31076 9676 31484 9704
rect 31076 9664 31082 9676
rect 31478 9664 31484 9676
rect 31536 9664 31542 9716
rect 32122 9704 32128 9716
rect 31864 9676 32128 9704
rect 30452 9608 30972 9636
rect 31864 9636 31892 9676
rect 32122 9664 32128 9676
rect 32180 9664 32186 9716
rect 34422 9664 34428 9716
rect 34480 9664 34486 9716
rect 37366 9664 37372 9716
rect 37424 9704 37430 9716
rect 37424 9676 38700 9704
rect 37424 9664 37430 9676
rect 38672 9674 38700 9676
rect 34440 9636 34468 9664
rect 31864 9608 31984 9636
rect 34178 9608 34468 9636
rect 30668 9580 30696 9608
rect 30006 9528 30012 9580
rect 30064 9528 30070 9580
rect 30101 9571 30159 9577
rect 30101 9537 30113 9571
rect 30147 9568 30159 9571
rect 30282 9568 30288 9580
rect 30147 9540 30288 9568
rect 30147 9537 30159 9540
rect 30101 9531 30159 9537
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 30377 9572 30435 9577
rect 30377 9571 30512 9572
rect 30377 9537 30389 9571
rect 30423 9568 30512 9571
rect 30423 9544 30604 9568
rect 30423 9537 30435 9544
rect 30484 9540 30604 9544
rect 30377 9531 30435 9537
rect 27433 9503 27491 9509
rect 27433 9469 27445 9503
rect 27479 9469 27491 9503
rect 27433 9463 27491 9469
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 27448 9432 27476 9463
rect 29638 9460 29644 9512
rect 29696 9460 29702 9512
rect 29546 9432 29552 9444
rect 27448 9404 29552 9432
rect 27540 9376 27568 9404
rect 29546 9392 29552 9404
rect 29604 9392 29610 9444
rect 30024 9432 30052 9528
rect 30576 9512 30604 9540
rect 30650 9528 30656 9580
rect 30708 9528 30714 9580
rect 31294 9568 31300 9580
rect 31128 9540 31300 9568
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 31128 9500 31156 9540
rect 31294 9528 31300 9540
rect 31352 9528 31358 9580
rect 31665 9572 31723 9577
rect 31665 9571 31800 9572
rect 31665 9537 31677 9571
rect 31711 9568 31800 9571
rect 31846 9568 31852 9580
rect 31711 9544 31852 9568
rect 31711 9537 31723 9544
rect 31772 9540 31852 9544
rect 31665 9531 31723 9537
rect 30616 9472 31156 9500
rect 31205 9503 31263 9509
rect 30616 9460 30622 9472
rect 31205 9469 31217 9503
rect 31251 9500 31263 9503
rect 31680 9500 31708 9531
rect 31846 9528 31852 9540
rect 31904 9528 31910 9580
rect 31956 9577 31984 9608
rect 34698 9596 34704 9648
rect 34756 9636 34762 9648
rect 38672 9646 39068 9674
rect 39298 9664 39304 9716
rect 39356 9704 39362 9716
rect 39669 9707 39727 9713
rect 39669 9704 39681 9707
rect 39356 9676 39681 9704
rect 39356 9664 39362 9676
rect 39669 9673 39681 9676
rect 39715 9673 39727 9707
rect 39669 9667 39727 9673
rect 41601 9707 41659 9713
rect 41601 9673 41613 9707
rect 41647 9704 41659 9707
rect 41647 9676 42196 9704
rect 41647 9673 41659 9676
rect 41601 9667 41659 9673
rect 37461 9639 37519 9645
rect 37461 9636 37473 9639
rect 34756 9608 34928 9636
rect 34756 9596 34762 9608
rect 34900 9577 34928 9608
rect 35912 9608 37473 9636
rect 35912 9577 35940 9608
rect 37461 9605 37473 9608
rect 37507 9605 37519 9639
rect 37461 9599 37519 9605
rect 31941 9571 31999 9577
rect 31941 9537 31953 9571
rect 31987 9537 31999 9571
rect 31941 9531 31999 9537
rect 34885 9571 34943 9577
rect 34885 9537 34897 9571
rect 34931 9537 34943 9571
rect 34885 9531 34943 9537
rect 35897 9571 35955 9577
rect 35897 9537 35909 9571
rect 35943 9537 35955 9571
rect 36814 9568 36820 9580
rect 35897 9531 35955 9537
rect 36004 9540 36820 9568
rect 31251 9472 31708 9500
rect 31251 9469 31263 9472
rect 31205 9463 31263 9469
rect 34238 9460 34244 9512
rect 34296 9500 34302 9512
rect 36004 9509 36032 9540
rect 36814 9528 36820 9540
rect 36872 9528 36878 9580
rect 36906 9528 36912 9580
rect 36964 9528 36970 9580
rect 37093 9571 37151 9577
rect 37093 9537 37105 9571
rect 37139 9568 37151 9571
rect 37182 9568 37188 9580
rect 37139 9540 37188 9568
rect 37139 9537 37151 9540
rect 37093 9531 37151 9537
rect 37182 9528 37188 9540
rect 37240 9528 37246 9580
rect 38626 9574 38792 9602
rect 38626 9568 38654 9574
rect 38488 9540 38654 9568
rect 38764 9572 38792 9574
rect 38838 9572 38844 9580
rect 38764 9544 38844 9572
rect 34609 9503 34667 9509
rect 34609 9500 34621 9503
rect 34296 9472 34621 9500
rect 34296 9460 34302 9472
rect 34609 9469 34621 9472
rect 34655 9469 34667 9503
rect 34609 9463 34667 9469
rect 35989 9503 36047 9509
rect 35989 9469 36001 9503
rect 36035 9469 36047 9503
rect 35989 9463 36047 9469
rect 36265 9503 36323 9509
rect 36265 9469 36277 9503
rect 36311 9500 36323 9503
rect 37550 9500 37556 9512
rect 36311 9472 37556 9500
rect 36311 9469 36323 9472
rect 36265 9463 36323 9469
rect 37550 9460 37556 9472
rect 37608 9460 37614 9512
rect 37826 9460 37832 9512
rect 37884 9460 37890 9512
rect 38105 9503 38163 9509
rect 38105 9469 38117 9503
rect 38151 9469 38163 9503
rect 38105 9463 38163 9469
rect 30285 9435 30343 9441
rect 30285 9432 30297 9435
rect 30024 9404 30297 9432
rect 30285 9401 30297 9404
rect 30331 9432 30343 9435
rect 37093 9435 37151 9441
rect 30331 9404 31156 9432
rect 30331 9401 30343 9404
rect 30285 9395 30343 9401
rect 27430 9364 27436 9376
rect 27356 9336 27436 9364
rect 27430 9324 27436 9336
rect 27488 9324 27494 9376
rect 27522 9324 27528 9376
rect 27580 9324 27586 9376
rect 29914 9324 29920 9376
rect 29972 9364 29978 9376
rect 30558 9364 30564 9376
rect 29972 9336 30564 9364
rect 29972 9324 29978 9336
rect 30558 9324 30564 9336
rect 30616 9324 30622 9376
rect 31128 9373 31156 9404
rect 37093 9401 37105 9435
rect 37139 9432 37151 9435
rect 37844 9432 37872 9460
rect 37139 9404 37872 9432
rect 38120 9432 38148 9463
rect 38378 9460 38384 9512
rect 38436 9500 38442 9512
rect 38488 9509 38516 9540
rect 38838 9528 38844 9544
rect 38896 9528 38902 9580
rect 38933 9571 38991 9577
rect 38933 9537 38945 9571
rect 38979 9568 38991 9571
rect 39040 9568 39068 9646
rect 39114 9596 39120 9648
rect 39172 9596 39178 9648
rect 41874 9645 41880 9648
rect 41861 9639 41880 9645
rect 41861 9605 41873 9639
rect 41861 9599 41880 9605
rect 41874 9596 41880 9599
rect 41932 9596 41938 9648
rect 42061 9639 42119 9645
rect 42061 9605 42073 9639
rect 42107 9605 42119 9639
rect 42168 9636 42196 9676
rect 43162 9664 43168 9716
rect 43220 9664 43226 9716
rect 43180 9636 43208 9664
rect 42168 9608 43208 9636
rect 42061 9599 42119 9605
rect 38979 9540 39068 9568
rect 41417 9571 41475 9577
rect 38979 9537 38991 9540
rect 38933 9531 38991 9537
rect 41417 9537 41429 9571
rect 41463 9568 41475 9571
rect 41463 9540 41736 9568
rect 41463 9537 41475 9540
rect 41417 9531 41475 9537
rect 38473 9503 38531 9509
rect 38473 9500 38485 9503
rect 38436 9472 38485 9500
rect 38436 9460 38442 9472
rect 38473 9469 38485 9472
rect 38519 9469 38531 9503
rect 38473 9463 38531 9469
rect 38562 9460 38568 9512
rect 38620 9460 38626 9512
rect 38657 9503 38715 9509
rect 38657 9469 38669 9503
rect 38703 9500 38715 9503
rect 39850 9500 39856 9512
rect 38703 9472 39856 9500
rect 38703 9469 38715 9472
rect 38657 9463 38715 9469
rect 39850 9460 39856 9472
rect 39908 9500 39914 9512
rect 40221 9503 40279 9509
rect 40221 9500 40233 9503
rect 39908 9472 40233 9500
rect 39908 9460 39914 9472
rect 40221 9469 40233 9472
rect 40267 9469 40279 9503
rect 40221 9463 40279 9469
rect 39022 9432 39028 9444
rect 38120 9404 39028 9432
rect 37139 9401 37151 9404
rect 37093 9395 37151 9401
rect 39022 9392 39028 9404
rect 39080 9392 39086 9444
rect 41708 9441 41736 9540
rect 42076 9444 42104 9599
rect 42150 9528 42156 9580
rect 42208 9568 42214 9580
rect 42613 9571 42671 9577
rect 42613 9568 42625 9571
rect 42208 9540 42625 9568
rect 42208 9528 42214 9540
rect 42613 9537 42625 9540
rect 42659 9537 42671 9571
rect 42613 9531 42671 9537
rect 42702 9528 42708 9580
rect 42760 9568 42766 9580
rect 42797 9571 42855 9577
rect 42797 9568 42809 9571
rect 42760 9540 42809 9568
rect 42760 9528 42766 9540
rect 42797 9537 42809 9540
rect 42843 9537 42855 9571
rect 42797 9531 42855 9537
rect 41693 9435 41751 9441
rect 41693 9401 41705 9435
rect 41739 9401 41751 9435
rect 41693 9395 41751 9401
rect 42058 9392 42064 9444
rect 42116 9392 42122 9444
rect 31113 9367 31171 9373
rect 31113 9333 31125 9367
rect 31159 9333 31171 9367
rect 31113 9327 31171 9333
rect 31386 9324 31392 9376
rect 31444 9324 31450 9376
rect 31754 9324 31760 9376
rect 31812 9324 31818 9376
rect 33134 9324 33140 9376
rect 33192 9324 33198 9376
rect 38841 9367 38899 9373
rect 38841 9333 38853 9367
rect 38887 9364 38899 9367
rect 39114 9364 39120 9376
rect 38887 9336 39120 9364
rect 38887 9333 38899 9336
rect 38841 9327 38899 9333
rect 39114 9324 39120 9336
rect 39172 9324 39178 9376
rect 39298 9324 39304 9376
rect 39356 9324 39362 9376
rect 41877 9367 41935 9373
rect 41877 9333 41889 9367
rect 41923 9364 41935 9367
rect 42429 9367 42487 9373
rect 42429 9364 42441 9367
rect 41923 9336 42441 9364
rect 41923 9333 41935 9336
rect 41877 9327 41935 9333
rect 42429 9333 42441 9336
rect 42475 9333 42487 9367
rect 42429 9327 42487 9333
rect 1104 9274 45172 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 45172 9274
rect 1104 9200 45172 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 6914 9160 6920 9172
rect 1627 9132 6920 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12802 9160 12808 9172
rect 12032 9132 12808 9160
rect 12032 9120 12038 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 13412 9132 13461 9160
rect 13412 9120 13418 9132
rect 13449 9129 13461 9132
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 13814 9120 13820 9172
rect 13872 9120 13878 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14884 9132 14933 9160
rect 14884 9120 14890 9132
rect 14921 9129 14933 9132
rect 14967 9129 14979 9163
rect 14921 9123 14979 9129
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 17126 9160 17132 9172
rect 15151 9132 17132 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17770 9160 17776 9172
rect 17420 9132 17776 9160
rect 12986 9052 12992 9104
rect 13044 9052 13050 9104
rect 15473 9095 15531 9101
rect 13464 9064 14596 9092
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11572 8996 11989 9024
rect 11572 8984 11578 8996
rect 11977 8993 11989 8996
rect 12023 9024 12035 9027
rect 13004 9024 13032 9052
rect 12023 8996 13032 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12250 8956 12256 8968
rect 11848 8928 12256 8956
rect 11848 8916 11854 8928
rect 12250 8916 12256 8928
rect 12308 8956 12314 8968
rect 13464 8965 13492 9064
rect 13648 8996 13860 9024
rect 13648 8965 13676 8996
rect 13832 8968 13860 8996
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12308 8928 12357 8956
rect 12308 8916 12314 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 11698 8848 11704 8900
rect 11756 8848 11762 8900
rect 13740 8888 13768 8919
rect 13814 8916 13820 8968
rect 13872 8916 13878 8968
rect 13924 8965 13952 9064
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 14056 8996 14105 9024
rect 14056 8984 14062 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 13909 8959 13967 8965
rect 13909 8925 13921 8959
rect 13955 8925 13967 8959
rect 13909 8919 13967 8925
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8925 14243 8959
rect 14185 8919 14243 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14568 8956 14596 9064
rect 15473 9061 15485 9095
rect 15519 9092 15531 9095
rect 15519 9064 15608 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 15580 9024 15608 9064
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 15712 9064 16712 9092
rect 15712 9052 15718 9064
rect 16390 9024 16396 9036
rect 14700 8996 15516 9024
rect 15580 8996 16396 9024
rect 14700 8984 14706 8996
rect 15488 8965 15516 8996
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14568 8928 15301 8956
rect 14200 8888 14228 8919
rect 13740 8860 14228 8888
rect 13740 8832 13768 8860
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13078 8820 13084 8832
rect 12492 8792 13084 8820
rect 12492 8780 12498 8792
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13722 8780 13728 8832
rect 13780 8780 13786 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14476 8820 14504 8919
rect 14568 8900 14596 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8956 15531 8959
rect 15838 8956 15844 8968
rect 15519 8928 15844 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16482 8956 16488 8968
rect 16264 8928 16488 8956
rect 16264 8916 16270 8928
rect 16482 8916 16488 8928
rect 16540 8956 16546 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16540 8928 16589 8956
rect 16540 8916 16546 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16684 8956 16712 9064
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 16945 9095 17003 9101
rect 16945 9092 16957 9095
rect 16816 9064 16957 9092
rect 16816 9052 16822 9064
rect 16945 9061 16957 9064
rect 16991 9092 17003 9095
rect 17420 9092 17448 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18046 9120 18052 9172
rect 18104 9120 18110 9172
rect 19981 9163 20039 9169
rect 19981 9129 19993 9163
rect 20027 9160 20039 9163
rect 20346 9160 20352 9172
rect 20027 9132 20352 9160
rect 20027 9129 20039 9132
rect 19981 9123 20039 9129
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22520 9132 22968 9160
rect 22520 9120 22526 9132
rect 16991 9064 17448 9092
rect 17497 9095 17555 9101
rect 16991 9061 17003 9064
rect 16945 9055 17003 9061
rect 17497 9061 17509 9095
rect 17543 9092 17555 9095
rect 17954 9092 17960 9104
rect 17543 9064 17960 9092
rect 17543 9061 17555 9064
rect 17497 9055 17555 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 22373 9095 22431 9101
rect 19996 9064 20300 9092
rect 19996 9036 20024 9064
rect 17052 8996 17908 9024
rect 16761 8959 16819 8965
rect 16761 8956 16773 8959
rect 16684 8928 16773 8956
rect 16577 8919 16635 8925
rect 16761 8925 16773 8928
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 14550 8848 14556 8900
rect 14608 8848 14614 8900
rect 16666 8848 16672 8900
rect 16724 8848 16730 8900
rect 14642 8820 14648 8832
rect 13872 8792 14648 8820
rect 13872 8780 13878 8792
rect 14642 8780 14648 8792
rect 14700 8820 14706 8832
rect 14930 8823 14988 8829
rect 14930 8820 14942 8823
rect 14700 8792 14942 8820
rect 14700 8780 14706 8792
rect 14930 8789 14942 8792
rect 14976 8820 14988 8823
rect 15930 8820 15936 8832
rect 14976 8792 15936 8820
rect 14976 8789 14988 8792
rect 14930 8783 14988 8789
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 16865 8820 16893 8919
rect 17052 8832 17080 8996
rect 17402 8965 17408 8968
rect 17372 8959 17408 8965
rect 17372 8925 17384 8959
rect 17372 8919 17408 8925
rect 17402 8916 17408 8919
rect 17460 8916 17466 8968
rect 17880 8965 17908 8996
rect 19978 8984 19984 9036
rect 20036 8984 20042 9036
rect 20145 9027 20203 9033
rect 20145 8993 20157 9027
rect 20191 9024 20203 9027
rect 20191 8993 20208 9024
rect 20145 8987 20208 8993
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 17126 8848 17132 8900
rect 17184 8888 17190 8900
rect 17604 8888 17632 8919
rect 19518 8916 19524 8968
rect 19576 8916 19582 8968
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20180 8956 20208 8987
rect 20272 8965 20300 9064
rect 22373 9061 22385 9095
rect 22419 9092 22431 9095
rect 22554 9092 22560 9104
rect 22419 9064 22560 9092
rect 22419 9061 22431 9064
rect 22373 9055 22431 9061
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 19751 8928 20208 8956
rect 20257 8959 20315 8965
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20622 8956 20628 8968
rect 20395 8928 20628 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22940 8965 22968 9132
rect 23382 9120 23388 9172
rect 23440 9120 23446 9172
rect 25682 9120 25688 9172
rect 25740 9120 25746 9172
rect 25774 9120 25780 9172
rect 25832 9160 25838 9172
rect 25869 9163 25927 9169
rect 25869 9160 25881 9163
rect 25832 9132 25881 9160
rect 25832 9120 25838 9132
rect 25869 9129 25881 9132
rect 25915 9129 25927 9163
rect 25869 9123 25927 9129
rect 27338 9120 27344 9172
rect 27396 9120 27402 9172
rect 27522 9120 27528 9172
rect 27580 9120 27586 9172
rect 28074 9120 28080 9172
rect 28132 9120 28138 9172
rect 28442 9120 28448 9172
rect 28500 9160 28506 9172
rect 28721 9163 28779 9169
rect 28721 9160 28733 9163
rect 28500 9132 28733 9160
rect 28500 9120 28506 9132
rect 28721 9129 28733 9132
rect 28767 9129 28779 9163
rect 28721 9123 28779 9129
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9129 28963 9163
rect 28905 9123 28963 9129
rect 23400 9092 23428 9120
rect 25700 9092 25728 9120
rect 23400 9064 23980 9092
rect 23952 9033 23980 9064
rect 25148 9064 25728 9092
rect 26329 9095 26387 9101
rect 25148 9033 25176 9064
rect 26329 9061 26341 9095
rect 26375 9061 26387 9095
rect 27540 9092 27568 9120
rect 28920 9092 28948 9123
rect 30282 9120 30288 9172
rect 30340 9120 30346 9172
rect 30509 9163 30567 9169
rect 30509 9129 30521 9163
rect 30555 9160 30567 9163
rect 31386 9160 31392 9172
rect 30555 9132 31392 9160
rect 30555 9129 30567 9132
rect 30509 9123 30567 9129
rect 31386 9120 31392 9132
rect 31444 9120 31450 9172
rect 31754 9120 31760 9172
rect 31812 9160 31818 9172
rect 31849 9163 31907 9169
rect 31849 9160 31861 9163
rect 31812 9132 31861 9160
rect 31812 9120 31818 9132
rect 31849 9129 31861 9132
rect 31895 9129 31907 9163
rect 31849 9123 31907 9129
rect 32217 9163 32275 9169
rect 32217 9129 32229 9163
rect 32263 9160 32275 9163
rect 32398 9160 32404 9172
rect 32263 9132 32404 9160
rect 32263 9129 32275 9132
rect 32217 9123 32275 9129
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 33134 9120 33140 9172
rect 33192 9120 33198 9172
rect 37366 9120 37372 9172
rect 37424 9120 37430 9172
rect 37553 9163 37611 9169
rect 37553 9129 37565 9163
rect 37599 9160 37611 9163
rect 38562 9160 38568 9172
rect 37599 9132 38568 9160
rect 37599 9129 37611 9132
rect 37553 9123 37611 9129
rect 38562 9120 38568 9132
rect 38620 9120 38626 9172
rect 38930 9120 38936 9172
rect 38988 9120 38994 9172
rect 39298 9120 39304 9172
rect 39356 9160 39362 9172
rect 40037 9163 40095 9169
rect 40037 9160 40049 9163
rect 39356 9132 40049 9160
rect 39356 9120 39362 9132
rect 40037 9129 40049 9132
rect 40083 9129 40095 9163
rect 40037 9123 40095 9129
rect 41874 9120 41880 9172
rect 41932 9120 41938 9172
rect 30098 9092 30104 9104
rect 26329 9055 26387 9061
rect 26712 9064 27568 9092
rect 28736 9064 30104 9092
rect 23937 9027 23995 9033
rect 23124 8996 23796 9024
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22336 8928 22569 8956
rect 22336 8916 22342 8928
rect 22557 8925 22569 8928
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23124 8956 23152 8996
rect 23072 8928 23152 8956
rect 23072 8916 23078 8928
rect 23198 8916 23204 8968
rect 23256 8916 23262 8968
rect 23768 8956 23796 8996
rect 23937 8993 23949 9027
rect 23983 8993 23995 9027
rect 23937 8987 23995 8993
rect 25133 9027 25191 9033
rect 25133 8993 25145 9027
rect 25179 8993 25191 9027
rect 25133 8987 25191 8993
rect 25314 8984 25320 9036
rect 25372 9024 25378 9036
rect 26142 9024 26148 9036
rect 25372 8996 26148 9024
rect 25372 8984 25378 8996
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 24394 8956 24400 8968
rect 23768 8928 24400 8956
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 26344 8956 26372 9055
rect 26712 8965 26740 9064
rect 26973 9027 27031 9033
rect 26973 8993 26985 9027
rect 27019 9024 27031 9027
rect 27338 9024 27344 9036
rect 27019 8996 27344 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 27338 8984 27344 8996
rect 27396 9024 27402 9036
rect 28261 9027 28319 9033
rect 27396 8996 28120 9024
rect 27396 8984 27402 8996
rect 25096 8928 26372 8956
rect 26697 8959 26755 8965
rect 25096 8916 25102 8928
rect 26697 8925 26709 8959
rect 26743 8925 26755 8959
rect 26697 8919 26755 8925
rect 27522 8916 27528 8968
rect 27580 8916 27586 8968
rect 28092 8965 28120 8996
rect 28261 8993 28273 9027
rect 28307 8993 28319 9027
rect 28261 8987 28319 8993
rect 28077 8959 28135 8965
rect 28077 8925 28089 8959
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 17184 8860 17632 8888
rect 19536 8888 19564 8916
rect 19797 8891 19855 8897
rect 19797 8888 19809 8891
rect 19536 8860 19809 8888
rect 17184 8848 17190 8860
rect 19797 8857 19809 8860
rect 19843 8857 19855 8891
rect 19797 8851 19855 8857
rect 19981 8891 20039 8897
rect 19981 8857 19993 8891
rect 20027 8857 20039 8891
rect 19981 8851 20039 8857
rect 16816 8792 16893 8820
rect 16816 8780 16822 8792
rect 17034 8780 17040 8832
rect 17092 8780 17098 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17313 8823 17371 8829
rect 17313 8820 17325 8823
rect 17276 8792 17325 8820
rect 17276 8780 17282 8792
rect 17313 8789 17325 8792
rect 17359 8789 17371 8823
rect 17313 8783 17371 8789
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17644 8792 17693 8820
rect 17644 8780 17650 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 19996 8820 20024 8851
rect 20070 8848 20076 8900
rect 20128 8848 20134 8900
rect 20530 8848 20536 8900
rect 20588 8848 20594 8900
rect 22186 8848 22192 8900
rect 22244 8888 22250 8900
rect 22649 8891 22707 8897
rect 22649 8888 22661 8891
rect 22244 8860 22661 8888
rect 22244 8848 22250 8860
rect 22649 8857 22661 8860
rect 22695 8857 22707 8891
rect 22649 8851 22707 8857
rect 22741 8891 22799 8897
rect 22741 8857 22753 8891
rect 22787 8888 22799 8891
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 22787 8860 23121 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 23750 8848 23756 8900
rect 23808 8888 23814 8900
rect 25593 8891 25651 8897
rect 23808 8860 25268 8888
rect 23808 8848 23814 8860
rect 20548 8820 20576 8848
rect 25240 8832 25268 8860
rect 25593 8857 25605 8891
rect 25639 8888 25651 8891
rect 25774 8888 25780 8900
rect 25639 8860 25780 8888
rect 25639 8857 25651 8860
rect 25593 8851 25651 8857
rect 25774 8848 25780 8860
rect 25832 8848 25838 8900
rect 26789 8891 26847 8897
rect 26789 8857 26801 8891
rect 26835 8888 26847 8891
rect 28166 8888 28172 8900
rect 26835 8860 28172 8888
rect 26835 8857 26847 8860
rect 26789 8851 26847 8857
rect 28166 8848 28172 8860
rect 28224 8848 28230 8900
rect 28276 8888 28304 8987
rect 28350 8916 28356 8968
rect 28408 8916 28414 8968
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8956 28503 8959
rect 28534 8956 28540 8968
rect 28491 8928 28540 8956
rect 28491 8925 28503 8928
rect 28445 8919 28503 8925
rect 28534 8916 28540 8928
rect 28592 8956 28598 8968
rect 28736 8956 28764 9064
rect 30098 9052 30104 9064
rect 30156 9052 30162 9104
rect 30834 9052 30840 9104
rect 30892 9052 30898 9104
rect 30193 9027 30251 9033
rect 30193 9024 30205 9027
rect 28592 8928 28764 8956
rect 28828 8996 30205 9024
rect 28592 8916 28598 8928
rect 28828 8888 28856 8996
rect 30193 8993 30205 8996
rect 30239 9024 30251 9027
rect 30239 8996 30328 9024
rect 30239 8993 30251 8996
rect 30193 8987 30251 8993
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8956 29607 8959
rect 29638 8956 29644 8968
rect 29595 8928 29644 8956
rect 29595 8925 29607 8928
rect 29549 8919 29607 8925
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 29730 8916 29736 8968
rect 29788 8916 29794 8968
rect 29822 8916 29828 8968
rect 29880 8916 29886 8968
rect 29963 8959 30021 8965
rect 29963 8956 29975 8959
rect 29932 8946 29975 8956
rect 28902 8897 28908 8900
rect 28276 8860 28856 8888
rect 28889 8891 28908 8897
rect 28889 8857 28901 8891
rect 28889 8851 28908 8857
rect 28902 8848 28908 8851
rect 28960 8848 28966 8900
rect 29089 8891 29147 8897
rect 29089 8888 29101 8891
rect 29012 8860 29101 8888
rect 29012 8832 29040 8860
rect 29089 8857 29101 8860
rect 29135 8857 29147 8891
rect 29089 8851 29147 8857
rect 29178 8848 29184 8900
rect 29236 8888 29242 8900
rect 29840 8888 29868 8916
rect 29914 8894 29920 8946
rect 29972 8925 29975 8946
rect 30009 8925 30021 8959
rect 30300 8953 30328 8996
rect 30466 8984 30472 9036
rect 30524 9024 30530 9036
rect 31570 9024 31576 9036
rect 30524 8996 31064 9024
rect 30524 8984 30530 8996
rect 30452 8953 30696 8956
rect 30300 8928 30696 8953
rect 30300 8925 30480 8928
rect 29972 8919 30021 8925
rect 29972 8894 29978 8919
rect 29236 8860 29868 8888
rect 29236 8848 29242 8860
rect 30190 8848 30196 8900
rect 30248 8888 30254 8900
rect 30668 8897 30696 8928
rect 30742 8916 30748 8968
rect 30800 8916 30806 8968
rect 30929 8959 30987 8965
rect 30929 8956 30941 8959
rect 30852 8928 30941 8956
rect 30852 8900 30880 8928
rect 30929 8925 30941 8928
rect 30975 8925 30987 8959
rect 30929 8919 30987 8925
rect 30437 8891 30495 8897
rect 30437 8888 30449 8891
rect 30248 8860 30449 8888
rect 30248 8848 30254 8860
rect 30437 8857 30449 8860
rect 30483 8857 30495 8891
rect 30437 8851 30495 8857
rect 30653 8891 30711 8897
rect 30653 8857 30665 8891
rect 30699 8857 30711 8891
rect 30653 8851 30711 8857
rect 19996 8792 20576 8820
rect 17681 8783 17739 8789
rect 23382 8780 23388 8832
rect 23440 8780 23446 8832
rect 23845 8823 23903 8829
rect 23845 8789 23857 8823
rect 23891 8820 23903 8823
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 23891 8792 24685 8820
rect 23891 8789 23903 8792
rect 23845 8783 23903 8789
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 28994 8780 29000 8832
rect 29052 8780 29058 8832
rect 29638 8780 29644 8832
rect 29696 8820 29702 8832
rect 30282 8820 30288 8832
rect 29696 8792 30288 8820
rect 29696 8780 29702 8792
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 30452 8820 30480 8851
rect 30834 8848 30840 8900
rect 30892 8848 30898 8900
rect 31036 8888 31064 8996
rect 31220 8996 31576 9024
rect 31220 8965 31248 8996
rect 31570 8984 31576 8996
rect 31628 9024 31634 9036
rect 33152 9024 33180 9120
rect 33505 9027 33563 9033
rect 33505 9024 33517 9027
rect 31628 8996 32076 9024
rect 33152 8996 33517 9024
rect 31628 8984 31634 8996
rect 31205 8959 31263 8965
rect 31205 8925 31217 8959
rect 31251 8925 31263 8959
rect 31205 8919 31263 8925
rect 31846 8916 31852 8968
rect 31904 8916 31910 8968
rect 32048 8965 32076 8996
rect 33505 8993 33517 8996
rect 33551 8993 33563 9027
rect 33505 8987 33563 8993
rect 32033 8959 32091 8965
rect 32033 8925 32045 8959
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32122 8916 32128 8968
rect 32180 8916 32186 8968
rect 32309 8959 32367 8965
rect 32309 8925 32321 8959
rect 32355 8925 32367 8959
rect 37384 8956 37412 9120
rect 38948 9092 38976 9120
rect 39853 9095 39911 9101
rect 39853 9092 39865 9095
rect 38948 9064 39865 9092
rect 39853 9061 39865 9064
rect 39899 9061 39911 9095
rect 39853 9055 39911 9061
rect 41690 8984 41696 9036
rect 41748 9024 41754 9036
rect 42702 9024 42708 9036
rect 41748 8996 41828 9024
rect 41748 8984 41754 8996
rect 38105 8959 38163 8965
rect 38105 8956 38117 8959
rect 37384 8928 38117 8956
rect 32309 8919 32367 8925
rect 38105 8925 38117 8928
rect 38151 8925 38163 8959
rect 38105 8919 38163 8925
rect 38289 8959 38347 8965
rect 38289 8925 38301 8959
rect 38335 8956 38347 8959
rect 38378 8956 38384 8968
rect 38335 8928 38384 8956
rect 38335 8925 38347 8928
rect 38289 8919 38347 8925
rect 31389 8891 31447 8897
rect 31389 8888 31401 8891
rect 31036 8860 31401 8888
rect 31389 8857 31401 8860
rect 31435 8857 31447 8891
rect 31389 8851 31447 8857
rect 31478 8848 31484 8900
rect 31536 8888 31542 8900
rect 32324 8888 32352 8919
rect 38378 8916 38384 8928
rect 38436 8916 38442 8968
rect 41800 8965 41828 8996
rect 41984 8996 42708 9024
rect 41984 8968 42012 8996
rect 42702 8984 42708 8996
rect 42760 8984 42766 9036
rect 41785 8959 41843 8965
rect 41785 8925 41797 8959
rect 41831 8925 41843 8959
rect 41785 8919 41843 8925
rect 41966 8916 41972 8968
rect 42024 8916 42030 8968
rect 42242 8916 42248 8968
rect 42300 8956 42306 8968
rect 42429 8959 42487 8965
rect 42429 8956 42441 8959
rect 42300 8928 42441 8956
rect 42300 8916 42306 8928
rect 42429 8925 42441 8928
rect 42475 8925 42487 8959
rect 42429 8919 42487 8925
rect 42610 8916 42616 8968
rect 42668 8916 42674 8968
rect 42797 8959 42855 8965
rect 42797 8925 42809 8959
rect 42843 8956 42855 8959
rect 42886 8956 42892 8968
rect 42843 8928 42892 8956
rect 42843 8925 42855 8928
rect 42797 8919 42855 8925
rect 42886 8916 42892 8928
rect 42944 8916 42950 8968
rect 31536 8860 32352 8888
rect 31536 8848 31542 8860
rect 36906 8848 36912 8900
rect 36964 8888 36970 8900
rect 37737 8891 37795 8897
rect 37737 8888 37749 8891
rect 36964 8860 37749 8888
rect 36964 8848 36970 8860
rect 37737 8857 37749 8860
rect 37783 8888 37795 8891
rect 39022 8888 39028 8900
rect 37783 8860 39028 8888
rect 37783 8857 37795 8860
rect 37737 8851 37795 8857
rect 39022 8848 39028 8860
rect 39080 8848 39086 8900
rect 39482 8848 39488 8900
rect 39540 8888 39546 8900
rect 40221 8891 40279 8897
rect 40221 8888 40233 8891
rect 39540 8860 40233 8888
rect 39540 8848 39546 8860
rect 40221 8857 40233 8860
rect 40267 8888 40279 8891
rect 42058 8888 42064 8900
rect 40267 8860 42064 8888
rect 40267 8857 40279 8860
rect 40221 8851 40279 8857
rect 42058 8848 42064 8860
rect 42116 8848 42122 8900
rect 42521 8891 42579 8897
rect 42521 8857 42533 8891
rect 42567 8888 42579 8891
rect 43070 8888 43076 8900
rect 42567 8860 43076 8888
rect 42567 8857 42579 8860
rect 42521 8851 42579 8857
rect 43070 8848 43076 8860
rect 43128 8848 43134 8900
rect 31110 8820 31116 8832
rect 30452 8792 31116 8820
rect 31110 8780 31116 8792
rect 31168 8780 31174 8832
rect 31570 8780 31576 8832
rect 31628 8780 31634 8832
rect 31662 8780 31668 8832
rect 31720 8780 31726 8832
rect 34146 8780 34152 8832
rect 34204 8780 34210 8832
rect 36814 8780 36820 8832
rect 36872 8820 36878 8832
rect 37090 8820 37096 8832
rect 36872 8792 37096 8820
rect 36872 8780 36878 8792
rect 37090 8780 37096 8792
rect 37148 8820 37154 8832
rect 37527 8823 37585 8829
rect 37527 8820 37539 8823
rect 37148 8792 37539 8820
rect 37148 8780 37154 8792
rect 37527 8789 37539 8792
rect 37573 8789 37585 8823
rect 37527 8783 37585 8789
rect 38289 8823 38347 8829
rect 38289 8789 38301 8823
rect 38335 8820 38347 8823
rect 39206 8820 39212 8832
rect 38335 8792 39212 8820
rect 38335 8789 38347 8792
rect 38289 8783 38347 8789
rect 39206 8780 39212 8792
rect 39264 8820 39270 8832
rect 40011 8823 40069 8829
rect 40011 8820 40023 8823
rect 39264 8792 40023 8820
rect 39264 8780 39270 8792
rect 40011 8789 40023 8792
rect 40057 8789 40069 8823
rect 40011 8783 40069 8789
rect 42981 8823 43039 8829
rect 42981 8789 42993 8823
rect 43027 8820 43039 8823
rect 43346 8820 43352 8832
rect 43027 8792 43352 8820
rect 43027 8789 43039 8792
rect 42981 8783 43039 8789
rect 43346 8780 43352 8792
rect 43404 8780 43410 8832
rect 1104 8730 45172 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 45172 8730
rect 1104 8656 45172 8678
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 15565 8619 15623 8625
rect 11756 8588 15424 8616
rect 11756 8576 11762 8588
rect 11900 8557 11928 8588
rect 11885 8551 11943 8557
rect 11885 8517 11897 8551
rect 11931 8517 11943 8551
rect 13722 8548 13728 8560
rect 11885 8511 11943 8517
rect 12544 8520 13728 8548
rect 12544 8492 12572 8520
rect 13722 8508 13728 8520
rect 13780 8548 13786 8560
rect 14826 8548 14832 8560
rect 13780 8520 14832 8548
rect 13780 8508 13786 8520
rect 14826 8508 14832 8520
rect 14884 8548 14890 8560
rect 15396 8548 15424 8588
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15654 8616 15660 8628
rect 15611 8588 15660 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 15988 8588 17233 8616
rect 15988 8576 15994 8588
rect 17221 8585 17233 8588
rect 17267 8616 17279 8619
rect 17589 8619 17647 8625
rect 17267 8588 17448 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 16482 8548 16488 8560
rect 14884 8520 15332 8548
rect 15396 8520 16488 8548
rect 14884 8508 14890 8520
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12526 8480 12532 8492
rect 12115 8452 12532 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 14366 8480 14372 8492
rect 14047 8452 14372 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 14366 8440 14372 8452
rect 14424 8480 14430 8492
rect 15102 8480 15108 8492
rect 14424 8452 15108 8480
rect 14424 8440 14430 8452
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 15304 8489 15332 8520
rect 16482 8508 16488 8520
rect 16540 8548 16546 8560
rect 17420 8548 17448 8588
rect 17589 8585 17601 8619
rect 17635 8616 17647 8619
rect 20070 8616 20076 8628
rect 17635 8588 20076 8616
rect 17635 8585 17647 8588
rect 17589 8579 17647 8585
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 22002 8616 22008 8628
rect 21867 8588 22008 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 23382 8576 23388 8628
rect 23440 8576 23446 8628
rect 24394 8576 24400 8628
rect 24452 8576 24458 8628
rect 24857 8619 24915 8625
rect 24857 8585 24869 8619
rect 24903 8616 24915 8619
rect 25038 8616 25044 8628
rect 24903 8588 25044 8616
rect 24903 8585 24915 8588
rect 24857 8579 24915 8585
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25222 8576 25228 8628
rect 25280 8576 25286 8628
rect 25590 8576 25596 8628
rect 25648 8616 25654 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 25648 8588 25697 8616
rect 25648 8576 25654 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 26326 8576 26332 8628
rect 26384 8616 26390 8628
rect 26973 8619 27031 8625
rect 26973 8616 26985 8619
rect 26384 8588 26985 8616
rect 26384 8576 26390 8588
rect 26973 8585 26985 8588
rect 27019 8585 27031 8619
rect 26973 8579 27031 8585
rect 27433 8619 27491 8625
rect 27433 8585 27445 8619
rect 27479 8616 27491 8619
rect 28166 8616 28172 8628
rect 27479 8588 28172 8616
rect 27479 8585 27491 8588
rect 27433 8579 27491 8585
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 28261 8619 28319 8625
rect 28261 8585 28273 8619
rect 28307 8616 28319 8619
rect 28350 8616 28356 8628
rect 28307 8588 28356 8616
rect 28307 8585 28319 8588
rect 28261 8579 28319 8585
rect 28350 8576 28356 8588
rect 28408 8576 28414 8628
rect 28442 8576 28448 8628
rect 28500 8576 28506 8628
rect 29086 8616 29092 8628
rect 28644 8588 29092 8616
rect 16540 8520 17356 8548
rect 17420 8520 17632 8548
rect 16540 8508 16546 8520
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 15470 8440 15476 8492
rect 15528 8440 15534 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 15580 8452 17049 8480
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 15580 8412 15608 8452
rect 17037 8449 17049 8452
rect 17083 8480 17095 8483
rect 17126 8480 17132 8492
rect 17083 8452 17132 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17328 8489 17356 8520
rect 17604 8492 17632 8520
rect 19886 8508 19892 8560
rect 19944 8548 19950 8560
rect 20622 8548 20628 8560
rect 19944 8520 20628 8548
rect 19944 8508 19950 8520
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 23400 8548 23428 8576
rect 28460 8548 28488 8576
rect 22020 8520 23428 8548
rect 28184 8520 28488 8548
rect 28537 8551 28595 8557
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 22020 8489 22048 8520
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8480 22155 8483
rect 24765 8483 24823 8489
rect 22143 8452 22232 8480
rect 22143 8449 22155 8452
rect 22097 8443 22155 8449
rect 22204 8424 22232 8452
rect 24765 8449 24777 8483
rect 24811 8480 24823 8483
rect 25593 8483 25651 8489
rect 25593 8480 25605 8483
rect 24811 8452 25605 8480
rect 24811 8449 24823 8452
rect 24765 8443 24823 8449
rect 25593 8449 25605 8452
rect 25639 8480 25651 8483
rect 26694 8480 26700 8492
rect 25639 8452 26700 8480
rect 25639 8449 25651 8452
rect 25593 8443 25651 8449
rect 26694 8440 26700 8452
rect 26752 8440 26758 8492
rect 27338 8440 27344 8492
rect 27396 8440 27402 8492
rect 28184 8489 28212 8520
rect 28537 8517 28549 8551
rect 28583 8548 28595 8551
rect 28644 8548 28672 8588
rect 29086 8576 29092 8588
rect 29144 8616 29150 8628
rect 29638 8616 29644 8628
rect 29144 8588 29644 8616
rect 29144 8576 29150 8588
rect 29638 8576 29644 8588
rect 29696 8576 29702 8628
rect 29822 8576 29828 8628
rect 29880 8616 29886 8628
rect 30834 8616 30840 8628
rect 29880 8588 30840 8616
rect 29880 8576 29886 8588
rect 30834 8576 30840 8588
rect 30892 8576 30898 8628
rect 31110 8576 31116 8628
rect 31168 8616 31174 8628
rect 31941 8619 31999 8625
rect 31941 8616 31953 8619
rect 31168 8588 31953 8616
rect 31168 8576 31174 8588
rect 31941 8585 31953 8588
rect 31987 8616 31999 8619
rect 32122 8616 32128 8628
rect 31987 8588 32128 8616
rect 31987 8585 31999 8588
rect 31941 8579 31999 8585
rect 32122 8576 32128 8588
rect 32180 8576 32186 8628
rect 34146 8576 34152 8628
rect 34204 8576 34210 8628
rect 42242 8616 42248 8628
rect 40420 8588 42248 8616
rect 31297 8551 31355 8557
rect 28583 8520 28672 8548
rect 28583 8517 28595 8520
rect 28537 8511 28595 8517
rect 28644 8489 28672 8520
rect 28828 8520 29224 8548
rect 28169 8483 28227 8489
rect 28169 8449 28181 8483
rect 28215 8449 28227 8483
rect 28169 8443 28227 8449
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8449 28411 8483
rect 28353 8443 28411 8449
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 14608 8384 15608 8412
rect 14608 8372 14614 8384
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 16942 8412 16948 8424
rect 15896 8384 16948 8412
rect 15896 8372 15902 8384
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 18966 8412 18972 8424
rect 17451 8384 18972 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 21818 8372 21824 8424
rect 21876 8372 21882 8424
rect 22186 8372 22192 8424
rect 22244 8372 22250 8424
rect 25041 8415 25099 8421
rect 25041 8381 25053 8415
rect 25087 8412 25099 8415
rect 25314 8412 25320 8424
rect 25087 8384 25320 8412
rect 25087 8381 25099 8384
rect 25041 8375 25099 8381
rect 25314 8372 25320 8384
rect 25372 8372 25378 8424
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 27246 8372 27252 8424
rect 27304 8412 27310 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 27304 8384 27537 8412
rect 27304 8372 27310 8384
rect 27525 8381 27537 8384
rect 27571 8381 27583 8415
rect 27525 8375 27583 8381
rect 27890 8372 27896 8424
rect 27948 8412 27954 8424
rect 27985 8415 28043 8421
rect 27985 8412 27997 8415
rect 27948 8384 27997 8412
rect 27948 8372 27954 8384
rect 27985 8381 27997 8384
rect 28031 8381 28043 8415
rect 28368 8412 28396 8443
rect 28828 8412 28856 8520
rect 29196 8492 29224 8520
rect 29472 8520 31248 8548
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8480 28963 8483
rect 28994 8480 29000 8492
rect 28951 8452 29000 8480
rect 28951 8449 28963 8452
rect 28905 8443 28963 8449
rect 28368 8384 28856 8412
rect 28920 8412 28948 8443
rect 28994 8440 29000 8452
rect 29052 8440 29058 8492
rect 29178 8440 29184 8492
rect 29236 8440 29242 8492
rect 29472 8489 29500 8520
rect 29457 8483 29515 8489
rect 29457 8449 29469 8483
rect 29503 8449 29515 8483
rect 29457 8443 29515 8449
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8480 29699 8483
rect 30006 8480 30012 8492
rect 29687 8452 30012 8480
rect 29687 8449 29699 8452
rect 29641 8443 29699 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 30116 8489 30144 8520
rect 30101 8483 30159 8489
rect 30101 8449 30113 8483
rect 30147 8449 30159 8483
rect 30101 8443 30159 8449
rect 30190 8440 30196 8492
rect 30248 8440 30254 8492
rect 30282 8440 30288 8492
rect 30340 8480 30346 8492
rect 30377 8483 30435 8489
rect 30377 8480 30389 8483
rect 30340 8452 30389 8480
rect 30340 8440 30346 8452
rect 30377 8449 30389 8452
rect 30423 8449 30435 8483
rect 30377 8443 30435 8449
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 30834 8440 30840 8492
rect 30892 8440 30898 8492
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8480 30987 8483
rect 31018 8480 31024 8492
rect 30975 8452 31024 8480
rect 30975 8449 30987 8452
rect 30929 8443 30987 8449
rect 31018 8440 31024 8452
rect 31076 8440 31082 8492
rect 31113 8483 31171 8489
rect 31113 8449 31125 8483
rect 31159 8449 31171 8483
rect 31220 8480 31248 8520
rect 31297 8517 31309 8551
rect 31343 8548 31355 8551
rect 34164 8548 34192 8576
rect 34241 8551 34299 8557
rect 34241 8548 34253 8551
rect 31343 8520 31754 8548
rect 34164 8520 34253 8548
rect 31343 8517 31355 8520
rect 31297 8511 31355 8517
rect 31726 8492 31754 8520
rect 34241 8517 34253 8520
rect 34287 8517 34299 8551
rect 34241 8511 34299 8517
rect 35989 8551 36047 8557
rect 35989 8517 36001 8551
rect 36035 8548 36047 8551
rect 36998 8548 37004 8560
rect 36035 8520 37004 8548
rect 36035 8517 36047 8520
rect 35989 8511 36047 8517
rect 36998 8508 37004 8520
rect 37056 8508 37062 8560
rect 40420 8492 40448 8588
rect 42242 8576 42248 8588
rect 42300 8576 42306 8628
rect 42610 8576 42616 8628
rect 42668 8616 42674 8628
rect 43165 8619 43223 8625
rect 43165 8616 43177 8619
rect 42668 8588 43177 8616
rect 42668 8576 42674 8588
rect 43165 8585 43177 8588
rect 43211 8585 43223 8619
rect 43165 8579 43223 8585
rect 41049 8551 41107 8557
rect 41049 8548 41061 8551
rect 40512 8520 41061 8548
rect 31570 8480 31576 8492
rect 31220 8452 31576 8480
rect 31113 8443 31171 8449
rect 30745 8415 30803 8421
rect 28920 8384 29868 8412
rect 27985 8375 28043 8381
rect 11422 8304 11428 8356
rect 11480 8344 11486 8356
rect 11701 8347 11759 8353
rect 11701 8344 11713 8347
rect 11480 8316 11713 8344
rect 11480 8304 11486 8316
rect 11701 8313 11713 8316
rect 11747 8344 11759 8347
rect 12176 8344 12204 8372
rect 11747 8316 12204 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 12268 8285 12296 8372
rect 14277 8347 14335 8353
rect 14277 8313 14289 8347
rect 14323 8344 14335 8347
rect 14918 8344 14924 8356
rect 14323 8316 14924 8344
rect 14323 8313 14335 8316
rect 14277 8307 14335 8313
rect 14918 8304 14924 8316
rect 14976 8344 14982 8356
rect 16758 8344 16764 8356
rect 14976 8316 16764 8344
rect 14976 8304 14982 8316
rect 16758 8304 16764 8316
rect 16816 8344 16822 8356
rect 19628 8344 19656 8372
rect 16816 8316 19656 8344
rect 16816 8304 16822 8316
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 26418 8344 26424 8356
rect 23440 8316 26424 8344
rect 23440 8304 23446 8316
rect 26418 8304 26424 8316
rect 26476 8344 26482 8356
rect 26476 8316 27384 8344
rect 26476 8304 26482 8316
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8245 12311 8279
rect 12253 8239 12311 8245
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 22278 8276 22284 8288
rect 17460 8248 22284 8276
rect 17460 8236 17466 8248
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 27356 8276 27384 8316
rect 27430 8304 27436 8356
rect 27488 8344 27494 8356
rect 28721 8347 28779 8353
rect 28721 8344 28733 8347
rect 27488 8316 28733 8344
rect 27488 8304 27494 8316
rect 28721 8313 28733 8316
rect 28767 8313 28779 8347
rect 29733 8347 29791 8353
rect 29733 8344 29745 8347
rect 28721 8307 28779 8313
rect 28828 8316 29745 8344
rect 28828 8276 28856 8316
rect 29733 8313 29745 8316
rect 29779 8313 29791 8347
rect 29840 8344 29868 8384
rect 30745 8381 30757 8415
rect 30791 8381 30803 8415
rect 30852 8412 30880 8440
rect 31128 8412 31156 8443
rect 31570 8440 31576 8452
rect 31628 8440 31634 8492
rect 31726 8483 31760 8492
rect 31726 8452 31739 8483
rect 31727 8449 31739 8452
rect 31727 8443 31760 8449
rect 31754 8440 31760 8443
rect 31812 8440 31818 8492
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8480 33471 8483
rect 40313 8483 40371 8489
rect 33459 8452 33824 8480
rect 33459 8449 33471 8452
rect 33413 8443 33471 8449
rect 33796 8421 33824 8452
rect 40313 8449 40325 8483
rect 40359 8480 40371 8483
rect 40402 8480 40408 8492
rect 40359 8452 40408 8480
rect 40359 8449 40371 8452
rect 40313 8443 40371 8449
rect 40402 8440 40408 8452
rect 40460 8440 40466 8492
rect 40512 8489 40540 8520
rect 41049 8517 41061 8520
rect 41095 8517 41107 8551
rect 41049 8511 41107 8517
rect 41690 8508 41696 8560
rect 41748 8548 41754 8560
rect 41877 8551 41935 8557
rect 41877 8548 41889 8551
rect 41748 8520 41889 8548
rect 41748 8508 41754 8520
rect 41877 8517 41889 8520
rect 41923 8517 41935 8551
rect 41877 8511 41935 8517
rect 41966 8508 41972 8560
rect 42024 8548 42030 8560
rect 42077 8551 42135 8557
rect 42077 8548 42089 8551
rect 42024 8520 42089 8548
rect 42024 8508 42030 8520
rect 42077 8517 42089 8520
rect 42123 8517 42135 8551
rect 42077 8511 42135 8517
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8449 40555 8483
rect 40497 8443 40555 8449
rect 40586 8440 40592 8492
rect 40644 8440 40650 8492
rect 30852 8384 31156 8412
rect 33781 8415 33839 8421
rect 30745 8375 30803 8381
rect 33781 8381 33793 8415
rect 33827 8381 33839 8415
rect 33781 8375 33839 8381
rect 30760 8344 30788 8375
rect 41414 8372 41420 8424
rect 41472 8412 41478 8424
rect 41601 8415 41659 8421
rect 41601 8412 41613 8415
rect 41472 8384 41613 8412
rect 41472 8372 41478 8384
rect 41601 8381 41613 8384
rect 41647 8381 41659 8415
rect 41601 8375 41659 8381
rect 42981 8415 43039 8421
rect 42981 8381 42993 8415
rect 43027 8381 43039 8415
rect 42981 8375 43039 8381
rect 31662 8344 31668 8356
rect 29840 8316 31668 8344
rect 29733 8307 29791 8313
rect 31662 8304 31668 8316
rect 31720 8304 31726 8356
rect 33965 8347 34023 8353
rect 33965 8313 33977 8347
rect 34011 8344 34023 8347
rect 34238 8344 34244 8356
rect 34011 8316 34244 8344
rect 34011 8313 34023 8316
rect 33965 8307 34023 8313
rect 34238 8304 34244 8316
rect 34296 8304 34302 8356
rect 42996 8344 43024 8375
rect 43714 8372 43720 8424
rect 43772 8372 43778 8424
rect 42168 8316 43024 8344
rect 27356 8248 28856 8276
rect 30466 8236 30472 8288
rect 30524 8236 30530 8288
rect 31478 8236 31484 8288
rect 31536 8236 31542 8288
rect 33594 8236 33600 8288
rect 33652 8236 33658 8288
rect 35897 8279 35955 8285
rect 35897 8245 35909 8279
rect 35943 8276 35955 8279
rect 36354 8276 36360 8288
rect 35943 8248 36360 8276
rect 35943 8245 35955 8248
rect 35897 8239 35955 8245
rect 36354 8236 36360 8248
rect 36412 8236 36418 8288
rect 40310 8236 40316 8288
rect 40368 8236 40374 8288
rect 40773 8279 40831 8285
rect 40773 8245 40785 8279
rect 40819 8276 40831 8279
rect 41230 8276 41236 8288
rect 40819 8248 41236 8276
rect 40819 8245 40831 8248
rect 40773 8239 40831 8245
rect 41230 8236 41236 8248
rect 41288 8236 41294 8288
rect 42058 8236 42064 8288
rect 42116 8276 42122 8288
rect 42168 8276 42196 8316
rect 42116 8248 42196 8276
rect 42116 8236 42122 8248
rect 42426 8236 42432 8288
rect 42484 8236 42490 8288
rect 1104 8186 45172 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 45172 8186
rect 1104 8112 45172 8134
rect 11698 8032 11704 8084
rect 11756 8032 11762 8084
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12066 8072 12072 8084
rect 12023 8044 12072 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12544 8044 13032 8072
rect 12544 8004 12572 8044
rect 11624 7976 12572 8004
rect 11624 7948 11652 7976
rect 12618 7964 12624 8016
rect 12676 7964 12682 8016
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12268 7908 12357 7936
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11808 7840 12173 7868
rect 11808 7812 11836 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 11790 7760 11796 7812
rect 11848 7760 11854 7812
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 12268 7800 12296 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7905 12495 7939
rect 13004 7936 13032 8044
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13722 8072 13728 8084
rect 13320 8044 13728 8072
rect 13320 8032 13326 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19518 8072 19524 8084
rect 18840 8044 19524 8072
rect 18840 8032 18846 8044
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 20070 8032 20076 8084
rect 20128 8072 20134 8084
rect 20128 8044 20300 8072
rect 20128 8032 20134 8044
rect 19610 7964 19616 8016
rect 19668 8004 19674 8016
rect 19668 7976 20208 8004
rect 19668 7964 19674 7976
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 13004 7908 13093 7936
rect 12437 7899 12495 7905
rect 13081 7905 13093 7908
rect 13127 7936 13139 7939
rect 13262 7936 13268 7948
rect 13127 7908 13268 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 12452 7870 12480 7899
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 15470 7896 15476 7948
rect 15528 7936 15534 7948
rect 19337 7939 19395 7945
rect 19337 7936 19349 7939
rect 15528 7908 19349 7936
rect 15528 7896 15534 7908
rect 19337 7905 19349 7908
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 19426 7896 19432 7948
rect 19484 7936 19490 7948
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 19484 7908 19809 7936
rect 19484 7896 19490 7908
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 19886 7896 19892 7948
rect 19944 7896 19950 7948
rect 12032 7772 12296 7800
rect 12360 7842 12480 7870
rect 12360 7800 12388 7842
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12728 7800 12756 7828
rect 12360 7772 12756 7800
rect 12912 7800 12940 7831
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 16632 7840 17601 7868
rect 16632 7828 16638 7840
rect 17589 7837 17601 7840
rect 17635 7868 17647 7871
rect 17678 7868 17684 7880
rect 17635 7840 17684 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 18138 7868 18144 7880
rect 17819 7840 18144 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 13170 7800 13176 7812
rect 12912 7772 13176 7800
rect 12032 7760 12038 7772
rect 13170 7760 13176 7772
rect 13228 7800 13234 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 13228 7772 13277 7800
rect 13228 7760 13234 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 17788 7800 17816 7831
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 18892 7840 19717 7868
rect 13265 7763 13323 7769
rect 14844 7772 17816 7800
rect 14844 7744 14872 7772
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 12250 7732 12256 7744
rect 11296 7704 12256 7732
rect 11296 7692 11302 7704
rect 12250 7692 12256 7704
rect 12308 7732 12314 7744
rect 13357 7735 13415 7741
rect 13357 7732 13369 7735
rect 12308 7704 13369 7732
rect 12308 7692 12314 7704
rect 13357 7701 13369 7704
rect 13403 7701 13415 7735
rect 13357 7695 13415 7701
rect 14826 7692 14832 7744
rect 14884 7692 14890 7744
rect 17678 7692 17684 7744
rect 17736 7692 17742 7744
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18892 7732 18920 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19904 7868 19932 7896
rect 20180 7877 20208 7976
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19904 7840 20085 7868
rect 19705 7831 19763 7837
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20272 7868 20300 8044
rect 21818 8032 21824 8084
rect 21876 8032 21882 8084
rect 23290 8032 23296 8084
rect 23348 8032 23354 8084
rect 23934 8032 23940 8084
rect 23992 8032 23998 8084
rect 25590 8032 25596 8084
rect 25648 8032 25654 8084
rect 26694 8032 26700 8084
rect 26752 8032 26758 8084
rect 27525 8075 27583 8081
rect 27525 8072 27537 8075
rect 26804 8044 27537 8072
rect 25608 8004 25636 8032
rect 26804 8004 26832 8044
rect 27525 8041 27537 8044
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 29730 8032 29736 8084
rect 29788 8072 29794 8084
rect 30190 8072 30196 8084
rect 29788 8044 30196 8072
rect 29788 8032 29794 8044
rect 30190 8032 30196 8044
rect 30248 8032 30254 8084
rect 31018 8032 31024 8084
rect 31076 8072 31082 8084
rect 31205 8075 31263 8081
rect 31205 8072 31217 8075
rect 31076 8044 31217 8072
rect 31076 8032 31082 8044
rect 31205 8041 31217 8044
rect 31251 8041 31263 8075
rect 40310 8072 40316 8084
rect 31205 8035 31263 8041
rect 39684 8044 40316 8072
rect 27338 8004 27344 8016
rect 25608 7976 26832 8004
rect 27080 7976 27344 8004
rect 20349 7871 20407 7877
rect 20349 7868 20361 7871
rect 20272 7840 20361 7868
rect 20165 7831 20223 7837
rect 20349 7837 20361 7840
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 19334 7760 19340 7812
rect 19392 7760 19398 7812
rect 18380 7704 18920 7732
rect 19352 7732 19380 7760
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19352 7704 19441 7732
rect 18380 7692 18386 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 19518 7692 19524 7744
rect 19576 7692 19582 7744
rect 19720 7732 19748 7831
rect 20438 7828 20444 7880
rect 20496 7828 20502 7880
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 22094 7868 22100 7880
rect 21683 7840 22100 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 27080 7877 27108 7976
rect 27338 7964 27344 7976
rect 27396 8004 27402 8016
rect 28353 8007 28411 8013
rect 28353 8004 28365 8007
rect 27396 7976 28365 8004
rect 27396 7964 27402 7976
rect 28353 7973 28365 7976
rect 28399 7973 28411 8007
rect 28353 7967 28411 7973
rect 36449 8007 36507 8013
rect 36449 7973 36461 8007
rect 36495 8004 36507 8007
rect 36630 8004 36636 8016
rect 36495 7976 36636 8004
rect 36495 7973 36507 7976
rect 36449 7967 36507 7973
rect 36630 7964 36636 7976
rect 36688 8004 36694 8016
rect 37001 8007 37059 8013
rect 37001 8004 37013 8007
rect 36688 7976 37013 8004
rect 36688 7964 36694 7976
rect 37001 7973 37013 7976
rect 37047 7973 37059 8007
rect 37001 7967 37059 7973
rect 27249 7939 27307 7945
rect 27249 7905 27261 7939
rect 27295 7936 27307 7939
rect 27522 7936 27528 7948
rect 27295 7908 27528 7936
rect 27295 7905 27307 7908
rect 27249 7899 27307 7905
rect 27522 7896 27528 7908
rect 27580 7936 27586 7948
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 27580 7908 28089 7936
rect 27580 7896 27586 7908
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28077 7899 28135 7905
rect 28721 7939 28779 7945
rect 28721 7905 28733 7939
rect 28767 7936 28779 7939
rect 29086 7936 29092 7948
rect 28767 7908 29092 7936
rect 28767 7905 28779 7908
rect 28721 7899 28779 7905
rect 29086 7896 29092 7908
rect 29144 7936 29150 7948
rect 29144 7908 29960 7936
rect 29144 7896 29150 7908
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 27065 7871 27123 7877
rect 24075 7840 24440 7868
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 19981 7803 20039 7809
rect 19981 7769 19993 7803
rect 20027 7800 20039 7803
rect 20456 7800 20484 7828
rect 20027 7772 20484 7800
rect 20027 7769 20039 7772
rect 19981 7763 20039 7769
rect 21450 7760 21456 7812
rect 21508 7760 21514 7812
rect 21542 7760 21548 7812
rect 21600 7800 21606 7812
rect 22005 7803 22063 7809
rect 22005 7800 22017 7803
rect 21600 7772 22017 7800
rect 21600 7760 21606 7772
rect 22005 7769 22017 7772
rect 22051 7769 22063 7803
rect 22005 7763 22063 7769
rect 24412 7744 24440 7840
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27890 7828 27896 7880
rect 27948 7828 27954 7880
rect 28534 7828 28540 7880
rect 28592 7828 28598 7880
rect 27157 7803 27215 7809
rect 27157 7769 27169 7803
rect 27203 7800 27215 7803
rect 27338 7800 27344 7812
rect 27203 7772 27344 7800
rect 27203 7769 27215 7772
rect 27157 7763 27215 7769
rect 27338 7760 27344 7772
rect 27396 7800 27402 7812
rect 29932 7809 29960 7908
rect 34698 7896 34704 7948
rect 34756 7896 34762 7948
rect 36832 7908 37136 7936
rect 31113 7871 31171 7877
rect 31113 7837 31125 7871
rect 31159 7837 31171 7871
rect 31113 7831 31171 7837
rect 31297 7871 31355 7877
rect 31297 7837 31309 7871
rect 31343 7868 31355 7871
rect 31478 7868 31484 7880
rect 31343 7840 31484 7868
rect 31343 7837 31355 7840
rect 31297 7831 31355 7837
rect 29917 7803 29975 7809
rect 27396 7772 29592 7800
rect 27396 7760 27402 7772
rect 20346 7732 20352 7744
rect 19720 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 24394 7692 24400 7744
rect 24452 7692 24458 7744
rect 27985 7735 28043 7741
rect 27985 7701 27997 7735
rect 28031 7732 28043 7735
rect 28074 7732 28080 7744
rect 28031 7704 28080 7732
rect 28031 7701 28043 7704
rect 27985 7695 28043 7701
rect 28074 7692 28080 7704
rect 28132 7692 28138 7744
rect 29564 7741 29592 7772
rect 29917 7769 29929 7803
rect 29963 7769 29975 7803
rect 29917 7763 29975 7769
rect 30466 7760 30472 7812
rect 30524 7760 30530 7812
rect 31128 7800 31156 7831
rect 31478 7828 31484 7840
rect 31536 7828 31542 7880
rect 31570 7828 31576 7880
rect 31628 7828 31634 7880
rect 36541 7871 36599 7877
rect 36541 7837 36553 7871
rect 36587 7837 36599 7871
rect 36541 7831 36599 7837
rect 31588 7800 31616 7828
rect 31128 7772 31616 7800
rect 34974 7760 34980 7812
rect 35032 7760 35038 7812
rect 36354 7800 36360 7812
rect 36202 7772 36360 7800
rect 36354 7760 36360 7772
rect 36412 7760 36418 7812
rect 29549 7735 29607 7741
rect 29549 7701 29561 7735
rect 29595 7701 29607 7735
rect 29549 7695 29607 7701
rect 29717 7735 29775 7741
rect 29717 7701 29729 7735
rect 29763 7732 29775 7735
rect 30484 7732 30512 7760
rect 36556 7744 36584 7831
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 36832 7877 36860 7908
rect 36817 7871 36875 7877
rect 36817 7837 36829 7871
rect 36863 7837 36875 7871
rect 36817 7831 36875 7837
rect 36906 7828 36912 7880
rect 36964 7828 36970 7880
rect 36924 7800 36952 7828
rect 37108 7812 37136 7908
rect 37752 7908 39528 7936
rect 37752 7880 37780 7908
rect 37734 7828 37740 7880
rect 37792 7828 37798 7880
rect 39298 7828 39304 7880
rect 39356 7828 39362 7880
rect 39500 7877 39528 7908
rect 39684 7877 39712 8044
rect 40310 8032 40316 8044
rect 40368 8032 40374 8084
rect 41877 8075 41935 8081
rect 41877 8041 41889 8075
rect 41923 8072 41935 8075
rect 42058 8072 42064 8084
rect 41923 8044 42064 8072
rect 41923 8041 41935 8044
rect 41877 8035 41935 8041
rect 42058 8032 42064 8044
rect 42116 8032 42122 8084
rect 39853 7939 39911 7945
rect 39853 7905 39865 7939
rect 39899 7936 39911 7939
rect 39899 7908 43668 7936
rect 39899 7905 39911 7908
rect 39853 7899 39911 7905
rect 43640 7880 43668 7908
rect 39485 7871 39543 7877
rect 39485 7837 39497 7871
rect 39531 7837 39543 7871
rect 39485 7831 39543 7837
rect 39669 7871 39727 7877
rect 39669 7837 39681 7871
rect 39715 7837 39727 7871
rect 39669 7831 39727 7837
rect 37001 7803 37059 7809
rect 37001 7800 37013 7803
rect 36924 7772 37013 7800
rect 37001 7769 37013 7772
rect 37047 7769 37059 7803
rect 37001 7763 37059 7769
rect 37090 7760 37096 7812
rect 37148 7760 37154 7812
rect 38654 7760 38660 7812
rect 38712 7800 38718 7812
rect 38712 7772 39160 7800
rect 38712 7760 38718 7772
rect 29763 7704 30512 7732
rect 29763 7701 29775 7704
rect 29717 7695 29775 7701
rect 36538 7692 36544 7744
rect 36596 7692 36602 7744
rect 36814 7692 36820 7744
rect 36872 7692 36878 7744
rect 37458 7692 37464 7744
rect 37516 7692 37522 7744
rect 37550 7692 37556 7744
rect 37608 7692 37614 7744
rect 37737 7735 37795 7741
rect 37737 7701 37749 7735
rect 37783 7732 37795 7735
rect 38746 7732 38752 7744
rect 37783 7704 38752 7732
rect 37783 7701 37795 7704
rect 37737 7695 37795 7701
rect 38746 7692 38752 7704
rect 38804 7692 38810 7744
rect 39132 7741 39160 7772
rect 39117 7735 39175 7741
rect 39117 7701 39129 7735
rect 39163 7701 39175 7735
rect 39500 7732 39528 7831
rect 41230 7828 41236 7880
rect 41288 7868 41294 7880
rect 41288 7854 42274 7868
rect 41288 7840 42288 7854
rect 41288 7828 41294 7840
rect 39577 7803 39635 7809
rect 39577 7769 39589 7803
rect 39623 7800 39635 7803
rect 40129 7803 40187 7809
rect 40129 7800 40141 7803
rect 39623 7772 40141 7800
rect 39623 7769 39635 7772
rect 39577 7763 39635 7769
rect 40129 7769 40141 7772
rect 40175 7769 40187 7803
rect 40129 7763 40187 7769
rect 40218 7732 40224 7744
rect 39500 7704 40224 7732
rect 39117 7695 39175 7701
rect 40218 7692 40224 7704
rect 40276 7692 40282 7744
rect 41414 7692 41420 7744
rect 41472 7732 41478 7744
rect 41601 7735 41659 7741
rect 41601 7732 41613 7735
rect 41472 7704 41613 7732
rect 41472 7692 41478 7704
rect 41601 7701 41613 7704
rect 41647 7701 41659 7735
rect 42260 7732 42288 7840
rect 43622 7828 43628 7880
rect 43680 7828 43686 7880
rect 42918 7772 43024 7800
rect 42996 7732 43024 7772
rect 43070 7760 43076 7812
rect 43128 7800 43134 7812
rect 43349 7803 43407 7809
rect 43349 7800 43361 7803
rect 43128 7772 43361 7800
rect 43128 7760 43134 7772
rect 43349 7769 43361 7772
rect 43395 7769 43407 7803
rect 43349 7763 43407 7769
rect 43438 7760 43444 7812
rect 43496 7760 43502 7812
rect 43456 7732 43484 7760
rect 42260 7704 43484 7732
rect 41601 7695 41659 7701
rect 1104 7642 45172 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 45172 7642
rect 1104 7568 45172 7590
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 12526 7528 12532 7540
rect 12124 7500 12532 7528
rect 12124 7488 12130 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13262 7488 13268 7540
rect 13320 7537 13326 7540
rect 13320 7531 13344 7537
rect 13332 7497 13344 7531
rect 13320 7491 13344 7497
rect 13320 7488 13326 7491
rect 13722 7488 13728 7540
rect 13780 7488 13786 7540
rect 14200 7500 14780 7528
rect 11149 7463 11207 7469
rect 11149 7429 11161 7463
rect 11195 7460 11207 7463
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 11195 7432 11805 7460
rect 11195 7429 11207 7432
rect 11149 7423 11207 7429
rect 11793 7429 11805 7432
rect 11839 7460 11851 7463
rect 12345 7463 12403 7469
rect 12345 7460 12357 7463
rect 11839 7432 12357 7460
rect 11839 7429 11851 7432
rect 11793 7423 11851 7429
rect 12345 7429 12357 7432
rect 12391 7429 12403 7463
rect 12345 7423 12403 7429
rect 13078 7420 13084 7472
rect 13136 7420 13142 7472
rect 14200 7460 14228 7500
rect 13372 7432 14228 7460
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 11698 7392 11704 7404
rect 11379 7364 11704 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 6914 7284 6920 7336
rect 6972 7284 6978 7336
rect 11072 7256 11100 7355
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12250 7392 12256 7404
rect 12207 7364 12256 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 13372 7392 13400 7432
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 14645 7463 14703 7469
rect 14645 7460 14657 7463
rect 14332 7432 14657 7460
rect 14332 7420 14338 7432
rect 14645 7429 14657 7432
rect 14691 7429 14703 7463
rect 14752 7460 14780 7500
rect 14826 7488 14832 7540
rect 14884 7488 14890 7540
rect 15470 7488 15476 7540
rect 15528 7488 15534 7540
rect 17402 7488 17408 7540
rect 17460 7488 17466 7540
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 18616 7500 19533 7528
rect 15746 7460 15752 7472
rect 14752 7432 15752 7460
rect 14645 7423 14703 7429
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 17696 7460 17724 7488
rect 17696 7432 18460 7460
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 12759 7364 13400 7392
rect 13464 7364 13553 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 13354 7256 13360 7268
rect 11072 7228 13360 7256
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 13464 7265 13492 7364
rect 13541 7361 13553 7364
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 14734 7352 14740 7404
rect 14792 7352 14798 7404
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 14976 7364 15301 7392
rect 14976 7352 14982 7364
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 16991 7364 17509 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 13449 7259 13507 7265
rect 13449 7225 13461 7259
rect 13495 7225 13507 7259
rect 14476 7256 14504 7352
rect 14752 7324 14780 7352
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14752 7296 15117 7324
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 17034 7284 17040 7336
rect 17092 7284 17098 7336
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 14826 7256 14832 7268
rect 14476 7228 14832 7256
rect 13449 7219 13507 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 17144 7256 17172 7287
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 17696 7324 17724 7355
rect 17954 7352 17960 7404
rect 18012 7352 18018 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18322 7392 18328 7404
rect 18187 7364 18328 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18432 7401 18460 7432
rect 18616 7401 18644 7500
rect 19521 7497 19533 7500
rect 19567 7528 19579 7531
rect 19978 7528 19984 7540
rect 19567 7500 19984 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19245 7463 19303 7469
rect 19245 7460 19257 7463
rect 19024 7432 19257 7460
rect 19024 7420 19030 7432
rect 19245 7429 19257 7432
rect 19291 7460 19303 7463
rect 19334 7460 19340 7472
rect 19291 7432 19340 7460
rect 19291 7429 19303 7432
rect 19245 7423 19303 7429
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 19812 7469 19840 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 24578 7528 24584 7540
rect 23216 7500 24584 7528
rect 19797 7463 19855 7469
rect 19797 7429 19809 7463
rect 19843 7460 19855 7463
rect 20165 7463 20223 7469
rect 19843 7432 19877 7460
rect 19843 7429 19855 7432
rect 19797 7423 19855 7429
rect 20165 7429 20177 7463
rect 20211 7460 20223 7463
rect 20346 7460 20352 7472
rect 20211 7432 20352 7460
rect 20211 7429 20223 7432
rect 20165 7423 20223 7429
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 20254 7352 20260 7404
rect 20312 7352 20318 7404
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 17696 7296 18245 7324
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7324 18751 7327
rect 19978 7324 19984 7336
rect 18739 7296 19984 7324
rect 18739 7293 18751 7296
rect 18693 7287 18751 7293
rect 17954 7256 17960 7268
rect 17144 7228 17960 7256
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 11330 7148 11336 7200
rect 11388 7148 11394 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 13228 7160 13277 7188
rect 13228 7148 13234 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16298 7188 16304 7200
rect 15804 7160 16304 7188
rect 15804 7148 15810 7160
rect 16298 7148 16304 7160
rect 16356 7188 16362 7200
rect 18524 7188 18552 7287
rect 19978 7284 19984 7296
rect 20036 7324 20042 7336
rect 20272 7324 20300 7352
rect 20036 7296 20300 7324
rect 20548 7324 20576 7488
rect 22005 7463 22063 7469
rect 22005 7429 22017 7463
rect 22051 7460 22063 7463
rect 23216 7460 23244 7500
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 24857 7531 24915 7537
rect 24857 7497 24869 7531
rect 24903 7528 24915 7531
rect 25314 7528 25320 7540
rect 24903 7500 25320 7528
rect 24903 7497 24915 7500
rect 24857 7491 24915 7497
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 26878 7488 26884 7540
rect 26936 7528 26942 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 26936 7500 26985 7528
rect 26936 7488 26942 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 27338 7488 27344 7540
rect 27396 7488 27402 7540
rect 27433 7531 27491 7537
rect 27433 7497 27445 7531
rect 27479 7528 27491 7531
rect 27890 7528 27896 7540
rect 27479 7500 27896 7528
rect 27479 7497 27491 7500
rect 27433 7491 27491 7497
rect 27890 7488 27896 7500
rect 27948 7488 27954 7540
rect 34974 7488 34980 7540
rect 35032 7488 35038 7540
rect 36630 7488 36636 7540
rect 36688 7488 36694 7540
rect 36722 7488 36728 7540
rect 36780 7528 36786 7540
rect 37001 7531 37059 7537
rect 37001 7528 37013 7531
rect 36780 7500 37013 7528
rect 36780 7488 36786 7500
rect 37001 7497 37013 7500
rect 37047 7497 37059 7531
rect 37001 7491 37059 7497
rect 37274 7488 37280 7540
rect 37332 7528 37338 7540
rect 37332 7500 41414 7528
rect 37332 7488 37338 7500
rect 22051 7432 23244 7460
rect 22051 7429 22063 7432
rect 22005 7423 22063 7429
rect 23842 7420 23848 7472
rect 23900 7420 23906 7472
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21177 7355 21235 7361
rect 21560 7364 21925 7392
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20548 7296 20913 7324
rect 20036 7284 20042 7296
rect 20272 7256 20300 7296
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 21082 7284 21088 7336
rect 21140 7284 21146 7336
rect 21192 7268 21220 7355
rect 21174 7256 21180 7268
rect 20272 7228 21180 7256
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 21560 7265 21588 7364
rect 21913 7361 21925 7364
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 23860 7392 23888 7420
rect 23523 7364 23888 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 24854 7352 24860 7404
rect 24912 7352 24918 7404
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7392 25559 7395
rect 25958 7392 25964 7404
rect 25547 7364 25964 7392
rect 25547 7361 25559 7364
rect 25501 7355 25559 7361
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7324 23259 7327
rect 23566 7324 23572 7336
rect 23247 7296 23572 7324
rect 23247 7293 23259 7296
rect 23201 7287 23259 7293
rect 23566 7284 23572 7296
rect 23624 7324 23630 7336
rect 24394 7324 24400 7336
rect 23624 7296 24400 7324
rect 23624 7284 23630 7296
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 25777 7327 25835 7333
rect 25777 7293 25789 7327
rect 25823 7324 25835 7327
rect 25866 7324 25872 7336
rect 25823 7296 25872 7324
rect 25823 7293 25835 7296
rect 25777 7287 25835 7293
rect 25866 7284 25872 7296
rect 25924 7284 25930 7336
rect 27522 7284 27528 7336
rect 27580 7284 27586 7336
rect 34992 7324 35020 7488
rect 35805 7395 35863 7401
rect 35805 7361 35817 7395
rect 35851 7392 35863 7395
rect 36173 7395 36231 7401
rect 36173 7392 36185 7395
rect 35851 7364 36185 7392
rect 35851 7361 35863 7364
rect 35805 7355 35863 7361
rect 36173 7361 36185 7364
rect 36219 7361 36231 7395
rect 36648 7392 36676 7488
rect 37016 7432 37582 7460
rect 37016 7404 37044 7432
rect 38746 7420 38752 7472
rect 38804 7460 38810 7472
rect 39206 7460 39212 7472
rect 38804 7432 39212 7460
rect 38804 7420 38810 7432
rect 39206 7420 39212 7432
rect 39264 7460 39270 7472
rect 39264 7432 39344 7460
rect 39264 7420 39270 7432
rect 36725 7395 36783 7401
rect 36725 7392 36737 7395
rect 36648 7364 36737 7392
rect 36173 7355 36231 7361
rect 36725 7361 36737 7364
rect 36771 7361 36783 7395
rect 36725 7355 36783 7361
rect 35437 7327 35495 7333
rect 35437 7324 35449 7327
rect 34992 7296 35449 7324
rect 35437 7293 35449 7296
rect 35483 7293 35495 7327
rect 35437 7287 35495 7293
rect 35897 7327 35955 7333
rect 35897 7293 35909 7327
rect 35943 7293 35955 7327
rect 35897 7287 35955 7293
rect 21545 7259 21603 7265
rect 21545 7225 21557 7259
rect 21591 7225 21603 7259
rect 21545 7219 21603 7225
rect 16356 7160 18552 7188
rect 16356 7148 16362 7160
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20220 7160 20453 7188
rect 20220 7148 20226 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20441 7151 20499 7157
rect 23382 7148 23388 7200
rect 23440 7148 23446 7200
rect 35912 7188 35940 7287
rect 36740 7256 36768 7355
rect 36906 7352 36912 7404
rect 36964 7352 36970 7404
rect 36998 7352 37004 7404
rect 37056 7352 37062 7404
rect 37093 7395 37151 7401
rect 37093 7361 37105 7395
rect 37139 7392 37151 7395
rect 37366 7392 37372 7404
rect 37139 7364 37372 7392
rect 37139 7361 37151 7364
rect 37093 7355 37151 7361
rect 37366 7352 37372 7364
rect 37424 7352 37430 7404
rect 39114 7352 39120 7404
rect 39172 7352 39178 7404
rect 39316 7401 39344 7432
rect 39592 7432 39988 7460
rect 39592 7404 39620 7432
rect 39301 7395 39359 7401
rect 39301 7361 39313 7395
rect 39347 7361 39359 7395
rect 39301 7355 39359 7361
rect 39574 7352 39580 7404
rect 39632 7352 39638 7404
rect 39960 7401 39988 7432
rect 40218 7420 40224 7472
rect 40276 7420 40282 7472
rect 41386 7460 41414 7500
rect 41690 7488 41696 7540
rect 41748 7528 41754 7540
rect 42242 7528 42248 7540
rect 41748 7500 42248 7528
rect 41748 7488 41754 7500
rect 42242 7488 42248 7500
rect 42300 7528 42306 7540
rect 42613 7531 42671 7537
rect 42613 7528 42625 7531
rect 42300 7500 42625 7528
rect 42300 7488 42306 7500
rect 42613 7497 42625 7500
rect 42659 7497 42671 7531
rect 42613 7491 42671 7497
rect 43622 7488 43628 7540
rect 43680 7528 43686 7540
rect 44269 7531 44327 7537
rect 44269 7528 44281 7531
rect 43680 7500 44281 7528
rect 43680 7488 43686 7500
rect 44269 7497 44281 7500
rect 44315 7497 44327 7531
rect 44269 7491 44327 7497
rect 42981 7463 43039 7469
rect 42981 7460 42993 7463
rect 41386 7432 42993 7460
rect 42981 7429 42993 7432
rect 43027 7429 43039 7463
rect 42981 7423 43039 7429
rect 39669 7395 39727 7401
rect 39669 7361 39681 7395
rect 39715 7361 39727 7395
rect 39669 7355 39727 7361
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 37277 7327 37335 7333
rect 37277 7293 37289 7327
rect 37323 7324 37335 7327
rect 37550 7324 37556 7336
rect 37323 7296 37556 7324
rect 37323 7293 37335 7296
rect 37277 7287 37335 7293
rect 37550 7284 37556 7296
rect 37608 7284 37614 7336
rect 38746 7284 38752 7336
rect 38804 7284 38810 7336
rect 39022 7284 39028 7336
rect 39080 7284 39086 7336
rect 39684 7268 39712 7355
rect 40402 7352 40408 7404
rect 40460 7352 40466 7404
rect 41322 7352 41328 7404
rect 41380 7352 41386 7404
rect 41509 7395 41567 7401
rect 41509 7361 41521 7395
rect 41555 7392 41567 7395
rect 41555 7364 41644 7392
rect 41555 7361 41567 7364
rect 41509 7355 41567 7361
rect 40589 7327 40647 7333
rect 40589 7293 40601 7327
rect 40635 7324 40647 7327
rect 41414 7324 41420 7336
rect 40635 7296 41420 7324
rect 40635 7293 40647 7296
rect 40589 7287 40647 7293
rect 41414 7284 41420 7296
rect 41472 7284 41478 7336
rect 37642 7256 37648 7268
rect 36740 7228 37648 7256
rect 37642 7216 37648 7228
rect 37700 7216 37706 7268
rect 39666 7216 39672 7268
rect 39724 7256 39730 7268
rect 41325 7259 41383 7265
rect 41325 7256 41337 7259
rect 39724 7228 41337 7256
rect 39724 7216 39730 7228
rect 41325 7225 41337 7228
rect 41371 7225 41383 7259
rect 41325 7219 41383 7225
rect 37734 7188 37740 7200
rect 35912 7160 37740 7188
rect 37734 7148 37740 7160
rect 37792 7148 37798 7200
rect 39482 7148 39488 7200
rect 39540 7188 39546 7200
rect 39577 7191 39635 7197
rect 39577 7188 39589 7191
rect 39540 7160 39589 7188
rect 39540 7148 39546 7160
rect 39577 7157 39589 7160
rect 39623 7157 39635 7191
rect 41432 7188 41460 7284
rect 41616 7265 41644 7364
rect 41782 7352 41788 7404
rect 41840 7352 41846 7404
rect 41969 7395 42027 7401
rect 41969 7361 41981 7395
rect 42015 7392 42027 7395
rect 42058 7392 42064 7404
rect 42015 7364 42064 7392
rect 42015 7361 42027 7364
rect 41969 7355 42027 7361
rect 42058 7352 42064 7364
rect 42116 7352 42122 7404
rect 42242 7352 42248 7404
rect 42300 7352 42306 7404
rect 42426 7352 42432 7404
rect 42484 7352 42490 7404
rect 42702 7352 42708 7404
rect 42760 7352 42766 7404
rect 41601 7259 41659 7265
rect 41601 7225 41613 7259
rect 41647 7225 41659 7259
rect 41601 7219 41659 7225
rect 42429 7259 42487 7265
rect 42429 7225 42441 7259
rect 42475 7256 42487 7259
rect 43714 7256 43720 7268
rect 42475 7228 43720 7256
rect 42475 7225 42487 7228
rect 42429 7219 42487 7225
rect 43714 7216 43720 7228
rect 43772 7216 43778 7268
rect 41785 7191 41843 7197
rect 41785 7188 41797 7191
rect 41432 7160 41797 7188
rect 39577 7151 39635 7157
rect 41785 7157 41797 7160
rect 41831 7157 41843 7191
rect 41785 7151 41843 7157
rect 1104 7098 45172 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 45172 7098
rect 1104 7024 45172 7046
rect 6914 6944 6920 6996
rect 6972 6944 6978 6996
rect 7947 6987 8005 6993
rect 7947 6953 7959 6987
rect 7993 6984 8005 6987
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 7993 6956 8953 6984
rect 7993 6953 8005 6956
rect 7947 6947 8005 6953
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 11606 6944 11612 6996
rect 11664 6944 11670 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 11756 6956 12633 6984
rect 11756 6944 11762 6956
rect 12621 6953 12633 6956
rect 12667 6984 12679 6987
rect 15930 6984 15936 6996
rect 12667 6956 15936 6984
rect 12667 6953 12679 6956
rect 12621 6947 12679 6953
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 16025 6987 16083 6993
rect 16025 6953 16037 6987
rect 16071 6984 16083 6987
rect 17037 6987 17095 6993
rect 16071 6956 16712 6984
rect 16071 6953 16083 6956
rect 16025 6947 16083 6953
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 6932 6848 6960 6944
rect 11624 6916 11652 6944
rect 11624 6888 12020 6916
rect 6503 6820 6960 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 11882 6808 11888 6860
rect 11940 6808 11946 6860
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 9953 6783 10011 6789
rect 9953 6780 9965 6783
rect 9824 6752 9965 6780
rect 9824 6740 9830 6752
rect 9953 6749 9965 6752
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11992 6789 12020 6888
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 14369 6919 14427 6925
rect 14369 6916 14381 6919
rect 12768 6888 14381 6916
rect 12768 6876 12774 6888
rect 14369 6885 14381 6888
rect 14415 6916 14427 6919
rect 15010 6916 15016 6928
rect 14415 6888 15016 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 16209 6919 16267 6925
rect 16209 6885 16221 6919
rect 16255 6916 16267 6919
rect 16255 6888 16620 6916
rect 16255 6885 16267 6888
rect 16209 6879 16267 6885
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13228 6820 13553 6848
rect 13228 6808 13234 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 15194 6848 15200 6860
rect 13541 6811 13599 6817
rect 13648 6820 15200 6848
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11388 6752 11529 6780
rect 11388 6740 11394 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12158 6740 12164 6792
rect 12216 6740 12222 6792
rect 13648 6780 13676 6820
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 16022 6848 16028 6860
rect 15611 6820 16028 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 12268 6752 13676 6780
rect 7282 6672 7288 6724
rect 7340 6672 7346 6724
rect 11701 6715 11759 6721
rect 11701 6681 11713 6715
rect 11747 6712 11759 6715
rect 12268 6712 12296 6752
rect 14090 6740 14096 6792
rect 14148 6740 14154 6792
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14642 6740 14648 6792
rect 14700 6740 14706 6792
rect 14918 6740 14924 6792
rect 14976 6740 14982 6792
rect 15654 6780 15660 6792
rect 15212 6752 15660 6780
rect 11747 6684 12296 6712
rect 11747 6681 11759 6684
rect 11701 6675 11759 6681
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 12529 6715 12587 6721
rect 12529 6681 12541 6715
rect 12575 6681 12587 6715
rect 12529 6675 12587 6681
rect 13081 6715 13139 6721
rect 13081 6681 13093 6715
rect 13127 6712 13139 6715
rect 13725 6715 13783 6721
rect 13127 6684 13676 6712
rect 13127 6681 13139 6684
rect 13081 6675 13139 6681
rect 6362 6604 6368 6656
rect 6420 6604 6426 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9640 6616 9781 6644
rect 9640 6604 9646 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12250 6644 12256 6656
rect 11848 6616 12256 6644
rect 11848 6604 11854 6616
rect 12250 6604 12256 6616
rect 12308 6644 12314 6656
rect 12544 6644 12572 6675
rect 12308 6616 12572 6644
rect 13357 6647 13415 6653
rect 12308 6604 12314 6616
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13538 6644 13544 6656
rect 13403 6616 13544 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 13648 6644 13676 6684
rect 13725 6681 13737 6715
rect 13771 6712 13783 6715
rect 13814 6712 13820 6724
rect 13771 6684 13820 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 14384 6712 14412 6740
rect 14936 6712 14964 6740
rect 13955 6684 14964 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 15212 6644 15240 6752
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16206 6789 16212 6792
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16197 6783 16212 6789
rect 16197 6749 16209 6783
rect 16197 6743 16212 6749
rect 15856 6712 15884 6743
rect 16206 6740 16212 6743
rect 16264 6740 16270 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 15304 6684 15884 6712
rect 15304 6656 15332 6684
rect 13648 6616 15240 6644
rect 15286 6604 15292 6656
rect 15344 6604 15350 6656
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16408 6644 16436 6743
rect 16482 6740 16488 6792
rect 16540 6740 16546 6792
rect 16592 6789 16620 6888
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16684 6712 16712 6956
rect 17037 6953 17049 6987
rect 17083 6984 17095 6987
rect 17218 6984 17224 6996
rect 17083 6956 17224 6984
rect 17083 6953 17095 6956
rect 17037 6947 17095 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 17770 6984 17776 6996
rect 17451 6956 17776 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 17954 6944 17960 6996
rect 18012 6944 18018 6996
rect 18782 6944 18788 6996
rect 18840 6944 18846 6996
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 21269 6987 21327 6993
rect 21269 6984 21281 6987
rect 21140 6956 21281 6984
rect 21140 6944 21146 6956
rect 21269 6953 21281 6956
rect 21315 6953 21327 6987
rect 21269 6947 21327 6953
rect 21450 6944 21456 6996
rect 21508 6944 21514 6996
rect 23566 6944 23572 6996
rect 23624 6944 23630 6996
rect 23842 6944 23848 6996
rect 23900 6984 23906 6996
rect 24029 6987 24087 6993
rect 24029 6984 24041 6987
rect 23900 6956 24041 6984
rect 23900 6944 23906 6956
rect 24029 6953 24041 6956
rect 24075 6953 24087 6987
rect 25038 6984 25044 6996
rect 24029 6947 24087 6953
rect 24872 6956 25044 6984
rect 18800 6916 18828 6944
rect 16776 6888 16988 6916
rect 16776 6789 16804 6888
rect 16960 6848 16988 6888
rect 17788 6888 18828 6916
rect 19812 6888 20024 6916
rect 17788 6848 17816 6888
rect 16960 6820 17816 6848
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 19812 6848 19840 6888
rect 17911 6820 19840 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 19996 6848 20024 6888
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 19996 6820 20177 6848
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6848 21143 6851
rect 21468 6848 21496 6944
rect 23584 6916 23612 6944
rect 23032 6888 23612 6916
rect 23032 6857 23060 6888
rect 21131 6820 21496 6848
rect 23017 6851 23075 6857
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 23017 6817 23029 6851
rect 23063 6817 23075 6851
rect 23566 6848 23572 6860
rect 23017 6811 23075 6817
rect 23216 6820 23572 6848
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 16850 6740 16856 6792
rect 16908 6740 16914 6792
rect 17310 6740 17316 6792
rect 17368 6740 17374 6792
rect 17402 6740 17408 6792
rect 17460 6780 17466 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17460 6752 17601 6780
rect 17460 6740 17466 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 17736 6752 18153 6780
rect 17736 6740 17742 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 19242 6740 19248 6792
rect 19300 6740 19306 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 16684 6684 18552 6712
rect 17402 6644 17408 6656
rect 15712 6616 17408 6644
rect 15712 6604 15718 6616
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18524 6644 18552 6684
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 18693 6715 18751 6721
rect 18693 6712 18705 6715
rect 18656 6684 18705 6712
rect 18656 6672 18662 6684
rect 18693 6681 18705 6684
rect 18739 6681 18751 6715
rect 19444 6712 19472 6743
rect 20254 6740 20260 6792
rect 20312 6789 20318 6792
rect 20312 6783 20340 6789
rect 20328 6749 20340 6783
rect 20312 6743 20340 6749
rect 20312 6740 20318 6743
rect 20438 6740 20444 6792
rect 20496 6740 20502 6792
rect 21174 6740 21180 6792
rect 21232 6740 21238 6792
rect 23216 6789 23244 6820
rect 23566 6808 23572 6820
rect 23624 6848 23630 6860
rect 23860 6848 23888 6944
rect 24872 6848 24900 6956
rect 25038 6944 25044 6956
rect 25096 6944 25102 6996
rect 25314 6944 25320 6996
rect 25372 6984 25378 6996
rect 27246 6984 27252 6996
rect 25372 6956 27252 6984
rect 25372 6944 25378 6956
rect 27246 6944 27252 6956
rect 27304 6984 27310 6996
rect 27341 6987 27399 6993
rect 27341 6984 27353 6987
rect 27304 6956 27353 6984
rect 27304 6944 27310 6956
rect 27341 6953 27353 6956
rect 27387 6953 27399 6987
rect 27341 6947 27399 6953
rect 33594 6944 33600 6996
rect 33652 6984 33658 6996
rect 33793 6987 33851 6993
rect 33793 6984 33805 6987
rect 33652 6956 33805 6984
rect 33652 6944 33658 6956
rect 33793 6953 33805 6956
rect 33839 6953 33851 6987
rect 33793 6947 33851 6953
rect 35056 6987 35114 6993
rect 35056 6953 35068 6987
rect 35102 6984 35114 6987
rect 36814 6984 36820 6996
rect 35102 6956 36820 6984
rect 35102 6953 35114 6956
rect 35056 6947 35114 6953
rect 36814 6944 36820 6956
rect 36872 6944 36878 6996
rect 37277 6987 37335 6993
rect 37277 6953 37289 6987
rect 37323 6984 37335 6987
rect 37366 6984 37372 6996
rect 37323 6956 37372 6984
rect 37323 6953 37335 6956
rect 37277 6947 37335 6953
rect 37366 6944 37372 6956
rect 37424 6944 37430 6996
rect 39025 6987 39083 6993
rect 39025 6953 39037 6987
rect 39071 6984 39083 6987
rect 39298 6984 39304 6996
rect 39071 6956 39304 6984
rect 39071 6953 39083 6956
rect 39025 6947 39083 6953
rect 39298 6944 39304 6956
rect 39356 6944 39362 6996
rect 43530 6984 43536 6996
rect 43088 6956 43536 6984
rect 23624 6820 23888 6848
rect 24044 6820 24900 6848
rect 24964 6888 25912 6916
rect 23624 6808 23630 6820
rect 24044 6789 24072 6820
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 23201 6783 23259 6789
rect 23201 6749 23213 6783
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 23385 6783 23443 6789
rect 23385 6749 23397 6783
rect 23431 6780 23443 6783
rect 23477 6783 23535 6789
rect 23477 6780 23489 6783
rect 23431 6752 23489 6780
rect 23431 6749 23443 6752
rect 23385 6743 23443 6749
rect 23477 6749 23489 6752
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 18693 6675 18751 6681
rect 18800 6684 19472 6712
rect 18800 6644 18828 6684
rect 18524 6616 18828 6644
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 21376 6644 21404 6743
rect 23860 6712 23888 6743
rect 24302 6740 24308 6792
rect 24360 6740 24366 6792
rect 24394 6740 24400 6792
rect 24452 6780 24458 6792
rect 24964 6789 24992 6888
rect 25884 6860 25912 6888
rect 42794 6876 42800 6928
rect 42852 6876 42858 6928
rect 43088 6860 43116 6956
rect 43530 6944 43536 6956
rect 43588 6944 43594 6996
rect 25409 6851 25467 6857
rect 25409 6817 25421 6851
rect 25455 6848 25467 6851
rect 25774 6848 25780 6860
rect 25455 6820 25780 6848
rect 25455 6817 25467 6820
rect 25409 6811 25467 6817
rect 25774 6808 25780 6820
rect 25832 6808 25838 6860
rect 25866 6808 25872 6860
rect 25924 6848 25930 6860
rect 25924 6820 26924 6848
rect 25924 6808 25930 6820
rect 24949 6783 25007 6789
rect 24949 6780 24961 6783
rect 24452 6752 24961 6780
rect 24452 6740 24458 6752
rect 24949 6749 24961 6752
rect 24995 6749 25007 6783
rect 24949 6743 25007 6749
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 24320 6712 24348 6740
rect 24854 6712 24860 6724
rect 23860 6684 24860 6712
rect 24854 6672 24860 6684
rect 24912 6712 24918 6724
rect 25240 6712 25268 6743
rect 25958 6740 25964 6792
rect 26016 6780 26022 6792
rect 26896 6789 26924 6820
rect 31018 6808 31024 6860
rect 31076 6848 31082 6860
rect 31573 6851 31631 6857
rect 31573 6848 31585 6851
rect 31076 6820 31585 6848
rect 31076 6808 31082 6820
rect 31573 6817 31585 6820
rect 31619 6817 31631 6851
rect 31573 6811 31631 6817
rect 36541 6851 36599 6857
rect 36541 6817 36553 6851
rect 36587 6848 36599 6851
rect 36725 6851 36783 6857
rect 36725 6848 36737 6851
rect 36587 6820 36737 6848
rect 36587 6817 36599 6820
rect 36541 6811 36599 6817
rect 36725 6817 36737 6820
rect 36771 6848 36783 6851
rect 37458 6848 37464 6860
rect 36771 6820 37464 6848
rect 36771 6817 36783 6820
rect 36725 6811 36783 6817
rect 37458 6808 37464 6820
rect 37516 6808 37522 6860
rect 37550 6808 37556 6860
rect 37608 6808 37614 6860
rect 42429 6851 42487 6857
rect 42429 6817 42441 6851
rect 42475 6848 42487 6851
rect 42702 6848 42708 6860
rect 42475 6820 42708 6848
rect 42475 6817 42487 6820
rect 42429 6811 42487 6817
rect 42702 6808 42708 6820
rect 42760 6808 42766 6860
rect 42886 6808 42892 6860
rect 42944 6808 42950 6860
rect 43070 6808 43076 6860
rect 43128 6808 43134 6860
rect 43346 6808 43352 6860
rect 43404 6808 43410 6860
rect 26421 6783 26479 6789
rect 26421 6780 26433 6783
rect 26016 6752 26433 6780
rect 26016 6740 26022 6752
rect 26421 6749 26433 6752
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 26881 6783 26939 6789
rect 26881 6749 26893 6783
rect 26927 6780 26939 6783
rect 27062 6780 27068 6792
rect 26927 6752 27068 6780
rect 26927 6749 26939 6752
rect 26881 6743 26939 6749
rect 27062 6740 27068 6752
rect 27120 6740 27126 6792
rect 27249 6783 27307 6789
rect 27249 6749 27261 6783
rect 27295 6780 27307 6783
rect 27522 6780 27528 6792
rect 27295 6752 27528 6780
rect 27295 6749 27307 6752
rect 27249 6743 27307 6749
rect 24912 6684 25268 6712
rect 24912 6672 24918 6684
rect 19208 6616 21404 6644
rect 19208 6604 19214 6616
rect 23474 6604 23480 6656
rect 23532 6644 23538 6656
rect 23661 6647 23719 6653
rect 23661 6644 23673 6647
rect 23532 6616 23673 6644
rect 23532 6604 23538 6616
rect 23661 6613 23673 6616
rect 23707 6644 23719 6647
rect 24762 6644 24768 6656
rect 23707 6616 24768 6644
rect 23707 6613 23719 6616
rect 23661 6607 23719 6613
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 25038 6604 25044 6656
rect 25096 6644 25102 6656
rect 25976 6644 26004 6740
rect 26789 6715 26847 6721
rect 26789 6681 26801 6715
rect 26835 6712 26847 6715
rect 27264 6712 27292 6743
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 30929 6783 30987 6789
rect 30929 6780 30941 6783
rect 30208 6752 30941 6780
rect 26835 6684 27292 6712
rect 26835 6681 26847 6684
rect 26789 6675 26847 6681
rect 30208 6656 30236 6752
rect 30929 6749 30941 6752
rect 30975 6780 30987 6783
rect 31389 6783 31447 6789
rect 31389 6780 31401 6783
rect 30975 6752 31401 6780
rect 30975 6749 30987 6752
rect 30929 6743 30987 6749
rect 31389 6749 31401 6752
rect 31435 6749 31447 6783
rect 31389 6743 31447 6749
rect 34057 6783 34115 6789
rect 34057 6749 34069 6783
rect 34103 6780 34115 6783
rect 34514 6780 34520 6792
rect 34103 6752 34520 6780
rect 34103 6749 34115 6752
rect 34057 6743 34115 6749
rect 34514 6740 34520 6752
rect 34572 6780 34578 6792
rect 34793 6783 34851 6789
rect 34793 6780 34805 6783
rect 34572 6752 34805 6780
rect 34572 6740 34578 6752
rect 34793 6749 34805 6752
rect 34839 6749 34851 6783
rect 34793 6743 34851 6749
rect 37918 6740 37924 6792
rect 37976 6780 37982 6792
rect 38841 6783 38899 6789
rect 38841 6780 38853 6783
rect 37976 6752 38853 6780
rect 37976 6740 37982 6752
rect 38841 6749 38853 6752
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 39114 6740 39120 6792
rect 39172 6780 39178 6792
rect 39209 6783 39267 6789
rect 39209 6780 39221 6783
rect 39172 6752 39221 6780
rect 39172 6740 39178 6752
rect 39209 6749 39221 6752
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 39393 6783 39451 6789
rect 39393 6749 39405 6783
rect 39439 6780 39451 6783
rect 39666 6780 39672 6792
rect 39439 6752 39672 6780
rect 39439 6749 39451 6752
rect 39393 6743 39451 6749
rect 39666 6740 39672 6752
rect 39724 6740 39730 6792
rect 31202 6672 31208 6724
rect 31260 6672 31266 6724
rect 36354 6712 36360 6724
rect 32232 6684 32614 6712
rect 36294 6684 36360 6712
rect 32232 6656 32260 6684
rect 36354 6672 36360 6684
rect 36412 6712 36418 6724
rect 36722 6712 36728 6724
rect 36412 6684 36728 6712
rect 36412 6672 36418 6684
rect 36722 6672 36728 6684
rect 36780 6712 36786 6724
rect 36998 6712 37004 6724
rect 36780 6684 37004 6712
rect 36780 6672 36786 6684
rect 36998 6672 37004 6684
rect 37056 6672 37062 6724
rect 39574 6672 39580 6724
rect 39632 6672 39638 6724
rect 43438 6672 43444 6724
rect 43496 6712 43502 6724
rect 43496 6684 43838 6712
rect 43496 6672 43502 6684
rect 25096 6616 26004 6644
rect 25096 6604 25102 6616
rect 30190 6604 30196 6656
rect 30248 6604 30254 6656
rect 31018 6604 31024 6656
rect 31076 6604 31082 6656
rect 32214 6604 32220 6656
rect 32272 6604 32278 6656
rect 32309 6647 32367 6653
rect 32309 6613 32321 6647
rect 32355 6644 32367 6647
rect 33042 6644 33048 6656
rect 32355 6616 33048 6644
rect 32355 6613 32367 6616
rect 32309 6607 32367 6613
rect 33042 6604 33048 6616
rect 33100 6604 33106 6656
rect 38194 6604 38200 6656
rect 38252 6604 38258 6656
rect 38286 6604 38292 6656
rect 38344 6604 38350 6656
rect 39206 6604 39212 6656
rect 39264 6644 39270 6656
rect 39301 6647 39359 6653
rect 39301 6644 39313 6647
rect 39264 6616 39313 6644
rect 39264 6604 39270 6616
rect 39301 6613 39313 6616
rect 39347 6613 39359 6647
rect 39301 6607 39359 6613
rect 44821 6647 44879 6653
rect 44821 6613 44833 6647
rect 44867 6644 44879 6647
rect 44867 6616 45232 6644
rect 44867 6613 44879 6616
rect 44821 6607 44879 6613
rect 1104 6554 45172 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 45172 6554
rect 1104 6480 45172 6502
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 5718 6440 5724 6452
rect 4479 6412 5724 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6362 6400 6368 6452
rect 6420 6400 6426 6452
rect 8159 6443 8217 6449
rect 8159 6409 8171 6443
rect 8205 6440 8217 6443
rect 9490 6440 9496 6452
rect 8205 6412 9496 6440
rect 8205 6409 8217 6412
rect 8159 6403 8217 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 13412 6412 14933 6440
rect 13412 6400 13418 6412
rect 14921 6409 14933 6412
rect 14967 6440 14979 6443
rect 15286 6440 15292 6452
rect 14967 6412 15292 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 17313 6443 17371 6449
rect 15427 6412 17080 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 5442 6332 5448 6384
rect 5500 6332 5506 6384
rect 6380 6304 6408 6400
rect 7282 6332 7288 6384
rect 7340 6332 7346 6384
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 14277 6375 14335 6381
rect 14277 6372 14289 6375
rect 13320 6344 14289 6372
rect 13320 6332 13326 6344
rect 14277 6341 14289 6344
rect 14323 6341 14335 6375
rect 14277 6335 14335 6341
rect 14476 6344 14780 6372
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6380 6276 6745 6304
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 9640 6276 9706 6304
rect 9640 6264 9646 6276
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14476 6313 14504 6344
rect 14752 6316 14780 6344
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 15252 6344 16344 6372
rect 15252 6332 15258 6344
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 13872 6276 14473 6304
rect 13872 6264 13878 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 5902 6196 5908 6248
rect 5960 6196 5966 6248
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 6227 6208 6377 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6365 6205 6377 6208
rect 6411 6236 6423 6239
rect 6914 6236 6920 6248
rect 6411 6208 6920 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 6196 6100 6224 6199
rect 6914 6196 6920 6208
rect 6972 6236 6978 6248
rect 8202 6236 8208 6248
rect 6972 6208 8208 6236
rect 6972 6196 6978 6208
rect 8202 6196 8208 6208
rect 8260 6236 8266 6248
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8260 6208 8309 6236
rect 8260 6196 8266 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8570 6196 8576 6248
rect 8628 6196 8634 6248
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6236 10103 6239
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10091 6208 10241 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 12158 6196 12164 6248
rect 12216 6236 12222 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12216 6208 13001 6236
rect 12216 6196 12222 6208
rect 12989 6205 13001 6208
rect 13035 6205 13047 6239
rect 13648 6236 13676 6264
rect 14090 6236 14096 6248
rect 13648 6208 14096 6236
rect 12989 6199 13047 6205
rect 3844 6072 6224 6100
rect 3844 6060 3850 6072
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10376 6072 10885 6100
rect 10376 6060 10382 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 13004 6100 13032 6199
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14568 6236 14596 6267
rect 14734 6264 14740 6316
rect 14792 6264 14798 6316
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14884 6276 15025 6304
rect 14884 6264 14890 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 14424 6208 14596 6236
rect 15028 6236 15056 6267
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 15930 6304 15936 6316
rect 15764 6276 15936 6304
rect 15488 6236 15516 6264
rect 15764 6245 15792 6276
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16316 6313 16344 6344
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16482 6304 16488 6316
rect 16347 6276 16488 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 15028 6208 15516 6236
rect 15565 6239 15623 6245
rect 14424 6196 14430 6208
rect 15565 6205 15577 6239
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16040 6236 16068 6264
rect 15887 6208 16068 6236
rect 16117 6239 16175 6245
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16117 6205 16129 6239
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 13354 6128 13360 6180
rect 13412 6128 13418 6180
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 15580 6168 15608 6199
rect 13504 6140 15608 6168
rect 15672 6168 15700 6199
rect 16132 6168 16160 6199
rect 16942 6196 16948 6248
rect 17000 6196 17006 6248
rect 17052 6236 17080 6412
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 17678 6440 17684 6452
rect 17359 6412 17684 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 19061 6443 19119 6449
rect 19061 6409 19073 6443
rect 19107 6440 19119 6443
rect 20254 6440 20260 6452
rect 19107 6412 20260 6440
rect 19107 6409 19119 6412
rect 19061 6403 19119 6409
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6440 23903 6443
rect 33870 6440 33876 6452
rect 23891 6412 24900 6440
rect 23891 6409 23903 6412
rect 23845 6403 23903 6409
rect 17494 6332 17500 6384
rect 17552 6332 17558 6384
rect 17126 6264 17132 6316
rect 17184 6264 17190 6316
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 17696 6304 17724 6400
rect 18506 6332 18512 6384
rect 18564 6372 18570 6384
rect 19245 6375 19303 6381
rect 19245 6372 19257 6375
rect 18564 6344 19257 6372
rect 18564 6332 18570 6344
rect 19245 6341 19257 6344
rect 19291 6341 19303 6375
rect 19245 6335 19303 6341
rect 19426 6332 19432 6384
rect 19484 6372 19490 6384
rect 19889 6375 19947 6381
rect 19889 6372 19901 6375
rect 19484 6344 19901 6372
rect 19484 6332 19490 6344
rect 19889 6341 19901 6344
rect 19935 6372 19947 6375
rect 20438 6372 20444 6384
rect 19935 6344 20444 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 17635 6276 17724 6304
rect 18708 6276 19073 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 18414 6236 18420 6248
rect 17052 6208 18420 6236
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 15672 6140 16160 6168
rect 16485 6171 16543 6177
rect 13504 6128 13510 6140
rect 13909 6103 13967 6109
rect 13909 6100 13921 6103
rect 13004 6072 13921 6100
rect 10873 6063 10931 6069
rect 13909 6069 13921 6072
rect 13955 6100 13967 6103
rect 14090 6100 14096 6112
rect 13955 6072 14096 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 15378 6100 15384 6112
rect 14792 6072 15384 6100
rect 14792 6060 14798 6072
rect 15378 6060 15384 6072
rect 15436 6100 15442 6112
rect 15672 6100 15700 6140
rect 16485 6137 16497 6171
rect 16531 6168 16543 6171
rect 18708 6168 18736 6276
rect 19061 6273 19073 6276
rect 19107 6304 19119 6307
rect 19150 6304 19156 6316
rect 19107 6276 19156 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 19392 6276 19472 6304
rect 19392 6264 19398 6276
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6236 18843 6239
rect 18874 6236 18880 6248
rect 18831 6208 18880 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 16531 6140 18736 6168
rect 18969 6171 19027 6177
rect 16531 6137 16543 6140
rect 16485 6131 16543 6137
rect 18969 6137 18981 6171
rect 19015 6168 19027 6171
rect 19058 6168 19064 6180
rect 19015 6140 19064 6168
rect 19015 6137 19027 6140
rect 18969 6131 19027 6137
rect 19058 6128 19064 6140
rect 19116 6128 19122 6180
rect 19444 6112 19472 6276
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 23566 6264 23572 6316
rect 23624 6264 23630 6316
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6304 23811 6307
rect 23860 6304 23888 6403
rect 24029 6375 24087 6381
rect 24029 6341 24041 6375
rect 24075 6372 24087 6375
rect 24302 6372 24308 6384
rect 24075 6344 24308 6372
rect 24075 6341 24087 6344
rect 24029 6335 24087 6341
rect 24302 6332 24308 6344
rect 24360 6332 24366 6384
rect 24872 6381 24900 6412
rect 25792 6412 33876 6440
rect 24857 6375 24915 6381
rect 24857 6341 24869 6375
rect 24903 6341 24915 6375
rect 24857 6335 24915 6341
rect 24949 6375 25007 6381
rect 24949 6341 24961 6375
rect 24995 6372 25007 6375
rect 25792 6372 25820 6412
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 33962 6400 33968 6452
rect 34020 6400 34026 6452
rect 36906 6400 36912 6452
rect 36964 6440 36970 6452
rect 37918 6449 37924 6452
rect 37277 6443 37335 6449
rect 37277 6440 37289 6443
rect 36964 6412 37289 6440
rect 36964 6400 36970 6412
rect 37277 6409 37289 6412
rect 37323 6440 37335 6443
rect 37914 6440 37924 6449
rect 37323 6412 37780 6440
rect 37879 6412 37924 6440
rect 37323 6409 37335 6412
rect 37277 6403 37335 6409
rect 24995 6344 25820 6372
rect 24995 6341 25007 6344
rect 24949 6335 25007 6341
rect 23799 6276 23888 6304
rect 23799 6273 23811 6276
rect 23753 6267 23811 6273
rect 24394 6264 24400 6316
rect 24452 6264 24458 6316
rect 24673 6307 24731 6313
rect 24673 6273 24685 6307
rect 24719 6273 24731 6307
rect 24673 6267 24731 6273
rect 24688 6236 24716 6267
rect 24762 6264 24768 6316
rect 24820 6304 24826 6316
rect 25792 6313 25820 6344
rect 33781 6375 33839 6381
rect 33781 6341 33793 6375
rect 33827 6372 33839 6375
rect 33980 6372 34008 6400
rect 33827 6344 34008 6372
rect 33827 6341 33839 6344
rect 33781 6335 33839 6341
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24820 6276 25053 6304
rect 24820 6264 24826 6276
rect 25041 6273 25053 6276
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 25777 6307 25835 6313
rect 25777 6273 25789 6307
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 30374 6264 30380 6316
rect 30432 6304 30438 6316
rect 34057 6307 34115 6313
rect 30432 6276 30590 6304
rect 32232 6276 32706 6304
rect 30432 6264 30438 6276
rect 24688 6208 25728 6236
rect 24854 6128 24860 6180
rect 24912 6168 24918 6180
rect 25317 6171 25375 6177
rect 25317 6168 25329 6171
rect 24912 6140 25329 6168
rect 24912 6128 24918 6140
rect 25317 6137 25329 6140
rect 25363 6137 25375 6171
rect 25317 6131 25375 6137
rect 15436 6072 15700 6100
rect 15436 6060 15442 6072
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 18598 6100 18604 6112
rect 15988 6072 18604 6100
rect 15988 6060 15994 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 19426 6060 19432 6112
rect 19484 6060 19490 6112
rect 23750 6060 23756 6112
rect 23808 6060 23814 6112
rect 23934 6060 23940 6112
rect 23992 6100 23998 6112
rect 24029 6103 24087 6109
rect 24029 6100 24041 6103
rect 23992 6072 24041 6100
rect 23992 6060 23998 6072
rect 24029 6069 24041 6072
rect 24075 6100 24087 6103
rect 25038 6100 25044 6112
rect 24075 6072 25044 6100
rect 24075 6069 24087 6072
rect 24029 6063 24087 6069
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 25222 6060 25228 6112
rect 25280 6060 25286 6112
rect 25700 6109 25728 6208
rect 29454 6196 29460 6248
rect 29512 6196 29518 6248
rect 30190 6196 30196 6248
rect 30248 6196 30254 6248
rect 31662 6196 31668 6248
rect 31720 6196 31726 6248
rect 31941 6239 31999 6245
rect 31941 6205 31953 6239
rect 31987 6205 31999 6239
rect 31941 6199 31999 6205
rect 29564 6140 30236 6168
rect 29564 6112 29592 6140
rect 25685 6103 25743 6109
rect 25685 6069 25697 6103
rect 25731 6100 25743 6103
rect 26142 6100 26148 6112
rect 25731 6072 26148 6100
rect 25731 6069 25743 6072
rect 25685 6063 25743 6069
rect 26142 6060 26148 6072
rect 26200 6060 26206 6112
rect 29546 6060 29552 6112
rect 29604 6060 29610 6112
rect 29914 6060 29920 6112
rect 29972 6100 29978 6112
rect 30101 6103 30159 6109
rect 30101 6100 30113 6103
rect 29972 6072 30113 6100
rect 29972 6060 29978 6072
rect 30101 6069 30113 6072
rect 30147 6069 30159 6103
rect 30208 6100 30236 6140
rect 31956 6100 31984 6199
rect 32232 6112 32260 6276
rect 34057 6273 34069 6307
rect 34103 6304 34115 6307
rect 34514 6304 34520 6316
rect 34103 6276 34520 6304
rect 34103 6273 34115 6276
rect 34057 6267 34115 6273
rect 34514 6264 34520 6276
rect 34572 6264 34578 6316
rect 36924 6313 36952 6400
rect 37090 6332 37096 6384
rect 37148 6332 37154 6384
rect 37445 6375 37503 6381
rect 37445 6341 37457 6375
rect 37491 6372 37503 6375
rect 37491 6344 37596 6372
rect 37491 6341 37503 6344
rect 37445 6335 37503 6341
rect 36909 6307 36967 6313
rect 36909 6273 36921 6307
rect 36955 6273 36967 6307
rect 37568 6304 37596 6344
rect 37642 6332 37648 6384
rect 37700 6332 37706 6384
rect 37752 6372 37780 6412
rect 37914 6403 37924 6412
rect 37918 6400 37924 6403
rect 37976 6400 37982 6452
rect 38194 6440 38200 6452
rect 38028 6412 38200 6440
rect 38028 6381 38056 6412
rect 38194 6400 38200 6412
rect 38252 6400 38258 6452
rect 38286 6400 38292 6452
rect 38344 6400 38350 6452
rect 41782 6400 41788 6452
rect 41840 6400 41846 6452
rect 42429 6443 42487 6449
rect 42429 6409 42441 6443
rect 42475 6440 42487 6443
rect 42702 6440 42708 6452
rect 42475 6412 42708 6440
rect 42475 6409 42487 6412
rect 42429 6403 42487 6409
rect 42702 6400 42708 6412
rect 42760 6400 42766 6452
rect 42794 6400 42800 6452
rect 42852 6440 42858 6452
rect 43073 6443 43131 6449
rect 43073 6440 43085 6443
rect 42852 6412 43085 6440
rect 42852 6400 42858 6412
rect 43073 6409 43085 6412
rect 43119 6409 43131 6443
rect 43073 6403 43131 6409
rect 44634 6400 44640 6452
rect 44692 6400 44698 6452
rect 45204 6440 45232 6616
rect 44744 6412 45232 6440
rect 38013 6375 38071 6381
rect 37752 6344 37964 6372
rect 37734 6304 37740 6316
rect 37568 6276 37740 6304
rect 36909 6267 36967 6273
rect 37734 6264 37740 6276
rect 37792 6264 37798 6316
rect 37829 6307 37887 6313
rect 37829 6273 37841 6307
rect 37875 6273 37887 6307
rect 37936 6304 37964 6344
rect 38013 6341 38025 6375
rect 38059 6341 38071 6375
rect 38013 6335 38071 6341
rect 38105 6307 38163 6313
rect 38105 6304 38117 6307
rect 37936 6276 38117 6304
rect 37829 6267 37887 6273
rect 38105 6273 38117 6276
rect 38151 6273 38163 6307
rect 38105 6267 38163 6273
rect 38197 6307 38255 6313
rect 38197 6273 38209 6307
rect 38243 6304 38255 6307
rect 38304 6304 38332 6400
rect 41800 6372 41828 6400
rect 44744 6372 44772 6412
rect 45278 6372 45284 6384
rect 41800 6344 44772 6372
rect 44836 6344 45284 6372
rect 38243 6276 38332 6304
rect 38243 6273 38255 6276
rect 38197 6267 38255 6273
rect 36725 6239 36783 6245
rect 36725 6205 36737 6239
rect 36771 6236 36783 6239
rect 37458 6236 37464 6248
rect 36771 6208 37464 6236
rect 36771 6205 36783 6208
rect 36725 6199 36783 6205
rect 37458 6196 37464 6208
rect 37516 6196 37522 6248
rect 37642 6196 37648 6248
rect 37700 6236 37706 6248
rect 37844 6236 37872 6267
rect 42242 6264 42248 6316
rect 42300 6304 42306 6316
rect 42720 6313 42748 6344
rect 42613 6307 42671 6313
rect 42613 6304 42625 6307
rect 42300 6276 42625 6304
rect 42300 6264 42306 6276
rect 42613 6273 42625 6276
rect 42659 6273 42671 6307
rect 42613 6267 42671 6273
rect 42705 6307 42763 6313
rect 42705 6273 42717 6307
rect 42751 6273 42763 6307
rect 42705 6267 42763 6273
rect 42797 6307 42855 6313
rect 42797 6273 42809 6307
rect 42843 6304 42855 6307
rect 42886 6304 42892 6316
rect 42843 6276 42892 6304
rect 42843 6273 42855 6276
rect 42797 6267 42855 6273
rect 38381 6239 38439 6245
rect 38381 6236 38393 6239
rect 37700 6208 37872 6236
rect 37936 6208 38393 6236
rect 37700 6196 37706 6208
rect 37936 6168 37964 6208
rect 38381 6205 38393 6208
rect 38427 6236 38439 6239
rect 38654 6236 38660 6248
rect 38427 6208 38660 6236
rect 38427 6205 38439 6208
rect 38381 6199 38439 6205
rect 38654 6196 38660 6208
rect 38712 6196 38718 6248
rect 38746 6196 38752 6248
rect 38804 6196 38810 6248
rect 42628 6236 42656 6267
rect 42886 6264 42892 6276
rect 42944 6304 42950 6316
rect 43548 6313 43576 6344
rect 44836 6313 44864 6344
rect 45278 6332 45284 6344
rect 45336 6332 45342 6384
rect 43349 6307 43407 6313
rect 43349 6304 43361 6307
rect 42944 6276 43361 6304
rect 42944 6264 42950 6276
rect 43349 6273 43361 6276
rect 43395 6273 43407 6307
rect 43349 6267 43407 6273
rect 43533 6307 43591 6313
rect 43533 6273 43545 6307
rect 43579 6273 43591 6307
rect 43533 6267 43591 6273
rect 44821 6307 44879 6313
rect 44821 6273 44833 6307
rect 44867 6273 44879 6307
rect 44821 6267 44879 6273
rect 43257 6239 43315 6245
rect 43257 6236 43269 6239
rect 42628 6208 43269 6236
rect 43257 6205 43269 6208
rect 43303 6205 43315 6239
rect 43257 6199 43315 6205
rect 43441 6239 43499 6245
rect 43441 6205 43453 6239
rect 43487 6205 43499 6239
rect 43441 6199 43499 6205
rect 37384 6140 37964 6168
rect 38105 6171 38163 6177
rect 30208 6072 31984 6100
rect 30101 6063 30159 6069
rect 32214 6060 32220 6112
rect 32272 6060 32278 6112
rect 32309 6103 32367 6109
rect 32309 6069 32321 6103
rect 32355 6100 32367 6103
rect 33134 6100 33140 6112
rect 32355 6072 33140 6100
rect 32355 6069 32367 6072
rect 32309 6063 32367 6069
rect 33134 6060 33140 6072
rect 33192 6060 33198 6112
rect 36538 6060 36544 6112
rect 36596 6100 36602 6112
rect 37384 6100 37412 6140
rect 38105 6137 38117 6171
rect 38151 6168 38163 6171
rect 38764 6168 38792 6196
rect 38151 6140 38792 6168
rect 38151 6137 38163 6140
rect 38105 6131 38163 6137
rect 42978 6128 42984 6180
rect 43036 6168 43042 6180
rect 43456 6168 43484 6199
rect 43036 6140 43484 6168
rect 43036 6128 43042 6140
rect 36596 6072 37412 6100
rect 37461 6103 37519 6109
rect 36596 6060 36602 6072
rect 37461 6069 37473 6103
rect 37507 6100 37519 6103
rect 37550 6100 37556 6112
rect 37507 6072 37556 6100
rect 37507 6069 37519 6072
rect 37461 6063 37519 6069
rect 37550 6060 37556 6072
rect 37608 6060 37614 6112
rect 1104 6010 45172 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 45172 6010
rect 1104 5936 45172 5958
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 5960 5868 6377 5896
rect 5960 5856 5966 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7282 5896 7288 5908
rect 6779 5868 7288 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 3786 5692 3792 5704
rect 3292 5664 3792 5692
rect 3292 5652 3298 5664
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 5583 5695 5641 5701
rect 5583 5661 5595 5695
rect 5629 5692 5641 5695
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5629 5664 5733 5692
rect 5629 5661 5641 5664
rect 5583 5655 5641 5661
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5442 5624 5448 5636
rect 5198 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5624 5506 5636
rect 6748 5624 6776 5859
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8628 5868 8953 5896
rect 8628 5856 8634 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 12032 5868 13553 5896
rect 12032 5856 12038 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14424 5868 14657 5896
rect 14424 5856 14430 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 15378 5856 15384 5908
rect 15436 5856 15442 5908
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5865 15991 5899
rect 15933 5859 15991 5865
rect 9582 5828 9588 5840
rect 8404 5800 9588 5828
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6972 5732 7021 5760
rect 6972 5720 6978 5732
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 8404 5678 8432 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 11839 5831 11897 5837
rect 11839 5797 11851 5831
rect 11885 5828 11897 5831
rect 12250 5828 12256 5840
rect 11885 5800 12256 5828
rect 11885 5797 11897 5800
rect 11839 5791 11897 5797
rect 12250 5788 12256 5800
rect 12308 5828 12314 5840
rect 13998 5828 14004 5840
rect 12308 5800 14004 5828
rect 12308 5788 12314 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 15948 5828 15976 5859
rect 16942 5856 16948 5908
rect 17000 5856 17006 5908
rect 17957 5899 18015 5905
rect 17957 5865 17969 5899
rect 18003 5896 18015 5899
rect 18230 5896 18236 5908
rect 18003 5868 18236 5896
rect 18003 5865 18015 5868
rect 17957 5859 18015 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 19242 5856 19248 5908
rect 19300 5856 19306 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20864 5868 21005 5896
rect 20864 5856 20870 5868
rect 20993 5865 21005 5868
rect 21039 5865 21051 5899
rect 20993 5859 21051 5865
rect 23750 5856 23756 5908
rect 23808 5856 23814 5908
rect 23842 5856 23848 5908
rect 23900 5896 23906 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23900 5868 24409 5896
rect 23900 5856 23906 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 24397 5859 24455 5865
rect 25222 5856 25228 5908
rect 25280 5896 25286 5908
rect 25758 5899 25816 5905
rect 25758 5896 25770 5899
rect 25280 5868 25770 5896
rect 25280 5856 25286 5868
rect 25758 5865 25770 5868
rect 25804 5865 25816 5899
rect 25758 5859 25816 5865
rect 26142 5856 26148 5908
rect 26200 5896 26206 5908
rect 29365 5899 29423 5905
rect 26200 5868 29224 5896
rect 26200 5856 26206 5868
rect 14148 5800 15976 5828
rect 14148 5788 14154 5800
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5729 8815 5763
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 8757 5723 8815 5729
rect 9692 5732 10057 5760
rect 8772 5692 8800 5723
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 8772 5664 9505 5692
rect 9493 5661 9505 5664
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9692 5636 9720 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 14642 5760 14648 5772
rect 13412 5732 14648 5760
rect 13412 5720 13418 5732
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5760 15071 5763
rect 15286 5760 15292 5772
rect 15059 5732 15292 5760
rect 15059 5729 15071 5732
rect 15013 5723 15071 5729
rect 15286 5720 15292 5732
rect 15344 5760 15350 5772
rect 16117 5763 16175 5769
rect 15344 5732 15792 5760
rect 15344 5720 15350 5732
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 13630 5692 13636 5704
rect 13096 5664 13636 5692
rect 13096 5636 13124 5664
rect 13630 5652 13636 5664
rect 13688 5692 13694 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13688 5664 13737 5692
rect 13688 5652 13694 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 5500 5596 6776 5624
rect 6825 5627 6883 5633
rect 5500 5584 5506 5596
rect 6825 5593 6837 5627
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 7285 5627 7343 5633
rect 7285 5593 7297 5627
rect 7331 5624 7343 5627
rect 7558 5624 7564 5636
rect 7331 5596 7564 5624
rect 7331 5593 7343 5596
rect 7285 5587 7343 5593
rect 6840 5556 6868 5587
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 9674 5584 9680 5636
rect 9732 5584 9738 5636
rect 10962 5584 10968 5636
rect 11020 5584 11026 5636
rect 13078 5584 13084 5636
rect 13136 5584 13142 5636
rect 13740 5624 13768 5655
rect 13906 5652 13912 5704
rect 13964 5652 13970 5704
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14274 5692 14280 5704
rect 14056 5664 14280 5692
rect 14056 5652 14062 5664
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14660 5692 14688 5720
rect 15194 5692 15200 5704
rect 14660 5664 15200 5692
rect 14553 5655 14611 5661
rect 14568 5624 14596 5655
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 15657 5695 15715 5701
rect 15519 5664 15608 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 15580 5636 15608 5664
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15764 5692 15792 5732
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16163 5732 16405 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16393 5729 16405 5732
rect 16439 5760 16451 5763
rect 16960 5760 16988 5856
rect 16439 5732 16988 5760
rect 16439 5729 16451 5732
rect 16393 5723 16451 5729
rect 17586 5720 17592 5772
rect 17644 5720 17650 5772
rect 16206 5692 16212 5704
rect 15764 5664 16212 5692
rect 15657 5655 15715 5661
rect 13740 5596 14596 5624
rect 15562 5584 15568 5636
rect 15620 5584 15626 5636
rect 9766 5556 9772 5568
rect 6840 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 14185 5559 14243 5565
rect 14185 5525 14197 5559
rect 14231 5556 14243 5559
rect 15102 5556 15108 5568
rect 14231 5528 15108 5556
rect 14231 5525 14243 5528
rect 14185 5519 14243 5525
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15672 5556 15700 5655
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 16540 5664 16589 5692
rect 16540 5652 16546 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 17604 5692 17632 5720
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 16577 5655 16635 5661
rect 17420 5664 17785 5692
rect 17420 5636 17448 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 16022 5584 16028 5636
rect 16080 5624 16086 5636
rect 16301 5627 16359 5633
rect 16301 5624 16313 5627
rect 16080 5596 16313 5624
rect 16080 5584 16086 5596
rect 16301 5593 16313 5596
rect 16347 5593 16359 5627
rect 16301 5587 16359 5593
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 17586 5584 17592 5636
rect 17644 5584 17650 5636
rect 15252 5528 15700 5556
rect 16485 5559 16543 5565
rect 15252 5516 15258 5528
rect 16485 5525 16497 5559
rect 16531 5556 16543 5559
rect 19260 5556 19288 5856
rect 23768 5760 23796 5856
rect 24302 5788 24308 5840
rect 24360 5828 24366 5840
rect 24360 5800 25268 5828
rect 24360 5788 24366 5800
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 23768 5732 24869 5760
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5729 25099 5763
rect 25041 5723 25099 5729
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5692 20959 5695
rect 21174 5692 21180 5704
rect 20947 5664 21180 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 23753 5695 23811 5701
rect 23753 5661 23765 5695
rect 23799 5692 23811 5695
rect 23934 5692 23940 5704
rect 23799 5664 23940 5692
rect 23799 5661 23811 5664
rect 23753 5655 23811 5661
rect 23934 5652 23940 5664
rect 23992 5652 23998 5704
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 24118 5692 24124 5704
rect 24075 5664 24124 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 24118 5652 24124 5664
rect 24176 5692 24182 5704
rect 24394 5692 24400 5704
rect 24176 5664 24400 5692
rect 24176 5652 24182 5664
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 24213 5627 24271 5633
rect 24213 5593 24225 5627
rect 24259 5624 24271 5627
rect 25056 5624 25084 5723
rect 25240 5701 25268 5800
rect 27617 5763 27675 5769
rect 27617 5760 27629 5763
rect 25516 5732 27629 5760
rect 25516 5704 25544 5732
rect 27617 5729 27629 5732
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 25225 5695 25283 5701
rect 25225 5661 25237 5695
rect 25271 5661 25283 5695
rect 25225 5655 25283 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 25424 5624 25452 5655
rect 25498 5652 25504 5704
rect 25556 5652 25562 5704
rect 27062 5652 27068 5704
rect 27120 5692 27126 5704
rect 27525 5695 27583 5701
rect 27525 5692 27537 5695
rect 27120 5664 27537 5692
rect 27120 5652 27126 5664
rect 27525 5661 27537 5664
rect 27571 5661 27583 5695
rect 27525 5655 27583 5661
rect 28994 5652 29000 5704
rect 29052 5652 29058 5704
rect 27338 5624 27344 5636
rect 24259 5596 24808 5624
rect 25056 5596 26188 5624
rect 27002 5596 27344 5624
rect 24259 5593 24271 5596
rect 24213 5587 24271 5593
rect 16531 5528 19288 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 23845 5559 23903 5565
rect 23845 5556 23857 5559
rect 23624 5528 23857 5556
rect 23624 5516 23630 5528
rect 23845 5525 23857 5528
rect 23891 5556 23903 5559
rect 24302 5556 24308 5568
rect 23891 5528 24308 5556
rect 23891 5525 23903 5528
rect 23845 5519 23903 5525
rect 24302 5516 24308 5528
rect 24360 5516 24366 5568
rect 24780 5565 24808 5596
rect 26160 5568 26188 5596
rect 27338 5584 27344 5596
rect 27396 5584 27402 5636
rect 27893 5627 27951 5633
rect 27893 5593 27905 5627
rect 27939 5593 27951 5627
rect 27893 5587 27951 5593
rect 24765 5559 24823 5565
rect 24765 5525 24777 5559
rect 24811 5525 24823 5559
rect 24765 5519 24823 5525
rect 25317 5559 25375 5565
rect 25317 5525 25329 5559
rect 25363 5556 25375 5559
rect 25498 5556 25504 5568
rect 25363 5528 25504 5556
rect 25363 5525 25375 5528
rect 25317 5519 25375 5525
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 26142 5516 26148 5568
rect 26200 5516 26206 5568
rect 27154 5516 27160 5568
rect 27212 5556 27218 5568
rect 27908 5556 27936 5587
rect 27212 5528 27936 5556
rect 29196 5556 29224 5868
rect 29365 5865 29377 5899
rect 29411 5896 29423 5899
rect 29454 5896 29460 5908
rect 29411 5868 29460 5896
rect 29411 5865 29423 5868
rect 29365 5859 29423 5865
rect 29454 5856 29460 5868
rect 29512 5856 29518 5908
rect 31018 5856 31024 5908
rect 31076 5856 31082 5908
rect 31202 5856 31208 5908
rect 31260 5896 31266 5908
rect 31297 5899 31355 5905
rect 31297 5896 31309 5899
rect 31260 5868 31309 5896
rect 31260 5856 31266 5868
rect 31297 5865 31309 5868
rect 31343 5865 31355 5899
rect 31297 5859 31355 5865
rect 31662 5856 31668 5908
rect 31720 5896 31726 5908
rect 32217 5899 32275 5905
rect 32217 5896 32229 5899
rect 31720 5868 32229 5896
rect 31720 5856 31726 5868
rect 32217 5865 32229 5868
rect 32263 5865 32275 5899
rect 32217 5859 32275 5865
rect 32306 5856 32312 5908
rect 32364 5856 32370 5908
rect 33042 5856 33048 5908
rect 33100 5856 33106 5908
rect 33134 5856 33140 5908
rect 33192 5896 33198 5908
rect 33689 5899 33747 5905
rect 33689 5896 33701 5899
rect 33192 5868 33701 5896
rect 33192 5856 33198 5868
rect 29825 5763 29883 5769
rect 29825 5729 29837 5763
rect 29871 5760 29883 5763
rect 29914 5760 29920 5772
rect 29871 5732 29920 5760
rect 29871 5729 29883 5732
rect 29825 5723 29883 5729
rect 29914 5720 29920 5732
rect 29972 5720 29978 5772
rect 31036 5760 31064 5856
rect 32140 5800 32628 5828
rect 32140 5760 32168 5800
rect 31036 5732 32168 5760
rect 29546 5652 29552 5704
rect 29604 5652 29610 5704
rect 31202 5652 31208 5704
rect 31260 5652 31266 5704
rect 31570 5652 31576 5704
rect 31628 5652 31634 5704
rect 31662 5652 31668 5704
rect 31720 5692 31726 5704
rect 32600 5701 32628 5800
rect 33060 5760 33088 5856
rect 33244 5837 33272 5868
rect 33689 5865 33701 5868
rect 33735 5865 33747 5899
rect 33689 5859 33747 5865
rect 33870 5856 33876 5908
rect 33928 5896 33934 5908
rect 34057 5899 34115 5905
rect 34057 5896 34069 5899
rect 33928 5868 34069 5896
rect 33928 5856 33934 5868
rect 34057 5865 34069 5868
rect 34103 5865 34115 5899
rect 34057 5859 34115 5865
rect 37829 5899 37887 5905
rect 37829 5865 37841 5899
rect 37875 5896 37887 5899
rect 39574 5896 39580 5908
rect 37875 5868 39580 5896
rect 37875 5865 37887 5868
rect 37829 5859 37887 5865
rect 39574 5856 39580 5868
rect 39632 5856 39638 5908
rect 33229 5831 33287 5837
rect 33229 5797 33241 5831
rect 33275 5797 33287 5831
rect 33229 5791 33287 5797
rect 33505 5763 33563 5769
rect 33505 5760 33517 5763
rect 33060 5732 33517 5760
rect 33505 5729 33517 5732
rect 33551 5760 33563 5763
rect 33551 5732 33640 5760
rect 33551 5729 33563 5732
rect 33505 5723 33563 5729
rect 33612 5701 33640 5732
rect 43070 5720 43076 5772
rect 43128 5720 43134 5772
rect 32493 5695 32551 5701
rect 32493 5692 32505 5695
rect 31720 5664 32505 5692
rect 31720 5652 31726 5664
rect 32493 5661 32505 5664
rect 32539 5661 32551 5695
rect 32493 5655 32551 5661
rect 32585 5695 32643 5701
rect 32585 5661 32597 5695
rect 32631 5661 32643 5695
rect 32585 5655 32643 5661
rect 33597 5695 33655 5701
rect 33597 5661 33609 5695
rect 33643 5661 33655 5695
rect 33597 5655 33655 5661
rect 37366 5652 37372 5704
rect 37424 5692 37430 5704
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 37424 5664 37841 5692
rect 37424 5652 37430 5664
rect 37829 5661 37841 5664
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 38010 5652 38016 5704
rect 38068 5652 38074 5704
rect 30374 5584 30380 5636
rect 30432 5584 30438 5636
rect 31220 5624 31248 5652
rect 32309 5627 32367 5633
rect 32309 5624 32321 5627
rect 31220 5596 32321 5624
rect 32309 5593 32321 5596
rect 32355 5593 32367 5627
rect 32309 5587 32367 5593
rect 43346 5584 43352 5636
rect 43404 5584 43410 5636
rect 43438 5584 43444 5636
rect 43496 5624 43502 5636
rect 43496 5596 43838 5624
rect 43496 5584 43502 5596
rect 33045 5559 33103 5565
rect 33045 5556 33057 5559
rect 29196 5528 33057 5556
rect 27212 5516 27218 5528
rect 33045 5525 33057 5528
rect 33091 5525 33103 5559
rect 33045 5519 33103 5525
rect 44818 5516 44824 5568
rect 44876 5516 44882 5568
rect 1104 5466 45172 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 45172 5466
rect 1104 5392 45172 5414
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 2740 5324 4016 5352
rect 2740 5312 2746 5324
rect 2501 5287 2559 5293
rect 2501 5253 2513 5287
rect 2547 5284 2559 5287
rect 2869 5287 2927 5293
rect 2869 5284 2881 5287
rect 2547 5256 2881 5284
rect 2547 5253 2559 5256
rect 2501 5247 2559 5253
rect 2869 5253 2881 5256
rect 2915 5253 2927 5287
rect 2869 5247 2927 5253
rect 3988 5216 4016 5324
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4212 5324 4445 5352
rect 4212 5312 4218 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 6914 5312 6920 5364
rect 6972 5312 6978 5364
rect 10042 5352 10048 5364
rect 8772 5324 10048 5352
rect 6932 5284 6960 5312
rect 8772 5293 8800 5324
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10468 5324 10885 5352
rect 10468 5312 10474 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 13688 5324 14381 5352
rect 13688 5312 13694 5324
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 14369 5315 14427 5321
rect 14553 5355 14611 5361
rect 14553 5321 14565 5355
rect 14599 5352 14611 5355
rect 14826 5352 14832 5364
rect 14599 5324 14832 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 20070 5352 20076 5364
rect 19812 5324 20076 5352
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 6932 5256 7021 5284
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 8757 5287 8815 5293
rect 8757 5253 8769 5287
rect 8803 5253 8815 5287
rect 8757 5247 8815 5253
rect 9582 5244 9588 5296
rect 9640 5244 9646 5296
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13964 5256 14197 5284
rect 13964 5244 13970 5256
rect 14185 5253 14197 5256
rect 14231 5284 14243 5287
rect 15562 5284 15568 5296
rect 14231 5256 15568 5284
rect 14231 5253 14243 5256
rect 14185 5247 14243 5253
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 19812 5293 19840 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 22572 5324 26280 5352
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5253 19855 5287
rect 19797 5247 19855 5253
rect 19978 5244 19984 5296
rect 20036 5284 20042 5296
rect 20036 5256 20286 5284
rect 20036 5244 20042 5256
rect 5442 5216 5448 5228
rect 3988 5202 5448 5216
rect 4002 5188 5448 5202
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 1854 5108 1860 5160
rect 1912 5108 1918 5160
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4387 5120 4997 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 9600 5148 9628 5244
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 10652 5188 10701 5216
rect 10652 5176 10658 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 12618 5216 12624 5228
rect 12207 5188 12624 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 10962 5148 10968 5160
rect 9600 5120 10968 5148
rect 4985 5111 5043 5117
rect 2608 5012 2636 5111
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11072 5148 11100 5179
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17092 5188 17509 5216
rect 17092 5176 17098 5188
rect 17497 5185 17509 5188
rect 17543 5216 17555 5219
rect 22005 5219 22063 5225
rect 17543 5188 20208 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 13170 5148 13176 5160
rect 11072 5120 13176 5148
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 19150 5148 19156 5160
rect 17635 5120 19156 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 20180 5148 20208 5188
rect 22005 5185 22017 5219
rect 22051 5216 22063 5219
rect 22186 5216 22192 5228
rect 22051 5188 22192 5216
rect 22051 5185 22063 5188
rect 22005 5179 22063 5185
rect 22186 5176 22192 5188
rect 22244 5176 22250 5228
rect 22572 5225 22600 5324
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 23477 5219 23535 5225
rect 23477 5185 23489 5219
rect 23523 5185 23535 5219
rect 23477 5179 23535 5185
rect 23753 5219 23811 5225
rect 23753 5185 23765 5219
rect 23799 5216 23811 5219
rect 23799 5188 24256 5216
rect 23799 5185 23811 5188
rect 23753 5179 23811 5185
rect 20806 5148 20812 5160
rect 20180 5120 20812 5148
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 21266 5108 21272 5160
rect 21324 5108 21330 5160
rect 21637 5151 21695 5157
rect 21637 5117 21649 5151
rect 21683 5148 21695 5151
rect 22094 5148 22100 5160
rect 21683 5120 22100 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 22094 5108 22100 5120
rect 22152 5148 22158 5160
rect 23290 5148 23296 5160
rect 22152 5120 23296 5148
rect 22152 5108 22158 5120
rect 23290 5108 23296 5120
rect 23348 5108 23354 5160
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18138 5080 18144 5092
rect 17911 5052 18144 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 23106 5040 23112 5092
rect 23164 5080 23170 5092
rect 23400 5080 23428 5179
rect 23492 5148 23520 5179
rect 23842 5148 23848 5160
rect 23492 5120 23848 5148
rect 23842 5108 23848 5120
rect 23900 5108 23906 5160
rect 23164 5052 23336 5080
rect 23400 5052 23796 5080
rect 23164 5040 23170 5052
rect 3234 5012 3240 5024
rect 2608 4984 3240 5012
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8895 5015 8953 5021
rect 8895 5012 8907 5015
rect 8352 4984 8907 5012
rect 8352 4972 8358 4984
rect 8895 4981 8907 4984
rect 8941 4981 8953 5015
rect 8895 4975 8953 4981
rect 11974 4972 11980 5024
rect 12032 4972 12038 5024
rect 14090 4972 14096 5024
rect 14148 5012 14154 5024
rect 14366 5012 14372 5024
rect 14148 4984 14372 5012
rect 14148 4972 14154 4984
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 20346 4972 20352 5024
rect 20404 5012 20410 5024
rect 21913 5015 21971 5021
rect 21913 5012 21925 5015
rect 20404 4984 21925 5012
rect 20404 4972 20410 4984
rect 21913 4981 21925 4984
rect 21959 4981 21971 5015
rect 21913 4975 21971 4981
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 23308 5012 23336 5052
rect 23768 5024 23796 5052
rect 24118 5040 24124 5092
rect 24176 5040 24182 5092
rect 24228 5080 24256 5188
rect 24302 5176 24308 5228
rect 24360 5216 24366 5228
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 24360 5188 24685 5216
rect 24360 5176 24366 5188
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 24765 5219 24823 5225
rect 24765 5185 24777 5219
rect 24811 5216 24823 5219
rect 24854 5216 24860 5228
rect 24811 5188 24860 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 24780 5080 24808 5179
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 25317 5219 25375 5225
rect 25317 5185 25329 5219
rect 25363 5185 25375 5219
rect 25317 5179 25375 5185
rect 24964 5148 24992 5179
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24964 5120 25145 5148
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 24228 5052 24808 5080
rect 24857 5083 24915 5089
rect 24857 5049 24869 5083
rect 24903 5080 24915 5083
rect 25222 5080 25228 5092
rect 24903 5052 25228 5080
rect 24903 5049 24915 5052
rect 24857 5043 24915 5049
rect 25222 5040 25228 5052
rect 25280 5040 25286 5092
rect 23661 5015 23719 5021
rect 23661 5012 23673 5015
rect 23308 4984 23673 5012
rect 23661 4981 23673 4984
rect 23707 4981 23719 5015
rect 23661 4975 23719 4981
rect 23750 4972 23756 5024
rect 23808 4972 23814 5024
rect 23842 4972 23848 5024
rect 23900 4972 23906 5024
rect 24136 5012 24164 5040
rect 24213 5015 24271 5021
rect 24213 5012 24225 5015
rect 24136 4984 24225 5012
rect 24213 4981 24225 4984
rect 24259 4981 24271 5015
rect 24213 4975 24271 4981
rect 24486 4972 24492 5024
rect 24544 4972 24550 5024
rect 25332 5012 25360 5179
rect 25406 5176 25412 5228
rect 25464 5216 25470 5228
rect 25777 5219 25835 5225
rect 25777 5216 25789 5219
rect 25464 5188 25789 5216
rect 25464 5176 25470 5188
rect 25777 5185 25789 5188
rect 25823 5185 25835 5219
rect 25777 5179 25835 5185
rect 26142 5176 26148 5228
rect 26200 5176 26206 5228
rect 25498 5108 25504 5160
rect 25556 5108 25562 5160
rect 25593 5151 25651 5157
rect 25593 5117 25605 5151
rect 25639 5148 25651 5151
rect 26160 5148 26188 5176
rect 25639 5120 26188 5148
rect 25639 5117 25651 5120
rect 25593 5111 25651 5117
rect 25409 5083 25467 5089
rect 25409 5049 25421 5083
rect 25455 5080 25467 5083
rect 25866 5080 25872 5092
rect 25455 5052 25872 5080
rect 25455 5049 25467 5052
rect 25409 5043 25467 5049
rect 25866 5040 25872 5052
rect 25924 5040 25930 5092
rect 25958 5040 25964 5092
rect 26016 5040 26022 5092
rect 25976 5012 26004 5040
rect 25332 4984 26004 5012
rect 26252 5012 26280 5324
rect 26970 5312 26976 5364
rect 27028 5352 27034 5364
rect 31297 5355 31355 5361
rect 27028 5324 29408 5352
rect 27028 5312 27034 5324
rect 29380 5284 29408 5324
rect 31297 5321 31309 5355
rect 31343 5352 31355 5355
rect 31570 5352 31576 5364
rect 31343 5324 31576 5352
rect 31343 5321 31355 5324
rect 31297 5315 31355 5321
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 35342 5312 35348 5364
rect 35400 5352 35406 5364
rect 38565 5355 38623 5361
rect 38565 5352 38577 5355
rect 35400 5324 38577 5352
rect 35400 5312 35406 5324
rect 38565 5321 38577 5324
rect 38611 5352 38623 5355
rect 38746 5352 38752 5364
rect 38611 5324 38752 5352
rect 38611 5321 38623 5324
rect 38565 5315 38623 5321
rect 38746 5312 38752 5324
rect 38804 5312 38810 5364
rect 41233 5355 41291 5361
rect 41233 5321 41245 5355
rect 41279 5352 41291 5355
rect 41322 5352 41328 5364
rect 41279 5324 41328 5352
rect 41279 5321 41291 5324
rect 41233 5315 41291 5321
rect 41322 5312 41328 5324
rect 41380 5312 41386 5364
rect 42150 5312 42156 5364
rect 42208 5352 42214 5364
rect 43165 5355 43223 5361
rect 42208 5324 42748 5352
rect 42208 5312 42214 5324
rect 29730 5284 29736 5296
rect 29380 5256 29736 5284
rect 29730 5244 29736 5256
rect 29788 5284 29794 5296
rect 30282 5284 30288 5296
rect 29788 5256 30288 5284
rect 29788 5244 29794 5256
rect 30282 5244 30288 5256
rect 30340 5244 30346 5296
rect 37274 5284 37280 5296
rect 31312 5256 37280 5284
rect 26970 5176 26976 5228
rect 27028 5216 27034 5228
rect 27065 5219 27123 5225
rect 27065 5216 27077 5219
rect 27028 5188 27077 5216
rect 27028 5176 27034 5188
rect 27065 5185 27077 5188
rect 27111 5185 27123 5219
rect 27065 5179 27123 5185
rect 31312 5160 31340 5256
rect 37274 5244 37280 5256
rect 37332 5244 37338 5296
rect 37384 5256 40066 5284
rect 42076 5256 42380 5284
rect 34606 5176 34612 5228
rect 34664 5216 34670 5228
rect 34701 5219 34759 5225
rect 34701 5216 34713 5219
rect 34664 5188 34713 5216
rect 34664 5176 34670 5188
rect 34701 5185 34713 5188
rect 34747 5185 34759 5219
rect 34701 5179 34759 5185
rect 34885 5219 34943 5225
rect 34885 5185 34897 5219
rect 34931 5216 34943 5219
rect 35434 5216 35440 5228
rect 34931 5188 35440 5216
rect 34931 5185 34943 5188
rect 34885 5179 34943 5185
rect 35434 5176 35440 5188
rect 35492 5176 35498 5228
rect 36357 5219 36415 5225
rect 36357 5216 36369 5219
rect 36004 5188 36369 5216
rect 29546 5108 29552 5160
rect 29604 5108 29610 5160
rect 29822 5108 29828 5160
rect 29880 5108 29886 5160
rect 31294 5108 31300 5160
rect 31352 5108 31358 5160
rect 36004 5148 36032 5188
rect 36357 5185 36369 5188
rect 36403 5216 36415 5219
rect 36538 5216 36544 5228
rect 36403 5188 36544 5216
rect 36403 5185 36415 5188
rect 36357 5179 36415 5185
rect 36538 5176 36544 5188
rect 36596 5176 36602 5228
rect 36722 5176 36728 5228
rect 36780 5216 36786 5228
rect 37384 5216 37412 5256
rect 36780 5188 37412 5216
rect 36780 5176 36786 5188
rect 38746 5176 38752 5228
rect 38804 5216 38810 5228
rect 39022 5216 39028 5228
rect 38804 5188 39028 5216
rect 38804 5176 38810 5188
rect 39022 5176 39028 5188
rect 39080 5216 39086 5228
rect 39206 5216 39212 5228
rect 39080 5188 39212 5216
rect 39080 5176 39086 5188
rect 39206 5176 39212 5188
rect 39264 5216 39270 5228
rect 41417 5219 41475 5225
rect 39264 5188 39344 5216
rect 39264 5176 39270 5188
rect 31726 5120 36032 5148
rect 27338 5040 27344 5092
rect 27396 5080 27402 5092
rect 28994 5080 29000 5092
rect 27396 5052 29000 5080
rect 27396 5040 27402 5052
rect 28994 5040 29000 5052
rect 29052 5040 29058 5092
rect 31726 5012 31754 5120
rect 36078 5108 36084 5160
rect 36136 5108 36142 5160
rect 39316 5157 39344 5188
rect 41417 5185 41429 5219
rect 41463 5216 41475 5219
rect 41506 5216 41512 5228
rect 41463 5188 41512 5216
rect 41463 5185 41475 5188
rect 41417 5179 41475 5185
rect 41506 5176 41512 5188
rect 41564 5176 41570 5228
rect 42076 5225 42104 5256
rect 41785 5219 41843 5225
rect 41785 5185 41797 5219
rect 41831 5185 41843 5219
rect 41785 5179 41843 5185
rect 41877 5219 41935 5225
rect 41877 5185 41889 5219
rect 41923 5216 41935 5219
rect 42061 5219 42119 5225
rect 42061 5216 42073 5219
rect 41923 5188 42073 5216
rect 41923 5185 41935 5188
rect 41877 5179 41935 5185
rect 42061 5185 42073 5188
rect 42107 5185 42119 5219
rect 42242 5216 42248 5228
rect 42061 5179 42119 5185
rect 42168 5188 42248 5216
rect 39301 5151 39359 5157
rect 39301 5117 39313 5151
rect 39347 5117 39359 5151
rect 39301 5111 39359 5117
rect 39574 5108 39580 5160
rect 39632 5108 39638 5160
rect 41046 5108 41052 5160
rect 41104 5148 41110 5160
rect 41800 5148 41828 5179
rect 41104 5120 41828 5148
rect 41104 5108 41110 5120
rect 36265 5083 36323 5089
rect 36265 5049 36277 5083
rect 36311 5080 36323 5083
rect 36446 5080 36452 5092
rect 36311 5052 36452 5080
rect 36311 5049 36323 5052
rect 36265 5043 36323 5049
rect 36446 5040 36452 5052
rect 36504 5040 36510 5092
rect 41690 5040 41696 5092
rect 41748 5080 41754 5092
rect 42168 5080 42196 5188
rect 42242 5176 42248 5188
rect 42300 5176 42306 5228
rect 41748 5052 42196 5080
rect 42352 5080 42380 5256
rect 42720 5157 42748 5324
rect 43165 5321 43177 5355
rect 43211 5352 43223 5355
rect 43346 5352 43352 5364
rect 43211 5324 43352 5352
rect 43211 5321 43223 5324
rect 43165 5315 43223 5321
rect 43346 5312 43352 5324
rect 43404 5312 43410 5364
rect 42797 5219 42855 5225
rect 42797 5185 42809 5219
rect 42843 5216 42855 5219
rect 43901 5219 43959 5225
rect 43901 5216 43913 5219
rect 42843 5188 43913 5216
rect 42843 5185 42855 5188
rect 42797 5179 42855 5185
rect 43901 5185 43913 5188
rect 43947 5185 43959 5219
rect 43901 5179 43959 5185
rect 42705 5151 42763 5157
rect 42705 5117 42717 5151
rect 42751 5117 42763 5151
rect 42705 5111 42763 5117
rect 42886 5108 42892 5160
rect 42944 5108 42950 5160
rect 44453 5151 44511 5157
rect 44453 5148 44465 5151
rect 42996 5120 44465 5148
rect 42904 5080 42932 5108
rect 42352 5052 42932 5080
rect 41748 5040 41754 5052
rect 42996 5024 43024 5120
rect 44453 5117 44465 5120
rect 44499 5148 44511 5151
rect 44818 5148 44824 5160
rect 44499 5120 44824 5148
rect 44499 5117 44511 5120
rect 44453 5111 44511 5117
rect 44818 5108 44824 5120
rect 44876 5108 44882 5160
rect 26252 4984 31754 5012
rect 34698 4972 34704 5024
rect 34756 4972 34762 5024
rect 36170 4972 36176 5024
rect 36228 4972 36234 5024
rect 41509 5015 41567 5021
rect 41509 4981 41521 5015
rect 41555 5012 41567 5015
rect 42978 5012 42984 5024
rect 41555 4984 42984 5012
rect 41555 4981 41567 4984
rect 41509 4975 41567 4981
rect 42978 4972 42984 4984
rect 43036 4972 43042 5024
rect 1104 4922 45172 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 45172 4922
rect 1104 4848 45172 4870
rect 1627 4811 1685 4817
rect 1627 4777 1639 4811
rect 1673 4808 1685 4811
rect 1854 4808 1860 4820
rect 1673 4780 1860 4808
rect 1673 4777 1685 4780
rect 1627 4771 1685 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10100 4780 17724 4808
rect 10100 4768 10106 4780
rect 13078 4749 13084 4752
rect 13035 4743 13084 4749
rect 13035 4709 13047 4743
rect 13081 4709 13084 4743
rect 13035 4703 13084 4709
rect 13078 4700 13084 4703
rect 13136 4700 13142 4752
rect 13170 4700 13176 4752
rect 13228 4700 13234 4752
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 3292 4644 3433 4672
rect 3292 4632 3298 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 8536 4644 9229 4672
rect 8536 4632 8542 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 10594 4672 10600 4684
rect 9217 4635 9275 4641
rect 9692 4644 10600 4672
rect 9692 4616 9720 4644
rect 10594 4632 10600 4644
rect 10652 4672 10658 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 10652 4644 11253 4672
rect 10652 4632 10658 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4672 11667 4675
rect 11974 4672 11980 4684
rect 11655 4644 11980 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13688 4644 13737 4672
rect 13688 4632 13694 4644
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 3050 4564 3056 4616
rect 3108 4564 3114 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8352 4576 8401 4604
rect 8352 4564 8358 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 9306 4564 9312 4616
rect 9364 4564 9370 4616
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 13596 4576 13676 4604
rect 13596 4564 13602 4576
rect 2682 4496 2688 4548
rect 2740 4496 2746 4548
rect 11974 4496 11980 4548
rect 12032 4496 12038 4548
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 7837 4471 7895 4477
rect 7837 4468 7849 4471
rect 7708 4440 7849 4468
rect 7708 4428 7714 4440
rect 7837 4437 7849 4440
rect 7883 4437 7895 4471
rect 7837 4431 7895 4437
rect 8938 4428 8944 4480
rect 8996 4428 9002 4480
rect 13538 4428 13544 4480
rect 13596 4428 13602 4480
rect 13648 4477 13676 4576
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 16850 4536 16856 4548
rect 16172 4508 16856 4536
rect 16172 4496 16178 4508
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 17696 4536 17724 4780
rect 20346 4768 20352 4820
rect 20404 4768 20410 4820
rect 21177 4811 21235 4817
rect 21177 4777 21189 4811
rect 21223 4808 21235 4811
rect 21266 4808 21272 4820
rect 21223 4780 21272 4808
rect 21223 4777 21235 4780
rect 21177 4771 21235 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 23198 4768 23204 4820
rect 23256 4768 23262 4820
rect 23566 4768 23572 4820
rect 23624 4768 23630 4820
rect 23753 4811 23811 4817
rect 23753 4777 23765 4811
rect 23799 4777 23811 4811
rect 23753 4771 23811 4777
rect 18690 4700 18696 4752
rect 18748 4740 18754 4752
rect 18785 4743 18843 4749
rect 18785 4740 18797 4743
rect 18748 4712 18797 4740
rect 18748 4700 18754 4712
rect 18785 4709 18797 4712
rect 18831 4709 18843 4743
rect 18785 4703 18843 4709
rect 18892 4712 19472 4740
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18693 4607 18751 4613
rect 18693 4604 18705 4607
rect 18012 4576 18705 4604
rect 18012 4564 18018 4576
rect 18693 4573 18705 4576
rect 18739 4604 18751 4607
rect 18892 4604 18920 4712
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4672 19027 4675
rect 19337 4675 19395 4681
rect 19337 4672 19349 4675
rect 19015 4644 19349 4672
rect 19015 4641 19027 4644
rect 18969 4635 19027 4641
rect 19337 4641 19349 4644
rect 19383 4641 19395 4675
rect 19337 4635 19395 4641
rect 18739 4576 18920 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19444 4613 19472 4712
rect 20364 4681 20392 4768
rect 20901 4743 20959 4749
rect 20901 4709 20913 4743
rect 20947 4709 20959 4743
rect 20901 4703 20959 4709
rect 20349 4675 20407 4681
rect 20349 4641 20361 4675
rect 20395 4641 20407 4675
rect 20349 4635 20407 4641
rect 20441 4675 20499 4681
rect 20441 4641 20453 4675
rect 20487 4672 20499 4675
rect 20806 4672 20812 4684
rect 20487 4644 20812 4672
rect 20487 4641 20499 4644
rect 20441 4635 20499 4641
rect 19245 4607 19303 4613
rect 19245 4604 19257 4607
rect 19208 4576 19257 4604
rect 19208 4564 19214 4576
rect 19245 4573 19257 4576
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20364 4604 20392 4635
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 19475 4576 20392 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20530 4564 20536 4616
rect 20588 4564 20594 4616
rect 20916 4604 20944 4703
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 22094 4672 22100 4684
rect 21867 4644 22100 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 22094 4632 22100 4644
rect 22152 4632 22158 4684
rect 22189 4675 22247 4681
rect 22189 4641 22201 4675
rect 22235 4672 22247 4675
rect 23216 4672 23244 4768
rect 23768 4684 23796 4771
rect 23842 4768 23848 4820
rect 23900 4768 23906 4820
rect 34698 4768 34704 4820
rect 34756 4768 34762 4820
rect 35700 4811 35758 4817
rect 35700 4777 35712 4811
rect 35746 4808 35758 4811
rect 36170 4808 36176 4820
rect 35746 4780 36176 4808
rect 35746 4777 35758 4780
rect 35700 4771 35758 4777
rect 36170 4768 36176 4780
rect 36228 4768 36234 4820
rect 37829 4811 37887 4817
rect 37829 4777 37841 4811
rect 37875 4808 37887 4811
rect 37918 4808 37924 4820
rect 37875 4780 37924 4808
rect 37875 4777 37887 4780
rect 37829 4771 37887 4777
rect 37918 4768 37924 4780
rect 37976 4768 37982 4820
rect 38010 4768 38016 4820
rect 38068 4768 38074 4820
rect 38473 4811 38531 4817
rect 38473 4777 38485 4811
rect 38519 4777 38531 4811
rect 38473 4771 38531 4777
rect 22235 4644 23244 4672
rect 22235 4641 22247 4644
rect 22189 4635 22247 4641
rect 23750 4632 23756 4684
rect 23808 4632 23814 4684
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20916 4576 21005 4604
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 21542 4564 21548 4616
rect 21600 4564 21606 4616
rect 23106 4564 23112 4616
rect 23164 4604 23170 4616
rect 23860 4604 23888 4768
rect 34716 4740 34744 4768
rect 38488 4740 38516 4771
rect 39574 4768 39580 4820
rect 39632 4808 39638 4820
rect 39945 4811 40003 4817
rect 39945 4808 39957 4811
rect 39632 4780 39957 4808
rect 39632 4768 39638 4780
rect 39945 4777 39957 4780
rect 39991 4777 40003 4811
rect 39945 4771 40003 4777
rect 40773 4811 40831 4817
rect 40773 4777 40785 4811
rect 40819 4808 40831 4811
rect 40862 4808 40868 4820
rect 40819 4780 40868 4808
rect 40819 4777 40831 4780
rect 40773 4771 40831 4777
rect 40862 4768 40868 4780
rect 40920 4768 40926 4820
rect 40957 4811 41015 4817
rect 40957 4777 40969 4811
rect 41003 4808 41015 4811
rect 41046 4808 41052 4820
rect 41003 4780 41052 4808
rect 41003 4777 41015 4780
rect 40957 4771 41015 4777
rect 41046 4768 41052 4780
rect 41104 4768 41110 4820
rect 42061 4811 42119 4817
rect 42061 4777 42073 4811
rect 42107 4808 42119 4811
rect 42150 4808 42156 4820
rect 42107 4780 42156 4808
rect 42107 4777 42119 4780
rect 42061 4771 42119 4777
rect 42150 4768 42156 4780
rect 42208 4768 42214 4820
rect 38746 4740 38752 4752
rect 34072 4712 34744 4740
rect 37384 4712 38752 4740
rect 33045 4675 33103 4681
rect 33045 4641 33057 4675
rect 33091 4672 33103 4675
rect 34072 4672 34100 4712
rect 33091 4644 34100 4672
rect 33091 4641 33103 4644
rect 33045 4635 33103 4641
rect 34514 4632 34520 4684
rect 34572 4672 34578 4684
rect 35342 4672 35348 4684
rect 34572 4644 35348 4672
rect 34572 4632 34578 4644
rect 35342 4632 35348 4644
rect 35400 4672 35406 4684
rect 35437 4675 35495 4681
rect 35437 4672 35449 4675
rect 35400 4644 35449 4672
rect 35400 4632 35406 4644
rect 35437 4641 35449 4644
rect 35483 4641 35495 4675
rect 35437 4635 35495 4641
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 23164 4576 23704 4604
rect 23860 4576 24041 4604
rect 23164 4564 23170 4576
rect 18601 4539 18659 4545
rect 18601 4536 18613 4539
rect 17696 4508 18613 4536
rect 18601 4505 18613 4508
rect 18647 4536 18659 4539
rect 21560 4536 21588 4564
rect 18647 4508 21588 4536
rect 22480 4508 22586 4536
rect 18647 4505 18659 4508
rect 18601 4499 18659 4505
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 16574 4468 16580 4480
rect 13679 4440 16580 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 18969 4471 19027 4477
rect 18969 4468 18981 4471
rect 18840 4440 18981 4468
rect 18840 4428 18846 4440
rect 18969 4437 18981 4440
rect 19015 4437 19027 4471
rect 18969 4431 19027 4437
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 22480 4468 22508 4508
rect 20036 4440 22508 4468
rect 23676 4468 23704 4576
rect 24029 4573 24041 4576
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 24854 4564 24860 4616
rect 24912 4564 24918 4616
rect 28534 4564 28540 4616
rect 28592 4604 28598 4616
rect 29546 4604 29552 4616
rect 28592 4576 29552 4604
rect 28592 4564 28598 4576
rect 29546 4564 29552 4576
rect 29604 4564 29610 4616
rect 31294 4564 31300 4616
rect 31352 4564 31358 4616
rect 32766 4564 32772 4616
rect 32824 4564 32830 4616
rect 37384 4613 37412 4712
rect 38746 4700 38752 4712
rect 38804 4740 38810 4752
rect 42245 4743 42303 4749
rect 38804 4712 39068 4740
rect 38804 4700 38810 4712
rect 38838 4632 38844 4684
rect 38896 4632 38902 4684
rect 39040 4681 39068 4712
rect 39592 4712 41920 4740
rect 39592 4684 39620 4712
rect 39025 4675 39083 4681
rect 39025 4641 39037 4675
rect 39071 4641 39083 4675
rect 39025 4635 39083 4641
rect 39574 4632 39580 4684
rect 39632 4632 39638 4684
rect 40313 4675 40371 4681
rect 40313 4672 40325 4675
rect 40144 4644 40325 4672
rect 35253 4607 35311 4613
rect 35253 4573 35265 4607
rect 35299 4573 35311 4607
rect 35253 4567 35311 4573
rect 37369 4607 37427 4613
rect 37369 4573 37381 4607
rect 37415 4573 37427 4607
rect 37369 4567 37427 4573
rect 37461 4607 37519 4613
rect 37461 4573 37473 4607
rect 37507 4573 37519 4607
rect 37461 4567 37519 4573
rect 23753 4539 23811 4545
rect 23753 4505 23765 4539
rect 23799 4536 23811 4539
rect 24872 4536 24900 4564
rect 23799 4508 24900 4536
rect 23799 4505 23811 4508
rect 23753 4499 23811 4505
rect 33778 4496 33784 4548
rect 33836 4496 33842 4548
rect 34701 4539 34759 4545
rect 34701 4536 34713 4539
rect 34348 4508 34713 4536
rect 23937 4471 23995 4477
rect 23937 4468 23949 4471
rect 23676 4440 23949 4468
rect 20036 4428 20042 4440
rect 23937 4437 23949 4440
rect 23983 4468 23995 4471
rect 25406 4468 25412 4480
rect 23983 4440 25412 4468
rect 23983 4437 23995 4440
rect 23937 4431 23995 4437
rect 25406 4428 25412 4440
rect 25464 4428 25470 4480
rect 33042 4428 33048 4480
rect 33100 4468 33106 4480
rect 34348 4468 34376 4508
rect 34701 4505 34713 4508
rect 34747 4505 34759 4539
rect 34701 4499 34759 4505
rect 33100 4440 34376 4468
rect 34517 4471 34575 4477
rect 33100 4428 33106 4440
rect 34517 4437 34529 4471
rect 34563 4468 34575 4471
rect 34606 4468 34612 4480
rect 34563 4440 34612 4468
rect 34563 4437 34575 4440
rect 34517 4431 34575 4437
rect 34606 4428 34612 4440
rect 34664 4468 34670 4480
rect 35268 4468 35296 4567
rect 36722 4496 36728 4548
rect 36780 4496 36786 4548
rect 37476 4536 37504 4567
rect 37826 4564 37832 4616
rect 37884 4564 37890 4616
rect 38856 4604 38884 4632
rect 39853 4607 39911 4613
rect 39853 4604 39865 4607
rect 38856 4576 39865 4604
rect 39853 4573 39865 4576
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 40034 4564 40040 4616
rect 40092 4564 40098 4616
rect 40144 4613 40172 4644
rect 40313 4641 40325 4644
rect 40359 4672 40371 4675
rect 40359 4644 41276 4672
rect 40359 4641 40371 4644
rect 40313 4635 40371 4641
rect 40129 4607 40187 4613
rect 40129 4573 40141 4607
rect 40175 4573 40187 4607
rect 40129 4567 40187 4573
rect 40497 4607 40555 4613
rect 40497 4573 40509 4607
rect 40543 4573 40555 4607
rect 40497 4567 40555 4573
rect 40681 4607 40739 4613
rect 40681 4573 40693 4607
rect 40727 4604 40739 4607
rect 41046 4604 41052 4616
rect 40727 4576 41052 4604
rect 40727 4573 40739 4576
rect 40681 4567 40739 4573
rect 37200 4508 37504 4536
rect 37200 4480 37228 4508
rect 38010 4496 38016 4548
rect 38068 4536 38074 4548
rect 38289 4539 38347 4545
rect 38289 4536 38301 4539
rect 38068 4508 38301 4536
rect 38068 4496 38074 4508
rect 38289 4505 38301 4508
rect 38335 4505 38347 4539
rect 38289 4499 38347 4505
rect 38672 4508 39804 4536
rect 34664 4440 35296 4468
rect 34664 4428 34670 4440
rect 36538 4428 36544 4480
rect 36596 4468 36602 4480
rect 37182 4468 37188 4480
rect 36596 4440 37188 4468
rect 36596 4428 36602 4440
rect 37182 4428 37188 4440
rect 37240 4428 37246 4480
rect 38194 4428 38200 4480
rect 38252 4468 38258 4480
rect 38672 4477 38700 4508
rect 38489 4471 38547 4477
rect 38489 4468 38501 4471
rect 38252 4440 38501 4468
rect 38252 4428 38258 4440
rect 38489 4437 38501 4440
rect 38535 4437 38547 4471
rect 38489 4431 38547 4437
rect 38657 4471 38715 4477
rect 38657 4437 38669 4471
rect 38703 4437 38715 4471
rect 38657 4431 38715 4437
rect 39298 4428 39304 4480
rect 39356 4468 39362 4480
rect 39669 4471 39727 4477
rect 39669 4468 39681 4471
rect 39356 4440 39681 4468
rect 39356 4428 39362 4440
rect 39669 4437 39681 4440
rect 39715 4437 39727 4471
rect 39776 4468 39804 4508
rect 40512 4468 40540 4567
rect 41046 4564 41052 4576
rect 41104 4564 41110 4616
rect 41248 4613 41276 4644
rect 41233 4607 41291 4613
rect 41233 4573 41245 4607
rect 41279 4573 41291 4607
rect 41233 4567 41291 4573
rect 41322 4564 41328 4616
rect 41380 4564 41386 4616
rect 41414 4564 41420 4616
rect 41472 4564 41478 4616
rect 40770 4496 40776 4548
rect 40828 4536 40834 4548
rect 41141 4539 41199 4545
rect 40828 4508 41092 4536
rect 40828 4496 40834 4508
rect 40678 4468 40684 4480
rect 39776 4440 40684 4468
rect 39669 4431 39727 4437
rect 40678 4428 40684 4440
rect 40736 4468 40742 4480
rect 40931 4471 40989 4477
rect 40931 4468 40943 4471
rect 40736 4440 40943 4468
rect 40736 4428 40742 4440
rect 40931 4437 40943 4440
rect 40977 4437 40989 4471
rect 41064 4468 41092 4508
rect 41141 4505 41153 4539
rect 41187 4536 41199 4539
rect 41506 4536 41512 4548
rect 41187 4508 41512 4536
rect 41187 4505 41199 4508
rect 41141 4499 41199 4505
rect 41506 4496 41512 4508
rect 41564 4536 41570 4548
rect 41892 4545 41920 4712
rect 42245 4709 42257 4743
rect 42291 4709 42303 4743
rect 42245 4703 42303 4709
rect 42260 4672 42288 4703
rect 42260 4644 43024 4672
rect 42242 4564 42248 4616
rect 42300 4604 42306 4616
rect 42996 4613 43024 4644
rect 42686 4607 42744 4613
rect 42300 4600 42656 4604
rect 42686 4600 42698 4607
rect 42300 4576 42698 4600
rect 42300 4564 42306 4576
rect 42628 4573 42698 4576
rect 42732 4604 42744 4607
rect 42981 4607 43039 4613
rect 42732 4573 42748 4604
rect 42628 4572 42748 4573
rect 42981 4573 42993 4607
rect 43027 4573 43039 4607
rect 42686 4567 42744 4572
rect 42981 4567 43039 4573
rect 41877 4539 41935 4545
rect 41564 4508 41828 4536
rect 41564 4496 41570 4508
rect 41690 4468 41696 4480
rect 41064 4440 41696 4468
rect 40931 4431 40989 4437
rect 41690 4428 41696 4440
rect 41748 4428 41754 4480
rect 41800 4468 41828 4508
rect 41877 4505 41889 4539
rect 41923 4505 41935 4539
rect 41877 4499 41935 4505
rect 41966 4496 41972 4548
rect 42024 4496 42030 4548
rect 42093 4539 42151 4545
rect 42093 4505 42105 4539
rect 42139 4536 42151 4539
rect 42337 4539 42395 4545
rect 42337 4536 42349 4539
rect 42139 4508 42349 4536
rect 42139 4505 42151 4508
rect 42093 4499 42151 4505
rect 42337 4505 42349 4508
rect 42383 4505 42395 4539
rect 42337 4499 42395 4505
rect 42521 4539 42579 4545
rect 42521 4505 42533 4539
rect 42567 4536 42579 4539
rect 42886 4536 42892 4548
rect 42567 4508 42892 4536
rect 42567 4505 42579 4508
rect 42521 4499 42579 4505
rect 42886 4496 42892 4508
rect 42944 4536 42950 4548
rect 43162 4536 43168 4548
rect 42944 4508 43168 4536
rect 42944 4496 42950 4508
rect 43162 4496 43168 4508
rect 43220 4496 43226 4548
rect 41984 4468 42012 4496
rect 41800 4440 42012 4468
rect 42794 4428 42800 4480
rect 42852 4428 42858 4480
rect 1104 4378 45172 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 45172 4378
rect 1104 4304 45172 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3108 4236 3801 4264
rect 3108 4224 3114 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 3789 4227 3847 4233
rect 12618 4224 12624 4276
rect 12676 4224 12682 4276
rect 19150 4224 19156 4276
rect 19208 4264 19214 4276
rect 20162 4264 20168 4276
rect 19208 4236 20168 4264
rect 19208 4224 19214 4236
rect 20162 4224 20168 4236
rect 20220 4264 20226 4276
rect 20220 4236 20300 4264
rect 20220 4224 20226 4236
rect 7282 4156 7288 4208
rect 7340 4156 7346 4208
rect 9674 4196 9680 4208
rect 9324 4168 9680 4196
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 6178 4128 6184 4140
rect 3292 4100 6184 4128
rect 3292 4088 3298 4100
rect 6178 4088 6184 4100
rect 6236 4128 6242 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6236 4100 6377 4128
rect 6236 4088 6242 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 9324 4137 9352 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 10962 4196 10968 4208
rect 10810 4168 10968 4196
rect 10962 4156 10968 4168
rect 11020 4196 11026 4208
rect 11974 4196 11980 4208
rect 11020 4168 11980 4196
rect 11020 4156 11026 4168
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 14108 4168 15056 4196
rect 14108 4140 14136 4168
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 8036 4100 9321 4128
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4614 4060 4620 4072
rect 4479 4032 4620 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 5534 4020 5540 4072
rect 5592 4020 5598 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7668 4060 7696 4088
rect 8036 4072 8064 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 15028 4137 15056 4168
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 16761 4199 16819 4205
rect 16761 4196 16773 4199
rect 15620 4168 16773 4196
rect 15620 4156 15626 4168
rect 16316 4140 16344 4168
rect 16761 4165 16773 4168
rect 16807 4165 16819 4199
rect 16761 4159 16819 4165
rect 18509 4199 18567 4205
rect 18509 4165 18521 4199
rect 18555 4196 18567 4199
rect 18782 4196 18788 4208
rect 18555 4168 18788 4196
rect 18555 4165 18567 4168
rect 18509 4159 18567 4165
rect 18782 4156 18788 4168
rect 18840 4156 18846 4208
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 6687 4032 7696 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8159 4032 8769 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11103 4032 12081 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12584 4032 13093 4060
rect 12584 4020 12590 4032
rect 13081 4029 13093 4032
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13630 4060 13636 4072
rect 13311 4032 13636 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8938 3992 8944 4004
rect 7800 3964 8944 3992
rect 7800 3952 7806 3964
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 14200 3992 14228 4091
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 16632 4100 17417 4128
rect 16632 4088 16638 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 19978 4128 19984 4140
rect 19668 4100 19984 4128
rect 19668 4088 19674 4100
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20272 4137 20300 4236
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 34238 4264 34244 4276
rect 29052 4236 29960 4264
rect 29052 4224 29058 4236
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 25590 4088 25596 4140
rect 25648 4088 25654 4140
rect 26050 4088 26056 4140
rect 26108 4128 26114 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26108 4100 26985 4128
rect 26108 4088 26114 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 27062 4088 27068 4140
rect 27120 4128 27126 4140
rect 27433 4131 27491 4137
rect 27433 4128 27445 4131
rect 27120 4100 27445 4128
rect 27120 4088 27126 4100
rect 27433 4097 27445 4100
rect 27479 4097 27491 4131
rect 29932 4128 29960 4236
rect 33152 4236 34244 4264
rect 32214 4128 32220 4140
rect 29932 4114 32220 4128
rect 29946 4100 32220 4114
rect 27433 4091 27491 4097
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 14332 4032 17509 4060
rect 14332 4020 14338 4032
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 14200 3964 14688 3992
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 6052 3896 6193 3924
rect 6052 3884 6058 3896
rect 6181 3893 6193 3896
rect 6227 3893 6239 3927
rect 6181 3887 6239 3893
rect 8202 3884 8208 3936
rect 8260 3884 8266 3936
rect 11514 3884 11520 3936
rect 11572 3884 11578 3936
rect 14550 3884 14556 3936
rect 14608 3884 14614 3936
rect 14660 3924 14688 3964
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 15194 3992 15200 4004
rect 14884 3964 15200 3992
rect 14884 3952 14890 3964
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 17512 3992 17540 4023
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 18104 4032 18245 4060
rect 18104 4020 18110 4032
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 18233 4023 18291 4029
rect 18340 4032 20177 4060
rect 18340 3992 18368 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20165 4023 20223 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20625 4063 20683 4069
rect 20625 4060 20637 4063
rect 20588 4032 20637 4060
rect 20588 4020 20594 4032
rect 20625 4029 20637 4032
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 28534 4020 28540 4072
rect 28592 4020 28598 4072
rect 28810 4020 28816 4072
rect 28868 4020 28874 4072
rect 30285 4063 30343 4069
rect 30285 4029 30297 4063
rect 30331 4060 30343 4063
rect 31386 4060 31392 4072
rect 30331 4032 31392 4060
rect 30331 4029 30343 4032
rect 30285 4023 30343 4029
rect 31386 4020 31392 4032
rect 31444 4020 31450 4072
rect 17512 3964 18368 3992
rect 19518 3952 19524 4004
rect 19576 3992 19582 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19576 3964 19993 3992
rect 19576 3952 19582 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 31864 3936 31892 4100
rect 32214 4088 32220 4100
rect 32272 4088 32278 4140
rect 32953 4131 33011 4137
rect 32953 4097 32965 4131
rect 32999 4128 33011 4131
rect 33042 4128 33048 4140
rect 32999 4100 33048 4128
rect 32999 4097 33011 4100
rect 32953 4091 33011 4097
rect 33042 4088 33048 4100
rect 33100 4088 33106 4140
rect 33152 4137 33180 4236
rect 34238 4224 34244 4236
rect 34296 4224 34302 4276
rect 34698 4264 34704 4276
rect 34440 4236 34704 4264
rect 34440 4205 34468 4236
rect 34698 4224 34704 4236
rect 34756 4224 34762 4276
rect 34885 4267 34943 4273
rect 34885 4233 34897 4267
rect 34931 4264 34943 4267
rect 35434 4264 35440 4276
rect 34931 4236 35440 4264
rect 34931 4233 34943 4236
rect 34885 4227 34943 4233
rect 35434 4224 35440 4236
rect 35492 4224 35498 4276
rect 36515 4267 36573 4273
rect 36515 4264 36527 4267
rect 36004 4236 36527 4264
rect 34425 4199 34483 4205
rect 34425 4165 34437 4199
rect 34471 4165 34483 4199
rect 34425 4159 34483 4165
rect 34532 4168 35388 4196
rect 33137 4131 33195 4137
rect 33137 4097 33149 4131
rect 33183 4097 33195 4131
rect 33137 4091 33195 4097
rect 34146 4088 34152 4140
rect 34204 4088 34210 4140
rect 34238 4088 34244 4140
rect 34296 4128 34302 4140
rect 34532 4128 34560 4168
rect 34296 4100 34560 4128
rect 34296 4088 34302 4100
rect 34606 4088 34612 4140
rect 34664 4088 34670 4140
rect 34716 4137 34744 4168
rect 35360 4137 35388 4168
rect 34701 4131 34759 4137
rect 34701 4097 34713 4131
rect 34747 4097 34759 4131
rect 34701 4091 34759 4097
rect 35161 4131 35219 4137
rect 35161 4097 35173 4131
rect 35207 4097 35219 4131
rect 35161 4091 35219 4097
rect 35345 4131 35403 4137
rect 35345 4097 35357 4131
rect 35391 4097 35403 4131
rect 35452 4128 35480 4224
rect 35894 4128 35900 4140
rect 35452 4100 35900 4128
rect 35345 4091 35403 4097
rect 33873 4063 33931 4069
rect 33873 4029 33885 4063
rect 33919 4060 33931 4063
rect 33962 4060 33968 4072
rect 33919 4032 33968 4060
rect 33919 4029 33931 4032
rect 33873 4023 33931 4029
rect 33962 4020 33968 4032
rect 34020 4060 34026 4072
rect 34333 4063 34391 4069
rect 34020 4032 34192 4060
rect 34020 4020 34026 4032
rect 33137 3995 33195 4001
rect 33137 3961 33149 3995
rect 33183 3992 33195 3995
rect 34054 3992 34060 4004
rect 33183 3964 34060 3992
rect 33183 3961 33195 3964
rect 33137 3955 33195 3961
rect 34054 3952 34060 3964
rect 34112 3952 34118 4004
rect 34164 3936 34192 4032
rect 34333 4029 34345 4063
rect 34379 4060 34391 4063
rect 34624 4060 34652 4088
rect 34379 4032 34652 4060
rect 34379 4029 34391 4032
rect 34333 4023 34391 4029
rect 35176 3992 35204 4091
rect 35360 4060 35388 4091
rect 35894 4088 35900 4100
rect 35952 4128 35958 4140
rect 36004 4137 36032 4236
rect 36515 4233 36527 4236
rect 36561 4233 36573 4267
rect 36515 4227 36573 4233
rect 36630 4224 36636 4276
rect 36688 4264 36694 4276
rect 37277 4267 37335 4273
rect 37277 4264 37289 4267
rect 36688 4236 37289 4264
rect 36688 4224 36694 4236
rect 37277 4233 37289 4236
rect 37323 4233 37335 4267
rect 37277 4227 37335 4233
rect 37826 4224 37832 4276
rect 37884 4224 37890 4276
rect 38657 4267 38715 4273
rect 38657 4233 38669 4267
rect 38703 4264 38715 4267
rect 38746 4264 38752 4276
rect 38703 4236 38752 4264
rect 38703 4233 38715 4236
rect 38657 4227 38715 4233
rect 38746 4224 38752 4236
rect 38804 4224 38810 4276
rect 40034 4224 40040 4276
rect 40092 4264 40098 4276
rect 40865 4267 40923 4273
rect 40865 4264 40877 4267
rect 40092 4236 40877 4264
rect 40092 4224 40098 4236
rect 40865 4233 40877 4236
rect 40911 4233 40923 4267
rect 40865 4227 40923 4233
rect 41414 4224 41420 4276
rect 41472 4264 41478 4276
rect 41601 4267 41659 4273
rect 41601 4264 41613 4267
rect 41472 4236 41613 4264
rect 41472 4224 41478 4236
rect 41601 4233 41613 4236
rect 41647 4233 41659 4267
rect 43438 4264 43444 4276
rect 41601 4227 41659 4233
rect 43088 4236 43444 4264
rect 36170 4156 36176 4208
rect 36228 4196 36234 4208
rect 36265 4199 36323 4205
rect 36265 4196 36277 4199
rect 36228 4168 36277 4196
rect 36228 4156 36234 4168
rect 36265 4165 36277 4168
rect 36311 4165 36323 4199
rect 36265 4159 36323 4165
rect 36725 4199 36783 4205
rect 36725 4165 36737 4199
rect 36771 4196 36783 4199
rect 37182 4196 37188 4208
rect 36771 4168 37188 4196
rect 36771 4165 36783 4168
rect 36725 4159 36783 4165
rect 35989 4131 36047 4137
rect 35989 4128 36001 4131
rect 35952 4100 36001 4128
rect 35952 4088 35958 4100
rect 35989 4097 36001 4100
rect 36035 4097 36047 4131
rect 35989 4091 36047 4097
rect 36081 4131 36139 4137
rect 36081 4097 36093 4131
rect 36127 4128 36139 4131
rect 36740 4128 36768 4159
rect 37182 4156 37188 4168
rect 37240 4196 37246 4208
rect 37844 4196 37872 4224
rect 40129 4199 40187 4205
rect 37240 4168 37872 4196
rect 38304 4168 38962 4196
rect 37240 4156 37246 4168
rect 36127 4100 36768 4128
rect 36909 4131 36967 4137
rect 36127 4097 36139 4100
rect 36081 4091 36139 4097
rect 36909 4097 36921 4131
rect 36955 4097 36967 4131
rect 36909 4091 36967 4097
rect 35710 4060 35716 4072
rect 35360 4032 35716 4060
rect 35710 4020 35716 4032
rect 35768 4020 35774 4072
rect 36446 4020 36452 4072
rect 36504 4060 36510 4072
rect 36924 4060 36952 4091
rect 37090 4088 37096 4140
rect 37148 4088 37154 4140
rect 38194 4128 38200 4140
rect 37200 4100 38200 4128
rect 37200 4060 37228 4100
rect 38194 4088 38200 4100
rect 38252 4088 38258 4140
rect 36504 4032 37228 4060
rect 36504 4020 36510 4032
rect 37274 4020 37280 4072
rect 37332 4060 37338 4072
rect 37829 4063 37887 4069
rect 37829 4060 37841 4063
rect 37332 4032 37841 4060
rect 37332 4020 37338 4032
rect 37829 4029 37841 4032
rect 37875 4029 37887 4063
rect 37829 4023 37887 4029
rect 38010 4020 38016 4072
rect 38068 4020 38074 4072
rect 34532 3964 35204 3992
rect 34532 3936 34560 3964
rect 36078 3952 36084 4004
rect 36136 3992 36142 4004
rect 36265 3995 36323 4001
rect 36265 3992 36277 3995
rect 36136 3964 36277 3992
rect 36136 3952 36142 3964
rect 36265 3961 36277 3964
rect 36311 3961 36323 3995
rect 36265 3955 36323 3961
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 14660 3896 17049 3924
rect 17037 3893 17049 3896
rect 17083 3924 17095 3927
rect 17402 3924 17408 3936
rect 17083 3896 17408 3924
rect 17083 3893 17095 3896
rect 17037 3887 17095 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17681 3927 17739 3933
rect 17681 3893 17693 3927
rect 17727 3924 17739 3927
rect 18690 3924 18696 3936
rect 17727 3896 18696 3924
rect 17727 3893 17739 3896
rect 17681 3887 17739 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 25774 3884 25780 3936
rect 25832 3884 25838 3936
rect 27154 3884 27160 3936
rect 27212 3884 27218 3936
rect 27249 3927 27307 3933
rect 27249 3893 27261 3927
rect 27295 3924 27307 3927
rect 27338 3924 27344 3936
rect 27295 3896 27344 3924
rect 27295 3893 27307 3896
rect 27249 3887 27307 3893
rect 27338 3884 27344 3896
rect 27396 3884 27402 3936
rect 31846 3884 31852 3936
rect 31904 3884 31910 3936
rect 33226 3884 33232 3936
rect 33284 3884 33290 3936
rect 33962 3884 33968 3936
rect 34020 3884 34026 3936
rect 34146 3884 34152 3936
rect 34204 3884 34210 3936
rect 34422 3884 34428 3936
rect 34480 3884 34486 3936
rect 34514 3884 34520 3936
rect 34572 3884 34578 3936
rect 35161 3927 35219 3933
rect 35161 3893 35173 3927
rect 35207 3924 35219 3927
rect 35526 3924 35532 3936
rect 35207 3896 35532 3924
rect 35207 3893 35219 3896
rect 35161 3887 35219 3893
rect 35526 3884 35532 3896
rect 35584 3884 35590 3936
rect 36357 3927 36415 3933
rect 36357 3893 36369 3927
rect 36403 3924 36415 3927
rect 36464 3924 36492 4020
rect 36722 3952 36728 4004
rect 36780 3952 36786 4004
rect 36906 3952 36912 4004
rect 36964 3952 36970 4004
rect 36403 3896 36492 3924
rect 36403 3893 36415 3896
rect 36357 3887 36415 3893
rect 36538 3884 36544 3936
rect 36596 3884 36602 3936
rect 36740 3924 36768 3952
rect 38304 3924 38332 4168
rect 40129 4165 40141 4199
rect 40175 4196 40187 4199
rect 43088 4196 43116 4236
rect 43438 4224 43444 4236
rect 43496 4224 43502 4276
rect 40175 4168 40632 4196
rect 40175 4165 40187 4168
rect 40129 4159 40187 4165
rect 40494 4088 40500 4140
rect 40552 4088 40558 4140
rect 40604 4137 40632 4168
rect 42352 4168 43194 4196
rect 42352 4140 42380 4168
rect 40589 4131 40647 4137
rect 40589 4097 40601 4131
rect 40635 4097 40647 4131
rect 40589 4091 40647 4097
rect 40678 4088 40684 4140
rect 40736 4128 40742 4140
rect 40773 4131 40831 4137
rect 40773 4128 40785 4131
rect 40736 4100 40785 4128
rect 40736 4088 40742 4100
rect 40773 4097 40785 4100
rect 40819 4097 40831 4131
rect 40773 4091 40831 4097
rect 40862 4088 40868 4140
rect 40920 4088 40926 4140
rect 40954 4088 40960 4140
rect 41012 4088 41018 4140
rect 41049 4131 41107 4137
rect 41049 4097 41061 4131
rect 41095 4097 41107 4131
rect 41049 4091 41107 4097
rect 41233 4131 41291 4137
rect 41233 4097 41245 4131
rect 41279 4128 41291 4131
rect 41322 4128 41328 4140
rect 41279 4100 41328 4128
rect 41279 4097 41291 4100
rect 41233 4091 41291 4097
rect 39114 4020 39120 4072
rect 39172 4060 39178 4072
rect 40405 4063 40463 4069
rect 40405 4060 40417 4063
rect 39172 4032 40417 4060
rect 39172 4020 39178 4032
rect 40405 4029 40417 4032
rect 40451 4029 40463 4063
rect 40880 4060 40908 4088
rect 41064 4060 41092 4091
rect 41322 4088 41328 4100
rect 41380 4088 41386 4140
rect 42334 4088 42340 4140
rect 42392 4088 42398 4140
rect 40880 4032 41092 4060
rect 40405 4023 40463 4029
rect 42058 4020 42064 4072
rect 42116 4060 42122 4072
rect 42153 4063 42211 4069
rect 42153 4060 42165 4063
rect 42116 4032 42165 4060
rect 42116 4020 42122 4032
rect 42153 4029 42165 4032
rect 42199 4029 42211 4063
rect 42153 4023 42211 4029
rect 42429 4063 42487 4069
rect 42429 4029 42441 4063
rect 42475 4029 42487 4063
rect 42429 4023 42487 4029
rect 42705 4063 42763 4069
rect 42705 4029 42717 4063
rect 42751 4060 42763 4063
rect 42794 4060 42800 4072
rect 42751 4032 42800 4060
rect 42751 4029 42763 4032
rect 42705 4023 42763 4029
rect 36740 3896 38332 3924
rect 38378 3884 38384 3936
rect 38436 3884 38442 3936
rect 41230 3884 41236 3936
rect 41288 3884 41294 3936
rect 42444 3924 42472 4023
rect 42794 4020 42800 4032
rect 42852 4020 42858 4072
rect 43162 4020 43168 4072
rect 43220 4060 43226 4072
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 43220 4032 44189 4060
rect 43220 4020 43226 4032
rect 44177 4029 44189 4032
rect 44223 4029 44235 4063
rect 44177 4023 44235 4029
rect 43070 3924 43076 3936
rect 42444 3896 43076 3924
rect 43070 3884 43076 3896
rect 43128 3884 43134 3936
rect 1104 3834 45172 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 45172 3834
rect 1104 3760 45172 3782
rect 7742 3720 7748 3732
rect 5460 3692 7748 3720
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 3881 3587 3939 3593
rect 3881 3584 3893 3587
rect 3292 3556 3893 3584
rect 3292 3544 3298 3556
rect 3881 3553 3893 3556
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 5460 3584 5488 3692
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 7947 3723 8005 3729
rect 7947 3689 7959 3723
rect 7993 3720 8005 3723
rect 8202 3720 8208 3732
rect 7993 3692 8208 3720
rect 7993 3689 8005 3692
rect 7947 3683 8005 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9306 3720 9312 3732
rect 8987 3692 9312 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9582 3680 9588 3732
rect 9640 3680 9646 3732
rect 10612 3692 12940 3720
rect 10612 3652 10640 3692
rect 9324 3624 10640 3652
rect 12912 3652 12940 3692
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 16298 3729 16304 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 13044 3692 13185 3720
rect 13044 3680 13050 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 16255 3723 16304 3729
rect 16255 3689 16267 3723
rect 16301 3689 16304 3723
rect 16255 3683 16304 3689
rect 16298 3680 16304 3683
rect 16356 3680 16362 3732
rect 19610 3720 19616 3732
rect 16684 3692 19616 3720
rect 12912 3624 14320 3652
rect 4295 3556 5488 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 5534 3544 5540 3596
rect 5592 3544 5598 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 5442 3516 5448 3528
rect 5276 3488 5448 3516
rect 5276 3434 5304 3488
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5552 3448 5580 3544
rect 5675 3451 5733 3457
rect 5675 3448 5687 3451
rect 5552 3420 5687 3448
rect 5675 3417 5687 3420
rect 5721 3417 5733 3451
rect 5675 3411 5733 3417
rect 7282 3408 7288 3460
rect 7340 3408 7346 3460
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 8018 3448 8024 3460
rect 7708 3420 8024 3448
rect 7708 3408 7714 3420
rect 8018 3408 8024 3420
rect 8076 3448 8082 3460
rect 8220 3448 8248 3547
rect 9324 3525 9352 3624
rect 12912 3596 12940 3624
rect 14292 3596 14320 3624
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3584 9459 3587
rect 9582 3584 9588 3596
rect 9447 3556 9588 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 9582 3544 9588 3556
rect 9640 3584 9646 3596
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9640 3556 10149 3584
rect 9640 3544 9646 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10594 3544 10600 3596
rect 10652 3544 10658 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11514 3584 11520 3596
rect 11011 3556 11520 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 12894 3544 12900 3596
rect 12952 3544 12958 3596
rect 14090 3544 14096 3596
rect 14148 3544 14154 3596
rect 14274 3544 14280 3596
rect 14332 3544 14338 3596
rect 16684 3584 16712 3692
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 24486 3680 24492 3732
rect 24544 3680 24550 3732
rect 25774 3680 25780 3732
rect 25832 3720 25838 3732
rect 26770 3723 26828 3729
rect 26770 3720 26782 3723
rect 25832 3692 26782 3720
rect 25832 3680 25838 3692
rect 26770 3689 26782 3692
rect 26816 3689 26828 3723
rect 28534 3720 28540 3732
rect 26770 3683 26828 3689
rect 28184 3692 28540 3720
rect 24504 3652 24532 3680
rect 23952 3624 24532 3652
rect 14660 3556 16712 3584
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 12802 3476 12808 3528
rect 12860 3476 12866 3528
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 8076 3420 8248 3448
rect 8076 3408 8082 3420
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6914 3380 6920 3392
rect 6503 3352 6920 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 9784 3380 9812 3476
rect 11974 3408 11980 3460
rect 12032 3408 12038 3460
rect 14660 3448 14688 3556
rect 16114 3476 16120 3528
rect 16172 3476 16178 3528
rect 12268 3434 14688 3448
rect 15841 3451 15899 3457
rect 12268 3420 14674 3434
rect 12268 3380 12296 3420
rect 15841 3417 15853 3451
rect 15887 3417 15899 3451
rect 16684 3434 16712 3556
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 18046 3584 18052 3596
rect 16908 3556 18052 3584
rect 16908 3544 16914 3556
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18601 3587 18659 3593
rect 18601 3553 18613 3587
rect 18647 3584 18659 3587
rect 18690 3584 18696 3596
rect 18647 3556 18696 3584
rect 18647 3553 18659 3556
rect 18601 3547 18659 3553
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 23952 3593 23980 3624
rect 23937 3587 23995 3593
rect 23937 3553 23949 3587
rect 23983 3553 23995 3587
rect 23937 3547 23995 3553
rect 24397 3587 24455 3593
rect 24397 3553 24409 3587
rect 24443 3584 24455 3587
rect 25682 3584 25688 3596
rect 24443 3556 25688 3584
rect 24443 3553 24455 3556
rect 24397 3547 24455 3553
rect 25682 3544 25688 3556
rect 25740 3584 25746 3596
rect 26510 3584 26516 3596
rect 25740 3556 26516 3584
rect 25740 3544 25746 3556
rect 26510 3544 26516 3556
rect 26568 3584 26574 3596
rect 28184 3584 28212 3692
rect 28534 3680 28540 3692
rect 28592 3720 28598 3732
rect 28592 3692 28672 3720
rect 28592 3680 28598 3692
rect 28261 3655 28319 3661
rect 28261 3621 28273 3655
rect 28307 3652 28319 3655
rect 28307 3624 28580 3652
rect 28307 3621 28319 3624
rect 28261 3615 28319 3621
rect 28552 3593 28580 3624
rect 26568 3556 28212 3584
rect 28537 3587 28595 3593
rect 26568 3544 26574 3556
rect 28537 3553 28549 3587
rect 28583 3553 28595 3587
rect 28644 3584 28672 3692
rect 28810 3680 28816 3732
rect 28868 3720 28874 3732
rect 29181 3723 29239 3729
rect 29181 3720 29193 3723
rect 28868 3692 29193 3720
rect 28868 3680 28874 3692
rect 29181 3689 29193 3692
rect 29227 3689 29239 3723
rect 29181 3683 29239 3689
rect 29822 3680 29828 3732
rect 29880 3680 29886 3732
rect 32674 3729 32680 3732
rect 32664 3723 32680 3729
rect 32664 3689 32676 3723
rect 32664 3683 32680 3689
rect 32674 3680 32680 3683
rect 32732 3680 32738 3732
rect 34514 3680 34520 3732
rect 34572 3680 34578 3732
rect 34606 3680 34612 3732
rect 34664 3720 34670 3732
rect 35618 3720 35624 3732
rect 34664 3692 35624 3720
rect 34664 3680 34670 3692
rect 35618 3680 35624 3692
rect 35676 3680 35682 3732
rect 37090 3680 37096 3732
rect 37148 3720 37154 3732
rect 37737 3723 37795 3729
rect 37737 3720 37749 3723
rect 37148 3692 37749 3720
rect 37148 3680 37154 3692
rect 37737 3689 37749 3692
rect 37783 3689 37795 3723
rect 37737 3683 37795 3689
rect 38378 3680 38384 3732
rect 38436 3680 38442 3732
rect 39485 3723 39543 3729
rect 39485 3689 39497 3723
rect 39531 3720 39543 3723
rect 40494 3720 40500 3732
rect 39531 3692 40500 3720
rect 39531 3689 39543 3692
rect 39485 3683 39543 3689
rect 40494 3680 40500 3692
rect 40552 3680 40558 3732
rect 33962 3612 33968 3664
rect 34020 3652 34026 3664
rect 37366 3652 37372 3664
rect 34020 3624 37372 3652
rect 34020 3612 34026 3624
rect 37366 3612 37372 3624
rect 37424 3612 37430 3664
rect 30466 3584 30472 3596
rect 28644 3556 30472 3584
rect 28537 3547 28595 3553
rect 30466 3544 30472 3556
rect 30524 3584 30530 3596
rect 32401 3587 32459 3593
rect 32401 3584 32413 3587
rect 30524 3556 32413 3584
rect 30524 3544 30530 3556
rect 32401 3553 32413 3556
rect 32447 3584 32459 3587
rect 32766 3584 32772 3596
rect 32447 3556 32772 3584
rect 32447 3553 32459 3556
rect 32401 3547 32459 3553
rect 32766 3544 32772 3556
rect 32824 3544 32830 3596
rect 33226 3544 33232 3596
rect 33284 3584 33290 3596
rect 33284 3556 34376 3584
rect 33284 3544 33290 3556
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17644 3488 17693 3516
rect 17644 3476 17650 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18196 3488 18521 3516
rect 18196 3476 18202 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23808 3488 23857 3516
rect 23808 3476 23814 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 25958 3476 25964 3528
rect 26016 3516 26022 3528
rect 26421 3519 26479 3525
rect 26421 3516 26433 3519
rect 26016 3488 26433 3516
rect 26016 3476 26022 3488
rect 26421 3485 26433 3488
rect 26467 3485 26479 3519
rect 28994 3516 29000 3528
rect 26421 3479 26479 3485
rect 28644 3488 29000 3516
rect 24673 3451 24731 3457
rect 24673 3448 24685 3451
rect 15841 3411 15899 3417
rect 24228 3420 24685 3448
rect 9784 3352 12296 3380
rect 12391 3383 12449 3389
rect 12391 3349 12403 3383
rect 12437 3380 12449 3383
rect 12710 3380 12716 3392
rect 12437 3352 12716 3380
rect 12437 3349 12449 3352
rect 12391 3343 12449 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 15856 3380 15884 3411
rect 13955 3352 15884 3380
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 17954 3380 17960 3392
rect 16172 3352 17960 3380
rect 16172 3340 16178 3352
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18138 3340 18144 3392
rect 18196 3340 18202 3392
rect 24228 3389 24256 3420
rect 24673 3417 24685 3420
rect 24719 3417 24731 3451
rect 25898 3420 27278 3448
rect 24673 3411 24731 3417
rect 24213 3383 24271 3389
rect 24213 3349 24225 3383
rect 24259 3349 24271 3383
rect 27172 3380 27200 3420
rect 28644 3380 28672 3488
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 30009 3519 30067 3525
rect 30009 3485 30021 3519
rect 30055 3516 30067 3519
rect 30558 3516 30564 3528
rect 30055 3488 30564 3516
rect 30055 3485 30067 3488
rect 30009 3479 30067 3485
rect 30558 3476 30564 3488
rect 30616 3476 30622 3528
rect 30834 3476 30840 3528
rect 30892 3476 30898 3528
rect 34348 3525 34376 3556
rect 34698 3544 34704 3596
rect 34756 3584 34762 3596
rect 35253 3587 35311 3593
rect 35253 3584 35265 3587
rect 34756 3556 35265 3584
rect 34756 3544 34762 3556
rect 35253 3553 35265 3556
rect 35299 3553 35311 3587
rect 35253 3547 35311 3553
rect 35434 3544 35440 3596
rect 35492 3544 35498 3596
rect 35894 3544 35900 3596
rect 35952 3544 35958 3596
rect 36906 3544 36912 3596
rect 36964 3544 36970 3596
rect 37182 3544 37188 3596
rect 37240 3544 37246 3596
rect 38396 3584 38424 3680
rect 39393 3587 39451 3593
rect 39393 3584 39405 3587
rect 38396 3556 39405 3584
rect 34241 3519 34299 3525
rect 34241 3485 34253 3519
rect 34287 3485 34299 3519
rect 34241 3479 34299 3485
rect 34333 3519 34391 3525
rect 34333 3485 34345 3519
rect 34379 3485 34391 3519
rect 34333 3479 34391 3485
rect 35805 3519 35863 3525
rect 35805 3485 35817 3519
rect 35851 3516 35863 3519
rect 36541 3519 36599 3525
rect 36541 3516 36553 3519
rect 35851 3488 36553 3516
rect 35851 3485 35863 3488
rect 35805 3479 35863 3485
rect 36541 3485 36553 3488
rect 36587 3485 36599 3519
rect 36541 3479 36599 3485
rect 31846 3408 31852 3460
rect 31904 3448 31910 3460
rect 34256 3448 34284 3479
rect 34422 3448 34428 3460
rect 31904 3420 33166 3448
rect 33980 3420 34428 3448
rect 31904 3408 31910 3420
rect 27172 3352 28672 3380
rect 32263 3383 32321 3389
rect 24213 3343 24271 3349
rect 32263 3349 32275 3383
rect 32309 3380 32321 3383
rect 33980 3380 34008 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 34517 3451 34575 3457
rect 34517 3417 34529 3451
rect 34563 3448 34575 3451
rect 34701 3451 34759 3457
rect 34701 3448 34713 3451
rect 34563 3420 34713 3448
rect 34563 3417 34575 3420
rect 34517 3411 34575 3417
rect 34701 3417 34713 3420
rect 34747 3417 34759 3451
rect 36924 3448 36952 3544
rect 37550 3476 37556 3528
rect 37608 3516 37614 3528
rect 38010 3516 38016 3528
rect 37608 3488 38016 3516
rect 37608 3476 37614 3488
rect 38010 3476 38016 3488
rect 38068 3516 38074 3528
rect 38672 3525 38700 3556
rect 39393 3553 39405 3556
rect 39439 3553 39451 3587
rect 39393 3547 39451 3553
rect 39574 3544 39580 3596
rect 39632 3544 39638 3596
rect 38289 3519 38347 3525
rect 38289 3516 38301 3519
rect 38068 3488 38301 3516
rect 38068 3476 38074 3488
rect 38289 3485 38301 3488
rect 38335 3485 38347 3519
rect 38289 3479 38347 3485
rect 38473 3519 38531 3525
rect 38473 3485 38485 3519
rect 38519 3485 38531 3519
rect 38473 3479 38531 3485
rect 38657 3519 38715 3525
rect 38657 3485 38669 3519
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 38488 3448 38516 3479
rect 39298 3476 39304 3528
rect 39356 3476 39362 3528
rect 36924 3420 38516 3448
rect 34701 3411 34759 3417
rect 32309 3352 34008 3380
rect 32309 3349 32321 3352
rect 32263 3343 32321 3349
rect 34146 3340 34152 3392
rect 34204 3380 34210 3392
rect 34606 3380 34612 3392
rect 34204 3352 34612 3380
rect 34204 3340 34210 3352
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 38562 3340 38568 3392
rect 38620 3340 38626 3392
rect 1104 3290 45172 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 45172 3290
rect 1104 3216 45172 3238
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4522 3176 4528 3188
rect 4479 3148 4528 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 6178 3136 6184 3188
rect 6236 3136 6242 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 12894 3176 12900 3188
rect 12851 3148 12900 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 5552 3108 5580 3136
rect 5474 3080 5580 3108
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 6012 3108 6040 3136
rect 5951 3080 6040 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 6196 3049 6224 3136
rect 9490 3108 9496 3120
rect 9062 3080 9496 3108
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 12820 3108 12848 3139
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 13780 3148 14381 3176
rect 13780 3136 13786 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 14369 3139 14427 3145
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 14608 3148 14749 3176
rect 14608 3136 14614 3148
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 14737 3139 14795 3145
rect 16945 3179 17003 3185
rect 16945 3145 16957 3179
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 18138 3176 18144 3188
rect 17359 3148 18144 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 12268 3080 12848 3108
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 7650 3040 7656 3052
rect 6227 3012 7656 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 9582 3000 9588 3052
rect 9640 3000 9646 3052
rect 12158 3000 12164 3052
rect 12216 3000 12222 3052
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7607 2944 8033 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 9447 2907 9505 2913
rect 9447 2873 9459 2907
rect 9493 2904 9505 2907
rect 9600 2904 9628 3000
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 12066 2972 12072 2984
rect 10275 2944 12072 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12268 2981 12296 3080
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 12710 3040 12716 3052
rect 12667 3012 12716 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 16301 3043 16359 3049
rect 13688 3012 15056 3040
rect 13688 3000 13694 3012
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2972 12587 2975
rect 13538 2972 13544 2984
rect 12575 2944 13544 2972
rect 12575 2941 12587 2944
rect 12529 2935 12587 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 14826 2932 14832 2984
rect 14884 2932 14890 2984
rect 15028 2981 15056 3012
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16960 3040 16988 3139
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 25590 3176 25596 3188
rect 22066 3148 25596 3176
rect 17402 3068 17408 3120
rect 17460 3068 17466 3120
rect 16347 3012 16988 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2972 15071 2975
rect 16114 2972 16120 2984
rect 15059 2944 16120 2972
rect 15059 2941 15071 2944
rect 15013 2935 15071 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17586 2932 17592 2984
rect 17644 2932 17650 2984
rect 22066 2972 22094 3148
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 26050 3136 26056 3188
rect 26108 3136 26114 3188
rect 26697 3179 26755 3185
rect 26697 3145 26709 3179
rect 26743 3176 26755 3179
rect 27062 3176 27068 3188
rect 26743 3148 27068 3176
rect 26743 3145 26755 3148
rect 26697 3139 26755 3145
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 27338 3176 27344 3188
rect 27264 3148 27344 3176
rect 27264 3117 27292 3148
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 28813 3179 28871 3185
rect 28813 3145 28825 3179
rect 28859 3176 28871 3179
rect 29362 3176 29368 3188
rect 28859 3148 29368 3176
rect 28859 3145 28871 3148
rect 28813 3139 28871 3145
rect 29362 3136 29368 3148
rect 29420 3136 29426 3188
rect 30466 3136 30472 3188
rect 30524 3136 30530 3188
rect 30558 3136 30564 3188
rect 30616 3176 30622 3188
rect 30653 3179 30711 3185
rect 30653 3176 30665 3179
rect 30616 3148 30665 3176
rect 30616 3136 30622 3148
rect 30653 3145 30665 3148
rect 30699 3145 30711 3179
rect 30653 3139 30711 3145
rect 30834 3136 30840 3188
rect 30892 3176 30898 3188
rect 31389 3179 31447 3185
rect 31389 3176 31401 3179
rect 30892 3148 31401 3176
rect 30892 3136 30898 3148
rect 31389 3145 31401 3148
rect 31435 3145 31447 3179
rect 31389 3139 31447 3145
rect 31726 3148 34560 3176
rect 27249 3111 27307 3117
rect 27249 3077 27261 3111
rect 27295 3077 27307 3111
rect 28994 3108 29000 3120
rect 28474 3080 29000 3108
rect 27249 3071 27307 3077
rect 28994 3068 29000 3080
rect 29052 3068 29058 3120
rect 29730 3068 29736 3120
rect 29788 3068 29794 3120
rect 30484 3108 30512 3136
rect 31726 3108 31754 3148
rect 34532 3120 34560 3148
rect 34698 3136 34704 3188
rect 34756 3176 34762 3188
rect 34993 3179 35051 3185
rect 34993 3176 35005 3179
rect 34756 3148 35005 3176
rect 34756 3136 34762 3148
rect 34993 3145 35005 3148
rect 35039 3145 35051 3179
rect 34993 3139 35051 3145
rect 35434 3136 35440 3188
rect 35492 3176 35498 3188
rect 37093 3179 37151 3185
rect 35492 3148 35664 3176
rect 35492 3136 35498 3148
rect 30484 3080 30604 3108
rect 26510 3000 26516 3052
rect 26568 3040 26574 3052
rect 30576 3049 30604 3080
rect 31128 3080 31754 3108
rect 26973 3043 27031 3049
rect 26973 3040 26985 3043
rect 26568 3012 26985 3040
rect 26568 3000 26574 3012
rect 26973 3009 26985 3012
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 30561 3043 30619 3049
rect 30561 3009 30573 3043
rect 30607 3009 30619 3043
rect 30561 3003 30619 3009
rect 17696 2944 22094 2972
rect 25593 2975 25651 2981
rect 9493 2876 9628 2904
rect 9493 2873 9505 2876
rect 9447 2867 9505 2873
rect 10502 2864 10508 2916
rect 10560 2864 10566 2916
rect 10689 2907 10747 2913
rect 10689 2873 10701 2907
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 10704 2836 10732 2867
rect 12802 2864 12808 2916
rect 12860 2904 12866 2916
rect 14844 2904 14872 2932
rect 12860 2876 14872 2904
rect 16485 2907 16543 2913
rect 12860 2864 12866 2876
rect 16485 2873 16497 2907
rect 16531 2904 16543 2907
rect 17512 2904 17540 2932
rect 16531 2876 17540 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 17696 2836 17724 2944
rect 25593 2941 25605 2975
rect 25639 2972 25651 2975
rect 26237 2975 26295 2981
rect 26237 2972 26249 2975
rect 25639 2944 26249 2972
rect 25639 2941 25651 2944
rect 25593 2935 25651 2941
rect 26237 2941 26249 2944
rect 26283 2972 26295 2975
rect 28721 2975 28779 2981
rect 26283 2944 28672 2972
rect 26283 2941 26295 2944
rect 26237 2935 26295 2941
rect 18046 2864 18052 2916
rect 18104 2904 18110 2916
rect 25608 2904 25636 2935
rect 18104 2876 25636 2904
rect 18104 2864 18110 2876
rect 25866 2864 25872 2916
rect 25924 2864 25930 2916
rect 26602 2864 26608 2916
rect 26660 2864 26666 2916
rect 28644 2904 28672 2944
rect 28721 2941 28733 2975
rect 28767 2972 28779 2975
rect 28994 2972 29000 2984
rect 28767 2944 29000 2972
rect 28767 2941 28779 2944
rect 28721 2935 28779 2941
rect 28994 2932 29000 2944
rect 29052 2932 29058 2984
rect 30282 2932 30288 2984
rect 30340 2932 30346 2984
rect 31128 2981 31156 3080
rect 33778 3068 33784 3120
rect 33836 3068 33842 3120
rect 34514 3068 34520 3120
rect 34572 3068 34578 3120
rect 34606 3068 34612 3120
rect 34664 3108 34670 3120
rect 34793 3111 34851 3117
rect 34793 3108 34805 3111
rect 34664 3080 34805 3108
rect 34664 3068 34670 3080
rect 34793 3077 34805 3080
rect 34839 3077 34851 3111
rect 35526 3108 35532 3120
rect 34793 3071 34851 3077
rect 34900 3080 35532 3108
rect 31481 3043 31539 3049
rect 31481 3009 31493 3043
rect 31527 3040 31539 3043
rect 32769 3043 32827 3049
rect 31527 3012 31754 3040
rect 31527 3009 31539 3012
rect 31481 3003 31539 3009
rect 31113 2975 31171 2981
rect 31113 2972 31125 2975
rect 30484 2944 31125 2972
rect 28644 2876 29316 2904
rect 10704 2808 17724 2836
rect 29288 2836 29316 2876
rect 30484 2836 30512 2944
rect 31113 2941 31125 2944
rect 31159 2941 31171 2975
rect 31113 2935 31171 2941
rect 30834 2864 30840 2916
rect 30892 2864 30898 2916
rect 29288 2808 30512 2836
rect 31726 2836 31754 3012
rect 32769 3009 32781 3043
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 32214 2836 32220 2848
rect 31726 2808 32220 2836
rect 32214 2796 32220 2808
rect 32272 2836 32278 2848
rect 32585 2839 32643 2845
rect 32585 2836 32597 2839
rect 32272 2808 32597 2836
rect 32272 2796 32278 2808
rect 32585 2805 32597 2808
rect 32631 2805 32643 2839
rect 32784 2836 32812 3003
rect 32858 3000 32864 3052
rect 32916 3040 32922 3052
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32916 3012 32965 3040
rect 32916 3000 32922 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 33229 2975 33287 2981
rect 33229 2941 33241 2975
rect 33275 2972 33287 2975
rect 34900 2972 34928 3080
rect 35526 3068 35532 3080
rect 35584 3068 35590 3120
rect 35636 3117 35664 3148
rect 37093 3145 37105 3179
rect 37139 3176 37151 3179
rect 37182 3176 37188 3188
rect 37139 3148 37188 3176
rect 37139 3145 37151 3148
rect 37093 3139 37151 3145
rect 37182 3136 37188 3148
rect 37240 3136 37246 3188
rect 37550 3136 37556 3188
rect 37608 3136 37614 3188
rect 39206 3136 39212 3188
rect 39264 3136 39270 3188
rect 41230 3176 41236 3188
rect 40604 3148 41236 3176
rect 35621 3111 35679 3117
rect 35621 3077 35633 3111
rect 35667 3077 35679 3111
rect 39224 3108 39252 3136
rect 40604 3117 40632 3148
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 42058 3136 42064 3188
rect 42116 3136 42122 3188
rect 40589 3111 40647 3117
rect 39224 3080 39344 3108
rect 35621 3071 35679 3077
rect 35342 3000 35348 3052
rect 35400 3000 35406 3052
rect 36722 3000 36728 3052
rect 36780 3040 36786 3052
rect 39316 3049 39344 3080
rect 40589 3077 40601 3111
rect 40635 3077 40647 3111
rect 42334 3108 42340 3120
rect 41814 3080 42340 3108
rect 40589 3071 40647 3077
rect 42334 3068 42340 3080
rect 42392 3068 42398 3120
rect 39301 3043 39359 3049
rect 36780 3012 37950 3040
rect 36780 3000 36786 3012
rect 39301 3009 39313 3043
rect 39347 3040 39359 3043
rect 40313 3043 40371 3049
rect 40313 3040 40325 3043
rect 39347 3012 40325 3040
rect 39347 3009 39359 3012
rect 39301 3003 39359 3009
rect 40313 3009 40325 3012
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 36740 2972 36768 3000
rect 33275 2944 34928 2972
rect 35452 2944 36768 2972
rect 33275 2941 33287 2944
rect 33229 2935 33287 2941
rect 34238 2864 34244 2916
rect 34296 2904 34302 2916
rect 35452 2904 35480 2944
rect 38562 2932 38568 2984
rect 38620 2972 38626 2984
rect 39025 2975 39083 2981
rect 39025 2972 39037 2975
rect 38620 2944 39037 2972
rect 38620 2932 38626 2944
rect 39025 2941 39037 2944
rect 39071 2941 39083 2975
rect 39025 2935 39083 2941
rect 34296 2876 35480 2904
rect 34296 2864 34302 2876
rect 34422 2836 34428 2848
rect 32784 2808 34428 2836
rect 32585 2799 32643 2805
rect 34422 2796 34428 2808
rect 34480 2836 34486 2848
rect 34977 2839 35035 2845
rect 34977 2836 34989 2839
rect 34480 2808 34989 2836
rect 34480 2796 34486 2808
rect 34977 2805 34989 2808
rect 35023 2805 35035 2839
rect 34977 2799 35035 2805
rect 35161 2839 35219 2845
rect 35161 2805 35173 2839
rect 35207 2836 35219 2839
rect 35710 2836 35716 2848
rect 35207 2808 35716 2836
rect 35207 2805 35219 2808
rect 35161 2799 35219 2805
rect 35710 2796 35716 2808
rect 35768 2796 35774 2848
rect 1104 2746 45172 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 45172 2746
rect 1104 2672 45172 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2632 8815 2635
rect 10502 2632 10508 2644
rect 8803 2604 10508 2632
rect 8803 2601 8815 2604
rect 8757 2595 8815 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 12066 2592 12072 2644
rect 12124 2592 12130 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 25866 2632 25872 2644
rect 17727 2604 25872 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 25866 2592 25872 2604
rect 25924 2592 25930 2644
rect 26602 2592 26608 2644
rect 26660 2632 26666 2644
rect 26697 2635 26755 2641
rect 26697 2632 26709 2635
rect 26660 2604 26709 2632
rect 26660 2592 26666 2604
rect 26697 2601 26709 2604
rect 26743 2601 26755 2635
rect 26697 2595 26755 2601
rect 30193 2635 30251 2641
rect 30193 2601 30205 2635
rect 30239 2632 30251 2635
rect 30282 2632 30288 2644
rect 30239 2604 30288 2632
rect 30239 2601 30251 2604
rect 30193 2595 30251 2601
rect 30282 2592 30288 2604
rect 30340 2592 30346 2644
rect 32674 2592 32680 2644
rect 32732 2592 32738 2644
rect 43898 2592 43904 2644
rect 43956 2592 43962 2644
rect 12084 2564 12112 2592
rect 18046 2564 18052 2576
rect 12084 2536 18052 2564
rect 18046 2524 18052 2536
rect 18104 2524 18110 2576
rect 7190 2456 7196 2508
rect 7248 2456 7254 2508
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8294 2496 8300 2508
rect 8251 2468 8300 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 29178 2456 29184 2508
rect 29236 2496 29242 2508
rect 29549 2499 29607 2505
rect 29549 2496 29561 2499
rect 29236 2468 29561 2496
rect 29236 2456 29242 2468
rect 29549 2465 29561 2468
rect 29595 2465 29607 2499
rect 29549 2459 29607 2465
rect 32214 2456 32220 2508
rect 32272 2456 32278 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7883 2400 8125 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 26510 2388 26516 2440
rect 26568 2388 26574 2440
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2428 32367 2431
rect 33226 2428 33232 2440
rect 32355 2400 33232 2428
rect 32355 2397 32367 2400
rect 32309 2391 32367 2397
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 44085 2431 44143 2437
rect 44085 2428 44097 2431
rect 43864 2400 44097 2428
rect 43864 2388 43870 2400
rect 44085 2397 44097 2400
rect 44131 2397 44143 2431
rect 44085 2391 44143 2397
rect 1104 2202 45172 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 45172 2202
rect 1104 2128 45172 2150
<< via1 >>
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 14832 46112 14884 46164
rect 940 45976 992 46028
rect 1676 45951 1728 45960
rect 1676 45917 1685 45951
rect 1685 45917 1719 45951
rect 1719 45917 1728 45951
rect 1676 45908 1728 45917
rect 6460 45908 6512 45960
rect 9864 45951 9916 45960
rect 9864 45917 9873 45951
rect 9873 45917 9907 45951
rect 9907 45917 9916 45951
rect 9864 45908 9916 45917
rect 14832 45951 14884 45960
rect 14832 45917 14841 45951
rect 14841 45917 14875 45951
rect 14875 45917 14884 45951
rect 14832 45908 14884 45917
rect 21824 46019 21876 46028
rect 21824 45985 21833 46019
rect 21833 45985 21867 46019
rect 21867 45985 21876 46019
rect 21824 45976 21876 45985
rect 24124 45976 24176 46028
rect 22192 45951 22244 45960
rect 22192 45917 22201 45951
rect 22201 45917 22235 45951
rect 22235 45917 22244 45951
rect 22192 45908 22244 45917
rect 23848 45908 23900 45960
rect 15936 45840 15988 45892
rect 27896 45908 27948 45960
rect 33140 45951 33192 45960
rect 33140 45917 33149 45951
rect 33149 45917 33183 45951
rect 33183 45917 33192 45951
rect 33140 45908 33192 45917
rect 41880 45908 41932 45960
rect 7472 45772 7524 45824
rect 8852 45772 8904 45824
rect 14004 45772 14056 45824
rect 24952 45772 25004 45824
rect 27528 45815 27580 45824
rect 27528 45781 27537 45815
rect 27537 45781 27571 45815
rect 27571 45781 27580 45815
rect 27528 45772 27580 45781
rect 41972 45883 42024 45892
rect 41972 45849 41981 45883
rect 41981 45849 42015 45883
rect 42015 45849 42024 45883
rect 41972 45840 42024 45849
rect 29092 45772 29144 45824
rect 32036 45772 32088 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 22192 45568 22244 45620
rect 27896 45611 27948 45620
rect 27896 45577 27923 45611
rect 27923 45577 27948 45611
rect 10048 45500 10100 45552
rect 10140 45432 10192 45484
rect 11704 45475 11756 45484
rect 11704 45441 11713 45475
rect 11713 45441 11747 45475
rect 11747 45441 11756 45475
rect 11704 45432 11756 45441
rect 13728 45500 13780 45552
rect 15936 45500 15988 45552
rect 16304 45500 16356 45552
rect 16488 45500 16540 45552
rect 13544 45475 13596 45484
rect 13544 45441 13578 45475
rect 13578 45441 13596 45475
rect 13544 45432 13596 45441
rect 9956 45407 10008 45416
rect 9956 45373 9965 45407
rect 9965 45373 9999 45407
rect 9999 45373 10008 45407
rect 9956 45364 10008 45373
rect 12532 45364 12584 45416
rect 9036 45271 9088 45280
rect 9036 45237 9045 45271
rect 9045 45237 9079 45271
rect 9079 45237 9088 45271
rect 9036 45228 9088 45237
rect 11520 45271 11572 45280
rect 11520 45237 11529 45271
rect 11529 45237 11563 45271
rect 11563 45237 11572 45271
rect 11520 45228 11572 45237
rect 14740 45271 14792 45280
rect 14740 45237 14749 45271
rect 14749 45237 14783 45271
rect 14783 45237 14792 45271
rect 14740 45228 14792 45237
rect 16580 45296 16632 45348
rect 16856 45432 16908 45484
rect 25872 45500 25924 45552
rect 27896 45568 27948 45577
rect 28080 45543 28132 45552
rect 28080 45509 28089 45543
rect 28089 45509 28123 45543
rect 28123 45509 28132 45543
rect 28080 45500 28132 45509
rect 18420 45475 18472 45484
rect 18420 45441 18429 45475
rect 18429 45441 18463 45475
rect 18463 45441 18472 45475
rect 18420 45432 18472 45441
rect 22008 45475 22060 45484
rect 22008 45441 22017 45475
rect 22017 45441 22051 45475
rect 22051 45441 22060 45475
rect 22008 45432 22060 45441
rect 23388 45432 23440 45484
rect 23940 45432 23992 45484
rect 24124 45432 24176 45484
rect 17316 45364 17368 45416
rect 23480 45407 23532 45416
rect 23480 45373 23489 45407
rect 23489 45373 23523 45407
rect 23523 45373 23532 45407
rect 23480 45364 23532 45373
rect 28540 45432 28592 45484
rect 26700 45364 26752 45416
rect 29644 45407 29696 45416
rect 29644 45373 29653 45407
rect 29653 45373 29687 45407
rect 29687 45373 29696 45407
rect 29644 45364 29696 45373
rect 29920 45407 29972 45416
rect 29920 45373 29929 45407
rect 29929 45373 29963 45407
rect 29963 45373 29972 45407
rect 29920 45364 29972 45373
rect 16212 45271 16264 45280
rect 16212 45237 16221 45271
rect 16221 45237 16255 45271
rect 16255 45237 16264 45271
rect 16212 45228 16264 45237
rect 17040 45228 17092 45280
rect 18236 45271 18288 45280
rect 18236 45237 18245 45271
rect 18245 45237 18279 45271
rect 18279 45237 18288 45271
rect 18236 45228 18288 45237
rect 22376 45228 22428 45280
rect 24032 45271 24084 45280
rect 24032 45237 24041 45271
rect 24041 45237 24075 45271
rect 24075 45237 24084 45271
rect 24032 45228 24084 45237
rect 25136 45228 25188 45280
rect 25504 45271 25556 45280
rect 25504 45237 25513 45271
rect 25513 45237 25547 45271
rect 25547 45237 25556 45271
rect 25504 45228 25556 45237
rect 26424 45228 26476 45280
rect 27160 45228 27212 45280
rect 30012 45271 30064 45280
rect 30012 45237 30021 45271
rect 30021 45237 30055 45271
rect 30055 45237 30064 45271
rect 30012 45228 30064 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 9036 45024 9088 45076
rect 11520 45024 11572 45076
rect 13544 45024 13596 45076
rect 8944 44931 8996 44940
rect 8944 44897 8953 44931
rect 8953 44897 8987 44931
rect 8987 44897 8996 44931
rect 8944 44888 8996 44897
rect 11980 44888 12032 44940
rect 12900 44888 12952 44940
rect 14464 44956 14516 45008
rect 16304 45024 16356 45076
rect 14740 44888 14792 44940
rect 15292 44888 15344 44940
rect 16212 44888 16264 44940
rect 18236 45024 18288 45076
rect 24032 45024 24084 45076
rect 28080 45024 28132 45076
rect 29644 45024 29696 45076
rect 30012 45024 30064 45076
rect 23572 44956 23624 45008
rect 8852 44820 8904 44872
rect 13820 44863 13872 44872
rect 13820 44829 13829 44863
rect 13829 44829 13863 44863
rect 13863 44829 13872 44863
rect 13820 44820 13872 44829
rect 10508 44752 10560 44804
rect 8576 44727 8628 44736
rect 8576 44693 8585 44727
rect 8585 44693 8619 44727
rect 8619 44693 8628 44727
rect 8576 44684 8628 44693
rect 10048 44684 10100 44736
rect 12164 44684 12216 44736
rect 13268 44684 13320 44736
rect 16672 44752 16724 44804
rect 17868 44752 17920 44804
rect 22192 44888 22244 44940
rect 21180 44820 21232 44872
rect 29092 44931 29144 44940
rect 29092 44897 29101 44931
rect 29101 44897 29135 44931
rect 29135 44897 29144 44931
rect 29092 44888 29144 44897
rect 23664 44820 23716 44872
rect 24124 44820 24176 44872
rect 24400 44863 24452 44872
rect 24400 44829 24409 44863
rect 24409 44829 24443 44863
rect 24443 44829 24452 44863
rect 24400 44820 24452 44829
rect 26240 44863 26292 44872
rect 26240 44829 26249 44863
rect 26249 44829 26283 44863
rect 26283 44829 26292 44863
rect 26240 44820 26292 44829
rect 20628 44752 20680 44804
rect 22652 44752 22704 44804
rect 23756 44752 23808 44804
rect 25136 44752 25188 44804
rect 26516 44795 26568 44804
rect 26516 44761 26525 44795
rect 26525 44761 26559 44795
rect 26559 44761 26568 44795
rect 26516 44752 26568 44761
rect 28540 44752 28592 44804
rect 16856 44684 16908 44736
rect 19064 44727 19116 44736
rect 19064 44693 19073 44727
rect 19073 44693 19107 44727
rect 19107 44693 19116 44727
rect 19064 44684 19116 44693
rect 23480 44684 23532 44736
rect 25688 44684 25740 44736
rect 28080 44727 28132 44736
rect 28080 44693 28089 44727
rect 28089 44693 28123 44727
rect 28123 44693 28132 44727
rect 28080 44684 28132 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 8944 44480 8996 44532
rect 9864 44480 9916 44532
rect 9956 44480 10008 44532
rect 10140 44523 10192 44532
rect 10140 44489 10149 44523
rect 10149 44489 10183 44523
rect 10183 44489 10192 44523
rect 10140 44480 10192 44489
rect 8576 44387 8628 44396
rect 8576 44353 8610 44387
rect 8610 44353 8628 44387
rect 8576 44344 8628 44353
rect 10692 44344 10744 44396
rect 11244 44412 11296 44464
rect 11704 44480 11756 44532
rect 12164 44480 12216 44532
rect 12900 44480 12952 44532
rect 14648 44480 14700 44532
rect 14832 44480 14884 44532
rect 17040 44523 17092 44532
rect 17040 44489 17049 44523
rect 17049 44489 17083 44523
rect 17083 44489 17092 44523
rect 17040 44480 17092 44489
rect 17316 44480 17368 44532
rect 22376 44480 22428 44532
rect 23480 44480 23532 44532
rect 23940 44480 23992 44532
rect 24216 44480 24268 44532
rect 26516 44480 26568 44532
rect 26700 44523 26752 44532
rect 26700 44489 26702 44523
rect 26702 44489 26736 44523
rect 26736 44489 26752 44523
rect 26700 44480 26752 44489
rect 9312 44276 9364 44328
rect 10508 44208 10560 44260
rect 12532 44276 12584 44328
rect 13176 44276 13228 44328
rect 15384 44387 15436 44396
rect 15384 44353 15418 44387
rect 15418 44353 15436 44387
rect 15384 44344 15436 44353
rect 22652 44412 22704 44464
rect 16672 44344 16724 44396
rect 17500 44344 17552 44396
rect 18880 44344 18932 44396
rect 13452 44276 13504 44328
rect 14464 44319 14516 44328
rect 14464 44285 14473 44319
rect 14473 44285 14507 44319
rect 14507 44285 14516 44319
rect 14464 44276 14516 44285
rect 8208 44140 8260 44192
rect 12440 44183 12492 44192
rect 12440 44149 12449 44183
rect 12449 44149 12483 44183
rect 12483 44149 12492 44183
rect 12440 44140 12492 44149
rect 13268 44140 13320 44192
rect 13728 44140 13780 44192
rect 17132 44319 17184 44328
rect 17132 44285 17141 44319
rect 17141 44285 17175 44319
rect 17175 44285 17184 44319
rect 17132 44276 17184 44285
rect 17316 44319 17368 44328
rect 17316 44285 17325 44319
rect 17325 44285 17359 44319
rect 17359 44285 17368 44319
rect 17316 44276 17368 44285
rect 14832 44208 14884 44260
rect 16672 44183 16724 44192
rect 16672 44149 16681 44183
rect 16681 44149 16715 44183
rect 16715 44149 16724 44183
rect 16672 44140 16724 44149
rect 18052 44208 18104 44260
rect 19616 44140 19668 44192
rect 25872 44387 25924 44396
rect 25872 44353 25881 44387
rect 25881 44353 25915 44387
rect 25915 44353 25924 44387
rect 25872 44344 25924 44353
rect 21180 44276 21232 44328
rect 25688 44276 25740 44328
rect 25136 44251 25188 44260
rect 25136 44217 25145 44251
rect 25145 44217 25179 44251
rect 25179 44217 25188 44251
rect 25136 44208 25188 44217
rect 26424 44412 26476 44464
rect 28080 44480 28132 44532
rect 26516 44387 26568 44396
rect 26516 44353 26525 44387
rect 26525 44353 26559 44387
rect 26559 44353 26568 44387
rect 26516 44344 26568 44353
rect 27160 44412 27212 44464
rect 27528 44412 27580 44464
rect 28540 44344 28592 44396
rect 45284 44344 45336 44396
rect 26976 44319 27028 44328
rect 26976 44285 26985 44319
rect 26985 44285 27019 44319
rect 27019 44285 27028 44319
rect 26976 44276 27028 44285
rect 44364 44276 44416 44328
rect 23388 44140 23440 44192
rect 25320 44183 25372 44192
rect 25320 44149 25329 44183
rect 25329 44149 25363 44183
rect 25363 44149 25372 44183
rect 25320 44140 25372 44149
rect 26516 44140 26568 44192
rect 27896 44140 27948 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 8208 43936 8260 43988
rect 10692 43936 10744 43988
rect 13820 43936 13872 43988
rect 15384 43936 15436 43988
rect 18420 43936 18472 43988
rect 18880 43936 18932 43988
rect 22192 43979 22244 43988
rect 22192 43945 22201 43979
rect 22201 43945 22235 43979
rect 22235 43945 22244 43979
rect 22192 43936 22244 43945
rect 23664 43979 23716 43988
rect 23664 43945 23673 43979
rect 23673 43945 23707 43979
rect 23707 43945 23716 43979
rect 23664 43936 23716 43945
rect 13176 43800 13228 43852
rect 11980 43775 12032 43784
rect 11980 43741 11989 43775
rect 11989 43741 12023 43775
rect 12023 43741 12032 43775
rect 11980 43732 12032 43741
rect 12440 43732 12492 43784
rect 14740 43732 14792 43784
rect 12532 43664 12584 43716
rect 12900 43664 12952 43716
rect 15292 43800 15344 43852
rect 16488 43800 16540 43852
rect 18880 43843 18932 43852
rect 18880 43809 18889 43843
rect 18889 43809 18923 43843
rect 18923 43809 18932 43843
rect 18880 43800 18932 43809
rect 16672 43732 16724 43784
rect 19616 43775 19668 43784
rect 19616 43741 19625 43775
rect 19625 43741 19659 43775
rect 19659 43741 19668 43775
rect 19616 43732 19668 43741
rect 17316 43664 17368 43716
rect 23572 43800 23624 43852
rect 26240 43800 26292 43852
rect 26976 43800 27028 43852
rect 29920 43800 29972 43852
rect 31852 43800 31904 43852
rect 33048 43800 33100 43852
rect 20444 43664 20496 43716
rect 8024 43596 8076 43648
rect 14464 43596 14516 43648
rect 14556 43639 14608 43648
rect 14556 43605 14565 43639
rect 14565 43605 14599 43639
rect 14599 43605 14608 43639
rect 14556 43596 14608 43605
rect 18420 43596 18472 43648
rect 19064 43596 19116 43648
rect 20076 43596 20128 43648
rect 23480 43732 23532 43784
rect 23756 43664 23808 43716
rect 25320 43732 25372 43784
rect 22652 43596 22704 43648
rect 30840 43664 30892 43716
rect 27712 43639 27764 43648
rect 27712 43605 27721 43639
rect 27721 43605 27755 43639
rect 27755 43605 27764 43639
rect 27712 43596 27764 43605
rect 28540 43596 28592 43648
rect 31944 43596 31996 43648
rect 33968 43596 34020 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 7748 43435 7800 43444
rect 7748 43401 7757 43435
rect 7757 43401 7791 43435
rect 7791 43401 7800 43435
rect 7748 43392 7800 43401
rect 8024 43392 8076 43444
rect 29920 43392 29972 43444
rect 7472 43324 7524 43376
rect 7932 43324 7984 43376
rect 8852 43324 8904 43376
rect 9312 43324 9364 43376
rect 32220 43324 32272 43376
rect 8300 43299 8352 43308
rect 8300 43265 8304 43299
rect 8304 43265 8338 43299
rect 8338 43265 8352 43299
rect 8300 43256 8352 43265
rect 8484 43299 8536 43308
rect 8484 43265 8493 43299
rect 8493 43265 8527 43299
rect 8527 43265 8536 43299
rect 8484 43256 8536 43265
rect 6920 43231 6972 43240
rect 6920 43197 6929 43231
rect 6929 43197 6963 43231
rect 6963 43197 6972 43231
rect 6920 43188 6972 43197
rect 8760 43299 8812 43308
rect 8760 43265 8769 43299
rect 8769 43265 8803 43299
rect 8803 43265 8812 43299
rect 8760 43256 8812 43265
rect 13360 43299 13412 43308
rect 13360 43265 13369 43299
rect 13369 43265 13403 43299
rect 13403 43265 13412 43299
rect 13360 43256 13412 43265
rect 20812 43256 20864 43308
rect 26792 43256 26844 43308
rect 26884 43256 26936 43308
rect 10692 43188 10744 43240
rect 16672 43231 16724 43240
rect 16672 43197 16681 43231
rect 16681 43197 16715 43231
rect 16715 43197 16724 43231
rect 16672 43188 16724 43197
rect 33876 43299 33928 43308
rect 33876 43265 33885 43299
rect 33885 43265 33919 43299
rect 33919 43265 33928 43299
rect 33876 43256 33928 43265
rect 33968 43231 34020 43240
rect 33968 43197 33977 43231
rect 33977 43197 34011 43231
rect 34011 43197 34020 43231
rect 33968 43188 34020 43197
rect 34244 43231 34296 43240
rect 34244 43197 34253 43231
rect 34253 43197 34287 43231
rect 34287 43197 34296 43231
rect 34244 43188 34296 43197
rect 35532 43256 35584 43308
rect 7472 43095 7524 43104
rect 7472 43061 7481 43095
rect 7481 43061 7515 43095
rect 7515 43061 7524 43095
rect 7472 43052 7524 43061
rect 8116 43095 8168 43104
rect 8116 43061 8125 43095
rect 8125 43061 8159 43095
rect 8159 43061 8168 43095
rect 8116 43052 8168 43061
rect 13176 43095 13228 43104
rect 13176 43061 13185 43095
rect 13185 43061 13219 43095
rect 13219 43061 13228 43095
rect 13176 43052 13228 43061
rect 17316 43095 17368 43104
rect 17316 43061 17325 43095
rect 17325 43061 17359 43095
rect 17359 43061 17368 43095
rect 17316 43052 17368 43061
rect 19156 43052 19208 43104
rect 21180 43052 21232 43104
rect 26976 43052 27028 43104
rect 31668 43052 31720 43104
rect 32220 43052 32272 43104
rect 35532 43052 35584 43104
rect 35716 43095 35768 43104
rect 35716 43061 35725 43095
rect 35725 43061 35759 43095
rect 35759 43061 35768 43095
rect 35716 43052 35768 43061
rect 36912 43052 36964 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 7472 42848 7524 42900
rect 14556 42848 14608 42900
rect 16672 42848 16724 42900
rect 17316 42848 17368 42900
rect 25228 42848 25280 42900
rect 28540 42848 28592 42900
rect 3884 42687 3936 42696
rect 3884 42653 3893 42687
rect 3893 42653 3927 42687
rect 3927 42653 3936 42687
rect 3884 42644 3936 42653
rect 4896 42687 4948 42696
rect 4896 42653 4905 42687
rect 4905 42653 4939 42687
rect 4939 42653 4948 42687
rect 4896 42644 4948 42653
rect 5356 42644 5408 42696
rect 8024 42712 8076 42764
rect 8116 42755 8168 42764
rect 8116 42721 8125 42755
rect 8125 42721 8159 42755
rect 8159 42721 8168 42755
rect 8116 42712 8168 42721
rect 8300 42712 8352 42764
rect 11796 42712 11848 42764
rect 14740 42712 14792 42764
rect 7840 42687 7892 42696
rect 7840 42653 7849 42687
rect 7849 42653 7883 42687
rect 7883 42653 7892 42687
rect 7840 42644 7892 42653
rect 8208 42644 8260 42696
rect 10600 42644 10652 42696
rect 12808 42644 12860 42696
rect 9036 42619 9088 42628
rect 9036 42585 9045 42619
rect 9045 42585 9079 42619
rect 9079 42585 9088 42619
rect 9036 42576 9088 42585
rect 11060 42576 11112 42628
rect 4160 42508 4212 42560
rect 4620 42508 4672 42560
rect 5448 42551 5500 42560
rect 5448 42517 5457 42551
rect 5457 42517 5491 42551
rect 5491 42517 5500 42551
rect 5448 42508 5500 42517
rect 6460 42508 6512 42560
rect 7472 42508 7524 42560
rect 9128 42508 9180 42560
rect 11704 42508 11756 42560
rect 13728 42644 13780 42696
rect 14648 42687 14700 42696
rect 14648 42653 14657 42687
rect 14657 42653 14691 42687
rect 14691 42653 14700 42687
rect 14648 42644 14700 42653
rect 13912 42576 13964 42628
rect 15568 42687 15620 42696
rect 15568 42653 15577 42687
rect 15577 42653 15611 42687
rect 15611 42653 15620 42687
rect 15568 42644 15620 42653
rect 18052 42687 18104 42696
rect 18052 42653 18061 42687
rect 18061 42653 18095 42687
rect 18095 42653 18104 42687
rect 18052 42644 18104 42653
rect 15844 42619 15896 42628
rect 13544 42508 13596 42560
rect 14096 42551 14148 42560
rect 14096 42517 14105 42551
rect 14105 42517 14139 42551
rect 14139 42517 14148 42551
rect 14096 42508 14148 42517
rect 14188 42508 14240 42560
rect 15844 42585 15853 42619
rect 15853 42585 15887 42619
rect 15887 42585 15896 42619
rect 15844 42576 15896 42585
rect 15752 42508 15804 42560
rect 16488 42576 16540 42628
rect 17500 42576 17552 42628
rect 22836 42712 22888 42764
rect 24400 42755 24452 42764
rect 24400 42721 24409 42755
rect 24409 42721 24443 42755
rect 24443 42721 24452 42755
rect 24400 42712 24452 42721
rect 26240 42712 26292 42764
rect 26700 42712 26752 42764
rect 31944 42848 31996 42900
rect 18788 42687 18840 42696
rect 18788 42653 18797 42687
rect 18797 42653 18831 42687
rect 18831 42653 18840 42687
rect 18788 42644 18840 42653
rect 19340 42687 19392 42696
rect 19340 42653 19349 42687
rect 19349 42653 19383 42687
rect 19383 42653 19392 42687
rect 19340 42644 19392 42653
rect 21180 42644 21232 42696
rect 22560 42644 22612 42696
rect 24032 42687 24084 42696
rect 24032 42653 24041 42687
rect 24041 42653 24075 42687
rect 24075 42653 24084 42687
rect 24032 42644 24084 42653
rect 17132 42508 17184 42560
rect 17592 42508 17644 42560
rect 18512 42551 18564 42560
rect 18512 42517 18521 42551
rect 18521 42517 18555 42551
rect 18555 42517 18564 42551
rect 18512 42508 18564 42517
rect 18696 42508 18748 42560
rect 19984 42551 20036 42560
rect 19984 42517 19993 42551
rect 19993 42517 20027 42551
rect 20027 42517 20036 42551
rect 19984 42508 20036 42517
rect 21548 42619 21600 42628
rect 21548 42585 21557 42619
rect 21557 42585 21591 42619
rect 21591 42585 21600 42619
rect 21548 42576 21600 42585
rect 23480 42508 23532 42560
rect 23848 42551 23900 42560
rect 23848 42517 23857 42551
rect 23857 42517 23891 42551
rect 23891 42517 23900 42551
rect 23848 42508 23900 42517
rect 25228 42576 25280 42628
rect 25504 42508 25556 42560
rect 27988 42619 28040 42628
rect 27988 42585 27997 42619
rect 27997 42585 28031 42619
rect 28031 42585 28040 42619
rect 27988 42576 28040 42585
rect 26148 42551 26200 42560
rect 26148 42517 26157 42551
rect 26157 42517 26191 42551
rect 26191 42517 26200 42551
rect 26148 42508 26200 42517
rect 26700 42551 26752 42560
rect 26700 42517 26709 42551
rect 26709 42517 26743 42551
rect 26743 42517 26752 42551
rect 26700 42508 26752 42517
rect 30012 42576 30064 42628
rect 31944 42712 31996 42764
rect 31024 42644 31076 42696
rect 31852 42644 31904 42696
rect 33048 42848 33100 42900
rect 32496 42780 32548 42832
rect 32680 42644 32732 42696
rect 30380 42508 30432 42560
rect 30656 42551 30708 42560
rect 30656 42517 30665 42551
rect 30665 42517 30699 42551
rect 30699 42517 30708 42551
rect 30656 42508 30708 42517
rect 30748 42508 30800 42560
rect 31760 42508 31812 42560
rect 32588 42576 32640 42628
rect 32496 42508 32548 42560
rect 33232 42687 33284 42696
rect 33232 42653 33267 42687
rect 33267 42653 33284 42687
rect 33232 42644 33284 42653
rect 35256 42755 35308 42764
rect 35256 42721 35265 42755
rect 35265 42721 35299 42755
rect 35299 42721 35308 42755
rect 35256 42712 35308 42721
rect 35716 42712 35768 42764
rect 33140 42508 33192 42560
rect 33324 42508 33376 42560
rect 34888 42508 34940 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 3884 42304 3936 42356
rect 5448 42304 5500 42356
rect 5356 42236 5408 42288
rect 6460 42304 6512 42356
rect 6920 42304 6972 42356
rect 6368 42211 6420 42220
rect 6368 42177 6377 42211
rect 6377 42177 6411 42211
rect 6411 42177 6420 42211
rect 6368 42168 6420 42177
rect 8484 42304 8536 42356
rect 8852 42347 8904 42356
rect 8852 42313 8861 42347
rect 8861 42313 8895 42347
rect 8895 42313 8904 42347
rect 8852 42304 8904 42313
rect 11060 42304 11112 42356
rect 11244 42304 11296 42356
rect 11888 42304 11940 42356
rect 13912 42304 13964 42356
rect 14096 42304 14148 42356
rect 15568 42347 15620 42356
rect 15568 42313 15577 42347
rect 15577 42313 15611 42347
rect 15611 42313 15620 42347
rect 15568 42304 15620 42313
rect 17132 42304 17184 42356
rect 19800 42304 19852 42356
rect 6736 42211 6788 42220
rect 6736 42177 6745 42211
rect 6745 42177 6779 42211
rect 6779 42177 6788 42211
rect 6736 42168 6788 42177
rect 3332 42100 3384 42152
rect 5356 42100 5408 42152
rect 6092 42143 6144 42152
rect 6092 42109 6101 42143
rect 6101 42109 6135 42143
rect 6135 42109 6144 42143
rect 6092 42100 6144 42109
rect 4712 42032 4764 42084
rect 5356 41964 5408 42016
rect 5448 41964 5500 42016
rect 7472 42211 7524 42220
rect 7472 42177 7481 42211
rect 7481 42177 7515 42211
rect 7515 42177 7524 42211
rect 7472 42168 7524 42177
rect 8300 42168 8352 42220
rect 8484 42168 8536 42220
rect 9128 42236 9180 42288
rect 10600 42236 10652 42288
rect 10784 42236 10836 42288
rect 11060 42168 11112 42220
rect 11980 42168 12032 42220
rect 13176 42236 13228 42288
rect 14464 42236 14516 42288
rect 13544 42168 13596 42220
rect 11520 42143 11572 42152
rect 11520 42109 11529 42143
rect 11529 42109 11563 42143
rect 11563 42109 11572 42143
rect 11520 42100 11572 42109
rect 13728 42143 13780 42152
rect 13728 42109 13737 42143
rect 13737 42109 13771 42143
rect 13771 42109 13780 42143
rect 13728 42100 13780 42109
rect 17592 42168 17644 42220
rect 18052 42236 18104 42288
rect 21548 42304 21600 42356
rect 23848 42304 23900 42356
rect 24032 42304 24084 42356
rect 26700 42304 26752 42356
rect 18696 42168 18748 42220
rect 8392 41964 8444 42016
rect 10692 42007 10744 42016
rect 10692 41973 10701 42007
rect 10701 41973 10735 42007
rect 10735 41973 10744 42007
rect 10692 41964 10744 41973
rect 11152 42007 11204 42016
rect 11152 41973 11161 42007
rect 11161 41973 11195 42007
rect 11195 41973 11204 42007
rect 11152 41964 11204 41973
rect 12256 41964 12308 42016
rect 14188 41964 14240 42016
rect 15292 41964 15344 42016
rect 17316 42143 17368 42152
rect 17316 42109 17325 42143
rect 17325 42109 17359 42143
rect 17359 42109 17368 42143
rect 17316 42100 17368 42109
rect 19156 42143 19208 42152
rect 19156 42109 19165 42143
rect 19165 42109 19199 42143
rect 19199 42109 19208 42143
rect 19156 42100 19208 42109
rect 19984 42100 20036 42152
rect 20628 42100 20680 42152
rect 15844 42032 15896 42084
rect 22284 42168 22336 42220
rect 23572 42236 23624 42288
rect 22652 42211 22704 42220
rect 22652 42177 22661 42211
rect 22661 42177 22695 42211
rect 22695 42177 22704 42211
rect 22652 42168 22704 42177
rect 22836 42211 22888 42220
rect 22836 42177 22845 42211
rect 22845 42177 22879 42211
rect 22879 42177 22888 42211
rect 22836 42168 22888 42177
rect 23112 42168 23164 42220
rect 22928 42100 22980 42152
rect 26332 42236 26384 42288
rect 26884 42236 26936 42288
rect 25044 42211 25096 42220
rect 25044 42177 25053 42211
rect 25053 42177 25087 42211
rect 25087 42177 25096 42211
rect 25044 42168 25096 42177
rect 26148 42168 26200 42220
rect 23296 42100 23348 42152
rect 26700 42168 26752 42220
rect 28540 42236 28592 42288
rect 30380 42236 30432 42288
rect 31484 42304 31536 42356
rect 31668 42304 31720 42356
rect 31760 42347 31812 42356
rect 31760 42313 31769 42347
rect 31769 42313 31803 42347
rect 31803 42313 31812 42347
rect 31760 42304 31812 42313
rect 32588 42304 32640 42356
rect 30564 42236 30616 42288
rect 33232 42236 33284 42288
rect 33784 42304 33836 42356
rect 34244 42304 34296 42356
rect 34888 42347 34940 42356
rect 34888 42313 34897 42347
rect 34897 42313 34931 42347
rect 34931 42313 34940 42347
rect 34888 42304 34940 42313
rect 33692 42279 33744 42288
rect 33692 42245 33701 42279
rect 33701 42245 33735 42279
rect 33735 42245 33744 42279
rect 33692 42236 33744 42245
rect 26792 42032 26844 42084
rect 18972 41964 19024 42016
rect 20536 41964 20588 42016
rect 22192 42007 22244 42016
rect 22192 41973 22201 42007
rect 22201 41973 22235 42007
rect 22235 41973 22244 42007
rect 22192 41964 22244 41973
rect 22284 41964 22336 42016
rect 22836 41964 22888 42016
rect 26700 42007 26752 42016
rect 26700 41973 26709 42007
rect 26709 41973 26743 42007
rect 26743 41973 26752 42007
rect 26700 41964 26752 41973
rect 30656 42168 30708 42220
rect 27252 42143 27304 42152
rect 27252 42109 27261 42143
rect 27261 42109 27295 42143
rect 27295 42109 27304 42143
rect 27252 42100 27304 42109
rect 29092 42143 29144 42152
rect 29092 42109 29101 42143
rect 29101 42109 29135 42143
rect 29135 42109 29144 42143
rect 29092 42100 29144 42109
rect 31852 42211 31904 42220
rect 31852 42177 31861 42211
rect 31861 42177 31895 42211
rect 31895 42177 31904 42211
rect 31852 42168 31904 42177
rect 31668 42100 31720 42152
rect 30196 42032 30248 42084
rect 30472 42032 30524 42084
rect 33324 42211 33376 42220
rect 33324 42177 33333 42211
rect 33333 42177 33367 42211
rect 33367 42177 33376 42211
rect 33324 42168 33376 42177
rect 34152 42236 34204 42288
rect 34704 42279 34756 42288
rect 34704 42245 34713 42279
rect 34713 42245 34747 42279
rect 34747 42245 34756 42279
rect 34704 42236 34756 42245
rect 34796 42236 34848 42288
rect 28356 41964 28408 42016
rect 30656 42007 30708 42016
rect 30656 41973 30665 42007
rect 30665 41973 30699 42007
rect 30699 41973 30708 42007
rect 30656 41964 30708 41973
rect 31208 41964 31260 42016
rect 35256 42168 35308 42220
rect 31760 41964 31812 42016
rect 32772 41964 32824 42016
rect 33508 41964 33560 42016
rect 34704 42032 34756 42084
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 3884 41760 3936 41812
rect 4620 41760 4672 41812
rect 4896 41760 4948 41812
rect 5356 41760 5408 41812
rect 6368 41760 6420 41812
rect 8300 41803 8352 41812
rect 8300 41769 8309 41803
rect 8309 41769 8343 41803
rect 8343 41769 8352 41803
rect 8300 41760 8352 41769
rect 8760 41760 8812 41812
rect 2780 41624 2832 41676
rect 3332 41624 3384 41676
rect 4344 41692 4396 41744
rect 1860 41599 1912 41608
rect 1860 41565 1869 41599
rect 1869 41565 1903 41599
rect 1903 41565 1912 41599
rect 1860 41556 1912 41565
rect 4804 41692 4856 41744
rect 5448 41624 5500 41676
rect 4252 41488 4304 41540
rect 4160 41463 4212 41472
rect 4160 41429 4169 41463
rect 4169 41429 4203 41463
rect 4203 41429 4212 41463
rect 4160 41420 4212 41429
rect 4988 41556 5040 41608
rect 5540 41556 5592 41608
rect 6460 41624 6512 41676
rect 10784 41760 10836 41812
rect 11152 41760 11204 41812
rect 11520 41803 11572 41812
rect 11520 41769 11529 41803
rect 11529 41769 11563 41803
rect 11563 41769 11572 41803
rect 11520 41760 11572 41769
rect 11704 41760 11756 41812
rect 12808 41760 12860 41812
rect 13360 41760 13412 41812
rect 17316 41803 17368 41812
rect 17316 41769 17325 41803
rect 17325 41769 17359 41803
rect 17359 41769 17368 41803
rect 17316 41760 17368 41769
rect 18512 41760 18564 41812
rect 18788 41760 18840 41812
rect 19340 41760 19392 41812
rect 5264 41488 5316 41540
rect 9128 41488 9180 41540
rect 11796 41692 11848 41744
rect 11888 41624 11940 41676
rect 13636 41667 13688 41676
rect 13636 41633 13645 41667
rect 13645 41633 13679 41667
rect 13679 41633 13688 41667
rect 13636 41624 13688 41633
rect 19800 41692 19852 41744
rect 14280 41624 14332 41676
rect 12256 41556 12308 41608
rect 14556 41556 14608 41608
rect 18328 41624 18380 41676
rect 9312 41463 9364 41472
rect 9312 41429 9321 41463
rect 9321 41429 9355 41463
rect 9355 41429 9364 41463
rect 9312 41420 9364 41429
rect 9404 41463 9456 41472
rect 9404 41429 9413 41463
rect 9413 41429 9447 41463
rect 9447 41429 9456 41463
rect 9404 41420 9456 41429
rect 10508 41488 10560 41540
rect 11060 41488 11112 41540
rect 15476 41488 15528 41540
rect 11244 41420 11296 41472
rect 13360 41420 13412 41472
rect 13728 41420 13780 41472
rect 15384 41463 15436 41472
rect 15384 41429 15393 41463
rect 15393 41429 15427 41463
rect 15427 41429 15436 41463
rect 16488 41556 16540 41608
rect 18788 41556 18840 41608
rect 16028 41488 16080 41540
rect 20076 41760 20128 41812
rect 20536 41760 20588 41812
rect 23296 41760 23348 41812
rect 26700 41760 26752 41812
rect 27252 41760 27304 41812
rect 29092 41760 29144 41812
rect 29828 41760 29880 41812
rect 30380 41760 30432 41812
rect 30472 41760 30524 41812
rect 30656 41760 30708 41812
rect 30840 41760 30892 41812
rect 20720 41556 20772 41608
rect 21180 41599 21232 41608
rect 21180 41565 21189 41599
rect 21189 41565 21223 41599
rect 21223 41565 21232 41599
rect 21180 41556 21232 41565
rect 23388 41624 23440 41676
rect 23940 41624 23992 41676
rect 31852 41760 31904 41812
rect 23112 41556 23164 41608
rect 23204 41556 23256 41608
rect 23480 41556 23532 41608
rect 26976 41599 27028 41608
rect 26976 41565 26985 41599
rect 26985 41565 27019 41599
rect 27019 41565 27028 41599
rect 26976 41556 27028 41565
rect 28356 41667 28408 41676
rect 28356 41633 28365 41667
rect 28365 41633 28399 41667
rect 28399 41633 28408 41667
rect 28356 41624 28408 41633
rect 30104 41624 30156 41676
rect 30288 41556 30340 41608
rect 30932 41624 30984 41676
rect 30748 41599 30800 41608
rect 30748 41565 30757 41599
rect 30757 41565 30791 41599
rect 30791 41565 30800 41599
rect 30748 41556 30800 41565
rect 31668 41624 31720 41676
rect 31944 41624 31996 41676
rect 32772 41667 32824 41676
rect 15384 41420 15436 41429
rect 17960 41420 18012 41472
rect 18972 41420 19024 41472
rect 21456 41531 21508 41540
rect 21456 41497 21465 41531
rect 21465 41497 21499 41531
rect 21499 41497 21508 41531
rect 21456 41488 21508 41497
rect 22744 41488 22796 41540
rect 22928 41488 22980 41540
rect 25044 41420 25096 41472
rect 26148 41420 26200 41472
rect 27252 41488 27304 41540
rect 29644 41420 29696 41472
rect 29828 41531 29880 41540
rect 29828 41497 29848 41531
rect 29848 41497 29880 41531
rect 29828 41488 29880 41497
rect 30472 41488 30524 41540
rect 30656 41531 30708 41540
rect 30656 41497 30665 41531
rect 30665 41497 30699 41531
rect 30699 41497 30708 41531
rect 30656 41488 30708 41497
rect 31208 41556 31260 41608
rect 31576 41599 31628 41608
rect 31576 41565 31585 41599
rect 31585 41565 31619 41599
rect 31619 41565 31628 41599
rect 31576 41556 31628 41565
rect 32772 41633 32781 41667
rect 32781 41633 32815 41667
rect 32815 41633 32824 41667
rect 32772 41624 32824 41633
rect 33140 41760 33192 41812
rect 33784 41760 33836 41812
rect 33048 41692 33100 41744
rect 34704 41692 34756 41744
rect 31392 41488 31444 41540
rect 32496 41599 32548 41608
rect 32496 41565 32505 41599
rect 32505 41565 32539 41599
rect 32539 41565 32548 41599
rect 32496 41556 32548 41565
rect 32680 41599 32732 41608
rect 32680 41565 32689 41599
rect 32689 41565 32723 41599
rect 32723 41565 32732 41599
rect 32680 41556 32732 41565
rect 33508 41556 33560 41608
rect 33784 41556 33836 41608
rect 34060 41599 34112 41608
rect 34060 41565 34069 41599
rect 34069 41565 34103 41599
rect 34103 41565 34112 41599
rect 34060 41556 34112 41565
rect 34152 41599 34204 41608
rect 34152 41565 34161 41599
rect 34161 41565 34195 41599
rect 34195 41565 34204 41599
rect 34152 41556 34204 41565
rect 34796 41624 34848 41676
rect 30380 41420 30432 41472
rect 33416 41531 33468 41540
rect 33416 41497 33425 41531
rect 33425 41497 33459 41531
rect 33459 41497 33468 41531
rect 33416 41488 33468 41497
rect 33600 41531 33652 41540
rect 33600 41497 33609 41531
rect 33609 41497 33643 41531
rect 33643 41497 33652 41531
rect 33600 41488 33652 41497
rect 31852 41420 31904 41472
rect 31944 41463 31996 41472
rect 31944 41429 31953 41463
rect 31953 41429 31987 41463
rect 31987 41429 31996 41463
rect 31944 41420 31996 41429
rect 34336 41488 34388 41540
rect 34704 41599 34756 41608
rect 34704 41565 34713 41599
rect 34713 41565 34747 41599
rect 34747 41565 34756 41599
rect 34704 41556 34756 41565
rect 35532 41531 35584 41540
rect 35532 41497 35557 41531
rect 35557 41497 35584 41531
rect 35532 41488 35584 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 2780 41216 2832 41268
rect 4160 41216 4212 41268
rect 4528 41216 4580 41268
rect 4988 41216 5040 41268
rect 9312 41216 9364 41268
rect 10508 41259 10560 41268
rect 10508 41225 10517 41259
rect 10517 41225 10551 41259
rect 10551 41225 10560 41259
rect 10508 41216 10560 41225
rect 11888 41259 11940 41268
rect 11888 41225 11897 41259
rect 11897 41225 11931 41259
rect 11931 41225 11940 41259
rect 11888 41216 11940 41225
rect 14188 41216 14240 41268
rect 5172 41148 5224 41200
rect 8024 41148 8076 41200
rect 10416 41148 10468 41200
rect 11244 41148 11296 41200
rect 3792 41012 3844 41064
rect 4160 41123 4212 41132
rect 4160 41089 4169 41123
rect 4169 41089 4203 41123
rect 4203 41089 4212 41123
rect 4160 41080 4212 41089
rect 4344 41123 4396 41132
rect 4344 41089 4352 41123
rect 4352 41089 4386 41123
rect 4386 41089 4396 41123
rect 4344 41080 4396 41089
rect 4528 41123 4580 41132
rect 4528 41089 4537 41123
rect 4537 41089 4571 41123
rect 4571 41089 4580 41123
rect 4528 41080 4580 41089
rect 4712 41123 4764 41132
rect 4712 41089 4719 41123
rect 4719 41089 4764 41123
rect 4712 41080 4764 41089
rect 4804 41123 4856 41132
rect 4804 41089 4813 41123
rect 4813 41089 4847 41123
rect 4847 41089 4856 41123
rect 4804 41080 4856 41089
rect 4988 41123 5040 41132
rect 4988 41089 5002 41123
rect 5002 41089 5036 41123
rect 5036 41089 5040 41123
rect 4988 41080 5040 41089
rect 8852 41080 8904 41132
rect 6092 41012 6144 41064
rect 8116 41055 8168 41064
rect 8116 41021 8125 41055
rect 8125 41021 8159 41055
rect 8159 41021 8168 41055
rect 8116 41012 8168 41021
rect 14280 41123 14332 41132
rect 11980 41055 12032 41064
rect 11980 41021 11989 41055
rect 11989 41021 12023 41055
rect 12023 41021 12032 41055
rect 11980 41012 12032 41021
rect 12164 41055 12216 41064
rect 12164 41021 12173 41055
rect 12173 41021 12207 41055
rect 12207 41021 12216 41055
rect 12164 41012 12216 41021
rect 14280 41089 14284 41123
rect 14284 41089 14318 41123
rect 14318 41089 14332 41123
rect 14280 41080 14332 41089
rect 14556 41080 14608 41132
rect 15292 41148 15344 41200
rect 15752 41259 15804 41268
rect 15752 41225 15761 41259
rect 15761 41225 15795 41259
rect 15795 41225 15804 41259
rect 15752 41216 15804 41225
rect 16028 41216 16080 41268
rect 18788 41259 18840 41268
rect 18788 41225 18797 41259
rect 18797 41225 18831 41259
rect 18831 41225 18840 41259
rect 18788 41216 18840 41225
rect 21180 41216 21232 41268
rect 21456 41216 21508 41268
rect 23480 41216 23532 41268
rect 17316 41148 17368 41200
rect 18328 41148 18380 41200
rect 14740 41123 14792 41132
rect 14740 41089 14749 41123
rect 14749 41089 14783 41123
rect 14783 41089 14792 41123
rect 14740 41080 14792 41089
rect 14648 40944 14700 40996
rect 15844 41055 15896 41064
rect 15844 41021 15853 41055
rect 15853 41021 15887 41055
rect 15887 41021 15896 41055
rect 15844 41012 15896 41021
rect 18696 41123 18748 41132
rect 18696 41089 18705 41123
rect 18705 41089 18739 41123
rect 18739 41089 18748 41123
rect 18696 41080 18748 41089
rect 20444 41148 20496 41200
rect 22192 41148 22244 41200
rect 3516 40876 3568 40928
rect 4252 40876 4304 40928
rect 5448 40876 5500 40928
rect 7472 40919 7524 40928
rect 7472 40885 7481 40919
rect 7481 40885 7515 40919
rect 7515 40885 7524 40919
rect 7472 40876 7524 40885
rect 13636 40876 13688 40928
rect 22560 41012 22612 41064
rect 22836 41123 22888 41132
rect 22836 41089 22845 41123
rect 22845 41089 22879 41123
rect 22879 41089 22888 41123
rect 22836 41080 22888 41089
rect 23296 41148 23348 41200
rect 25320 41216 25372 41268
rect 28264 41216 28316 41268
rect 30288 41216 30340 41268
rect 25228 41148 25280 41200
rect 26792 41148 26844 41200
rect 23204 41123 23256 41132
rect 23204 41089 23213 41123
rect 23213 41089 23247 41123
rect 23247 41089 23256 41123
rect 23204 41080 23256 41089
rect 23480 41080 23532 41132
rect 23664 41012 23716 41064
rect 26332 41080 26384 41132
rect 27252 41080 27304 41132
rect 24400 41055 24452 41064
rect 24400 41021 24409 41055
rect 24409 41021 24443 41055
rect 24443 41021 24452 41055
rect 24400 41012 24452 41021
rect 24676 41055 24728 41064
rect 24676 41021 24685 41055
rect 24685 41021 24719 41055
rect 24719 41021 24728 41055
rect 24676 41012 24728 41021
rect 28816 41191 28868 41200
rect 28816 41157 28825 41191
rect 28825 41157 28859 41191
rect 28859 41157 28868 41191
rect 28816 41148 28868 41157
rect 30840 41216 30892 41268
rect 31668 41216 31720 41268
rect 30932 41191 30984 41200
rect 30932 41157 30941 41191
rect 30941 41157 30975 41191
rect 30975 41157 30984 41191
rect 30932 41148 30984 41157
rect 31576 41148 31628 41200
rect 30564 41012 30616 41064
rect 31208 41080 31260 41132
rect 31852 41080 31904 41132
rect 32128 41123 32180 41132
rect 32128 41089 32137 41123
rect 32137 41089 32171 41123
rect 32171 41089 32180 41123
rect 32128 41080 32180 41089
rect 33692 41216 33744 41268
rect 34244 41216 34296 41268
rect 34796 41216 34848 41268
rect 35072 41216 35124 41268
rect 35532 41216 35584 41268
rect 32496 41148 32548 41200
rect 32404 41123 32456 41132
rect 32404 41089 32413 41123
rect 32413 41089 32447 41123
rect 32447 41089 32456 41123
rect 32404 41080 32456 41089
rect 33048 41148 33100 41200
rect 33600 41080 33652 41132
rect 30932 41012 30984 41064
rect 31116 41055 31168 41064
rect 31116 41021 31125 41055
rect 31125 41021 31159 41055
rect 31159 41021 31168 41055
rect 31116 41012 31168 41021
rect 31576 41055 31628 41064
rect 31576 41021 31585 41055
rect 31585 41021 31619 41055
rect 31619 41021 31628 41055
rect 31576 41012 31628 41021
rect 31944 41012 31996 41064
rect 20536 40876 20588 40928
rect 22652 40919 22704 40928
rect 22652 40885 22661 40919
rect 22661 40885 22695 40919
rect 22695 40885 22704 40919
rect 22652 40876 22704 40885
rect 24492 40876 24544 40928
rect 26516 40876 26568 40928
rect 27160 40876 27212 40928
rect 28264 40919 28316 40928
rect 28264 40885 28273 40919
rect 28273 40885 28307 40919
rect 28307 40885 28316 40919
rect 28264 40876 28316 40885
rect 28356 40876 28408 40928
rect 28540 40876 28592 40928
rect 30288 40919 30340 40928
rect 30288 40885 30297 40919
rect 30297 40885 30331 40919
rect 30331 40885 30340 40919
rect 30288 40876 30340 40885
rect 31208 40919 31260 40928
rect 31208 40885 31217 40919
rect 31217 40885 31251 40919
rect 31251 40885 31260 40919
rect 31208 40876 31260 40885
rect 31760 40944 31812 40996
rect 31392 40876 31444 40928
rect 33784 41080 33836 41132
rect 34704 41148 34756 41200
rect 34336 41123 34388 41132
rect 34336 41089 34345 41123
rect 34345 41089 34379 41123
rect 34379 41089 34388 41123
rect 34336 41080 34388 41089
rect 34520 41080 34572 41132
rect 34428 40876 34480 40928
rect 35808 40876 35860 40928
rect 35900 40876 35952 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 4620 40672 4672 40724
rect 6736 40672 6788 40724
rect 8760 40672 8812 40724
rect 11796 40672 11848 40724
rect 16120 40672 16172 40724
rect 17868 40672 17920 40724
rect 18696 40672 18748 40724
rect 22652 40672 22704 40724
rect 24676 40672 24728 40724
rect 1860 40536 1912 40588
rect 3608 40536 3660 40588
rect 4160 40536 4212 40588
rect 4804 40536 4856 40588
rect 6184 40536 6236 40588
rect 7472 40536 7524 40588
rect 8668 40579 8720 40588
rect 8668 40545 8677 40579
rect 8677 40545 8711 40579
rect 8711 40545 8720 40579
rect 8668 40536 8720 40545
rect 25320 40604 25372 40656
rect 28540 40672 28592 40724
rect 31300 40672 31352 40724
rect 31944 40672 31996 40724
rect 4620 40511 4672 40520
rect 4620 40477 4629 40511
rect 4629 40477 4663 40511
rect 4663 40477 4672 40511
rect 4620 40468 4672 40477
rect 5080 40468 5132 40520
rect 8024 40468 8076 40520
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 3332 40400 3384 40452
rect 4344 40400 4396 40452
rect 8576 40468 8628 40520
rect 11152 40511 11204 40520
rect 11152 40477 11161 40511
rect 11161 40477 11195 40511
rect 11195 40477 11204 40511
rect 11152 40468 11204 40477
rect 15936 40536 15988 40588
rect 10048 40400 10100 40452
rect 11796 40443 11848 40452
rect 11796 40409 11805 40443
rect 11805 40409 11839 40443
rect 11839 40409 11848 40443
rect 11796 40400 11848 40409
rect 11888 40443 11940 40452
rect 11888 40409 11897 40443
rect 11897 40409 11931 40443
rect 11931 40409 11940 40443
rect 11888 40400 11940 40409
rect 13728 40511 13780 40520
rect 13728 40477 13737 40511
rect 13737 40477 13771 40511
rect 13771 40477 13780 40511
rect 13728 40468 13780 40477
rect 14464 40468 14516 40520
rect 17500 40536 17552 40588
rect 19156 40536 19208 40588
rect 4068 40375 4120 40384
rect 4068 40341 4077 40375
rect 4077 40341 4111 40375
rect 4111 40341 4120 40375
rect 4068 40332 4120 40341
rect 8208 40332 8260 40384
rect 8300 40375 8352 40384
rect 8300 40341 8309 40375
rect 8309 40341 8343 40375
rect 8343 40341 8352 40375
rect 8300 40332 8352 40341
rect 8392 40332 8444 40384
rect 9220 40332 9272 40384
rect 12256 40375 12308 40384
rect 12256 40341 12265 40375
rect 12265 40341 12299 40375
rect 12299 40341 12308 40375
rect 12256 40332 12308 40341
rect 13912 40375 13964 40384
rect 13912 40341 13921 40375
rect 13921 40341 13955 40375
rect 13955 40341 13964 40375
rect 13912 40332 13964 40341
rect 16028 40332 16080 40384
rect 17684 40332 17736 40384
rect 20168 40511 20220 40520
rect 20168 40477 20177 40511
rect 20177 40477 20211 40511
rect 20211 40477 20220 40511
rect 20168 40468 20220 40477
rect 23664 40468 23716 40520
rect 20904 40332 20956 40384
rect 24124 40332 24176 40384
rect 26148 40511 26200 40520
rect 26148 40477 26157 40511
rect 26157 40477 26191 40511
rect 26191 40477 26200 40511
rect 26148 40468 26200 40477
rect 26884 40604 26936 40656
rect 26516 40579 26568 40588
rect 26516 40545 26525 40579
rect 26525 40545 26559 40579
rect 26559 40545 26568 40579
rect 26516 40536 26568 40545
rect 27804 40536 27856 40588
rect 31576 40536 31628 40588
rect 32404 40536 32456 40588
rect 27344 40468 27396 40520
rect 28264 40468 28316 40520
rect 35256 40511 35308 40520
rect 35256 40477 35265 40511
rect 35265 40477 35299 40511
rect 35299 40477 35308 40511
rect 35256 40468 35308 40477
rect 26332 40443 26384 40452
rect 26332 40409 26367 40443
rect 26367 40409 26384 40443
rect 26332 40400 26384 40409
rect 30748 40400 30800 40452
rect 35992 40468 36044 40520
rect 38016 40468 38068 40520
rect 26792 40332 26844 40384
rect 26884 40332 26936 40384
rect 27436 40375 27488 40384
rect 27436 40341 27445 40375
rect 27445 40341 27479 40375
rect 27479 40341 27488 40375
rect 27436 40332 27488 40341
rect 35532 40443 35584 40452
rect 35532 40409 35541 40443
rect 35541 40409 35575 40443
rect 35575 40409 35584 40443
rect 35532 40400 35584 40409
rect 35808 40400 35860 40452
rect 36912 40400 36964 40452
rect 35900 40375 35952 40384
rect 35900 40341 35909 40375
rect 35909 40341 35943 40375
rect 35943 40341 35952 40375
rect 35900 40332 35952 40341
rect 37188 40332 37240 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 1860 40128 1912 40180
rect 4068 40128 4120 40180
rect 8116 40128 8168 40180
rect 8576 40128 8628 40180
rect 8668 40128 8720 40180
rect 4344 40060 4396 40112
rect 8024 40060 8076 40112
rect 3608 40035 3660 40044
rect 3608 40001 3617 40035
rect 3617 40001 3651 40035
rect 3651 40001 3660 40035
rect 3608 39992 3660 40001
rect 6184 39992 6236 40044
rect 3516 39967 3568 39976
rect 3516 39933 3525 39967
rect 3525 39933 3559 39967
rect 3559 39933 3568 39967
rect 3516 39924 3568 39933
rect 3976 39924 4028 39976
rect 6644 39967 6696 39976
rect 6644 39933 6653 39967
rect 6653 39933 6687 39967
rect 6687 39933 6696 39967
rect 6644 39924 6696 39933
rect 8484 40035 8536 40044
rect 8484 40001 8493 40035
rect 8493 40001 8527 40035
rect 8527 40001 8536 40035
rect 8484 39992 8536 40001
rect 8576 40035 8628 40044
rect 8576 40001 8585 40035
rect 8585 40001 8619 40035
rect 8619 40001 8628 40035
rect 8576 39992 8628 40001
rect 9772 40128 9824 40180
rect 10416 40128 10468 40180
rect 11888 40128 11940 40180
rect 13728 40128 13780 40180
rect 12256 40060 12308 40112
rect 14648 40128 14700 40180
rect 17684 40128 17736 40180
rect 14464 40060 14516 40112
rect 16948 40060 17000 40112
rect 21180 40128 21232 40180
rect 22744 40128 22796 40180
rect 26240 40128 26292 40180
rect 27436 40128 27488 40180
rect 28172 40128 28224 40180
rect 28264 40128 28316 40180
rect 35256 40171 35308 40180
rect 35256 40137 35265 40171
rect 35265 40137 35299 40171
rect 35299 40137 35308 40171
rect 35256 40128 35308 40137
rect 35532 40128 35584 40180
rect 20628 40060 20680 40112
rect 11152 39992 11204 40044
rect 9220 39924 9272 39976
rect 10048 39924 10100 39976
rect 11060 39967 11112 39976
rect 11060 39933 11069 39967
rect 11069 39933 11103 39967
rect 11103 39933 11112 39967
rect 11060 39924 11112 39933
rect 6092 39831 6144 39840
rect 6092 39797 6101 39831
rect 6101 39797 6135 39831
rect 6135 39797 6144 39831
rect 6092 39788 6144 39797
rect 8116 39788 8168 39840
rect 10784 39788 10836 39840
rect 12440 39924 12492 39976
rect 12808 39967 12860 39976
rect 12808 39933 12817 39967
rect 12817 39933 12851 39967
rect 12851 39933 12860 39967
rect 12808 39924 12860 39933
rect 12992 39967 13044 39976
rect 12992 39933 13001 39967
rect 13001 39933 13035 39967
rect 13035 39933 13044 39967
rect 12992 39924 13044 39933
rect 13912 39924 13964 39976
rect 13544 39788 13596 39840
rect 13636 39788 13688 39840
rect 15384 39924 15436 39976
rect 15936 40035 15988 40044
rect 15936 40001 15946 40035
rect 15946 40001 15980 40035
rect 15980 40001 15988 40035
rect 15936 39992 15988 40001
rect 16120 40035 16172 40044
rect 16120 40001 16129 40035
rect 16129 40001 16163 40035
rect 16163 40001 16172 40035
rect 16120 39992 16172 40001
rect 16212 40035 16264 40044
rect 16212 40001 16221 40035
rect 16221 40001 16255 40035
rect 16255 40001 16264 40035
rect 16212 39992 16264 40001
rect 16028 39924 16080 39976
rect 17132 39992 17184 40044
rect 16948 39856 17000 39908
rect 20720 39992 20772 40044
rect 20904 40060 20956 40112
rect 23480 39992 23532 40044
rect 27620 40103 27672 40112
rect 27620 40069 27629 40103
rect 27629 40069 27663 40103
rect 27663 40069 27672 40103
rect 27620 40060 27672 40069
rect 20904 39967 20956 39976
rect 20904 39933 20913 39967
rect 20913 39933 20947 39967
rect 20947 39933 20956 39967
rect 20904 39924 20956 39933
rect 27160 40035 27212 40044
rect 27160 40001 27169 40035
rect 27169 40001 27203 40035
rect 27203 40001 27212 40035
rect 27160 39992 27212 40001
rect 27344 40035 27396 40044
rect 27344 40001 27353 40035
rect 27353 40001 27387 40035
rect 27387 40001 27396 40035
rect 27344 39992 27396 40001
rect 27896 39992 27948 40044
rect 30932 40060 30984 40112
rect 24584 39924 24636 39976
rect 26884 39924 26936 39976
rect 28264 39924 28316 39976
rect 34060 40060 34112 40112
rect 34336 39992 34388 40044
rect 40500 40060 40552 40112
rect 35900 39992 35952 40044
rect 40684 39992 40736 40044
rect 34428 39924 34480 39976
rect 35440 39924 35492 39976
rect 38016 39924 38068 39976
rect 39120 39967 39172 39976
rect 39120 39933 39129 39967
rect 39129 39933 39163 39967
rect 39163 39933 39172 39967
rect 39120 39924 39172 39933
rect 17592 39831 17644 39840
rect 17592 39797 17601 39831
rect 17601 39797 17635 39831
rect 17635 39797 17644 39831
rect 17592 39788 17644 39797
rect 18328 39788 18380 39840
rect 18788 39831 18840 39840
rect 18788 39797 18797 39831
rect 18797 39797 18831 39831
rect 18831 39797 18840 39831
rect 18788 39788 18840 39797
rect 21088 39788 21140 39840
rect 21548 39831 21600 39840
rect 21548 39797 21557 39831
rect 21557 39797 21591 39831
rect 21591 39797 21600 39831
rect 21548 39788 21600 39797
rect 23664 39788 23716 39840
rect 26332 39788 26384 39840
rect 26516 39788 26568 39840
rect 27528 39856 27580 39908
rect 30288 39788 30340 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3976 39584 4028 39636
rect 6184 39584 6236 39636
rect 6644 39584 6696 39636
rect 8024 39584 8076 39636
rect 8576 39584 8628 39636
rect 9772 39584 9824 39636
rect 12440 39584 12492 39636
rect 13544 39584 13596 39636
rect 4528 39516 4580 39568
rect 4804 39516 4856 39568
rect 8208 39516 8260 39568
rect 17132 39584 17184 39636
rect 20904 39584 20956 39636
rect 27528 39584 27580 39636
rect 27896 39584 27948 39636
rect 2596 39380 2648 39432
rect 6368 39448 6420 39500
rect 2504 39287 2556 39296
rect 2504 39253 2513 39287
rect 2513 39253 2547 39287
rect 2547 39253 2556 39287
rect 2504 39244 2556 39253
rect 3148 39244 3200 39296
rect 5908 39244 5960 39296
rect 8116 39380 8168 39432
rect 8024 39355 8076 39364
rect 8024 39321 8033 39355
rect 8033 39321 8067 39355
rect 8067 39321 8076 39355
rect 8024 39312 8076 39321
rect 8300 39423 8352 39432
rect 8300 39389 8309 39423
rect 8309 39389 8343 39423
rect 8343 39389 8352 39423
rect 8300 39380 8352 39389
rect 8392 39380 8444 39432
rect 8944 39423 8996 39432
rect 8944 39389 8953 39423
rect 8953 39389 8987 39423
rect 8987 39389 8996 39423
rect 8944 39380 8996 39389
rect 9036 39380 9088 39432
rect 18328 39516 18380 39568
rect 20352 39516 20404 39568
rect 10048 39491 10100 39500
rect 10048 39457 10057 39491
rect 10057 39457 10091 39491
rect 10091 39457 10100 39491
rect 10048 39448 10100 39457
rect 13636 39448 13688 39500
rect 15384 39491 15436 39500
rect 15384 39457 15393 39491
rect 15393 39457 15427 39491
rect 15427 39457 15436 39491
rect 15384 39448 15436 39457
rect 21640 39448 21692 39500
rect 24400 39491 24452 39500
rect 24400 39457 24409 39491
rect 24409 39457 24443 39491
rect 24443 39457 24452 39491
rect 24400 39448 24452 39457
rect 26792 39491 26844 39500
rect 26792 39457 26801 39491
rect 26801 39457 26835 39491
rect 26835 39457 26844 39491
rect 26792 39448 26844 39457
rect 30288 39516 30340 39568
rect 30012 39448 30064 39500
rect 10784 39380 10836 39432
rect 15108 39423 15160 39432
rect 15108 39389 15117 39423
rect 15117 39389 15151 39423
rect 15151 39389 15160 39423
rect 15108 39380 15160 39389
rect 17684 39423 17736 39432
rect 17684 39389 17693 39423
rect 17693 39389 17727 39423
rect 17727 39389 17736 39423
rect 17684 39380 17736 39389
rect 19432 39380 19484 39432
rect 22284 39423 22336 39432
rect 22284 39389 22293 39423
rect 22293 39389 22327 39423
rect 22327 39389 22336 39423
rect 22284 39380 22336 39389
rect 26424 39423 26476 39432
rect 26424 39389 26433 39423
rect 26433 39389 26467 39423
rect 26467 39389 26476 39423
rect 26424 39380 26476 39389
rect 29828 39423 29880 39432
rect 29828 39389 29837 39423
rect 29837 39389 29871 39423
rect 29871 39389 29880 39423
rect 29828 39380 29880 39389
rect 30380 39448 30432 39500
rect 32220 39491 32272 39500
rect 32220 39457 32229 39491
rect 32229 39457 32263 39491
rect 32263 39457 32272 39491
rect 32220 39448 32272 39457
rect 39304 39448 39356 39500
rect 30196 39380 30248 39432
rect 11520 39312 11572 39364
rect 14188 39312 14240 39364
rect 8116 39244 8168 39296
rect 8484 39244 8536 39296
rect 9036 39244 9088 39296
rect 13820 39287 13872 39296
rect 13820 39253 13829 39287
rect 13829 39253 13863 39287
rect 13863 39253 13872 39287
rect 13820 39244 13872 39253
rect 19984 39312 20036 39364
rect 17040 39244 17092 39296
rect 19156 39244 19208 39296
rect 20260 39287 20312 39296
rect 20260 39253 20269 39287
rect 20269 39253 20303 39287
rect 20303 39253 20312 39287
rect 20260 39244 20312 39253
rect 20720 39312 20772 39364
rect 22008 39355 22060 39364
rect 22008 39321 22017 39355
rect 22017 39321 22051 39355
rect 22051 39321 22060 39355
rect 22008 39312 22060 39321
rect 22652 39312 22704 39364
rect 24676 39355 24728 39364
rect 24676 39321 24685 39355
rect 24685 39321 24719 39355
rect 24719 39321 24728 39355
rect 24676 39312 24728 39321
rect 35624 39423 35676 39432
rect 35624 39389 35633 39423
rect 35633 39389 35667 39423
rect 35667 39389 35676 39423
rect 35624 39380 35676 39389
rect 35992 39423 36044 39432
rect 35992 39389 36001 39423
rect 36001 39389 36035 39423
rect 36035 39389 36044 39423
rect 35992 39380 36044 39389
rect 38016 39423 38068 39432
rect 38016 39389 38025 39423
rect 38025 39389 38059 39423
rect 38059 39389 38068 39423
rect 38016 39380 38068 39389
rect 38292 39380 38344 39432
rect 42064 39448 42116 39500
rect 21088 39244 21140 39296
rect 21180 39244 21232 39296
rect 23388 39244 23440 39296
rect 25688 39244 25740 39296
rect 26332 39287 26384 39296
rect 26332 39253 26341 39287
rect 26341 39253 26375 39287
rect 26375 39253 26384 39287
rect 26332 39244 26384 39253
rect 30012 39287 30064 39296
rect 30012 39253 30021 39287
rect 30021 39253 30055 39287
rect 30055 39253 30064 39287
rect 30012 39244 30064 39253
rect 30472 39287 30524 39296
rect 30472 39253 30481 39287
rect 30481 39253 30515 39287
rect 30515 39253 30524 39287
rect 30472 39244 30524 39253
rect 31484 39312 31536 39364
rect 35808 39355 35860 39364
rect 35808 39321 35817 39355
rect 35817 39321 35851 39355
rect 35851 39321 35860 39355
rect 35808 39312 35860 39321
rect 35900 39355 35952 39364
rect 35900 39321 35909 39355
rect 35909 39321 35943 39355
rect 35943 39321 35952 39355
rect 35900 39312 35952 39321
rect 37188 39312 37240 39364
rect 38752 39312 38804 39364
rect 39856 39423 39908 39432
rect 39856 39389 39865 39423
rect 39865 39389 39899 39423
rect 39899 39389 39908 39423
rect 39856 39380 39908 39389
rect 41788 39380 41840 39432
rect 40132 39355 40184 39364
rect 40132 39321 40141 39355
rect 40141 39321 40175 39355
rect 40175 39321 40184 39355
rect 40132 39312 40184 39321
rect 40684 39312 40736 39364
rect 34152 39244 34204 39296
rect 34336 39244 34388 39296
rect 36268 39287 36320 39296
rect 36268 39253 36277 39287
rect 36277 39253 36311 39287
rect 36311 39253 36320 39287
rect 36268 39244 36320 39253
rect 39488 39244 39540 39296
rect 40040 39244 40092 39296
rect 41696 39287 41748 39296
rect 41696 39253 41705 39287
rect 41705 39253 41739 39287
rect 41739 39253 41748 39287
rect 41696 39244 41748 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 2596 39083 2648 39092
rect 2596 39049 2605 39083
rect 2605 39049 2639 39083
rect 2639 39049 2648 39083
rect 2596 39040 2648 39049
rect 4620 39040 4672 39092
rect 8484 39040 8536 39092
rect 11520 39083 11572 39092
rect 11520 39049 11529 39083
rect 11529 39049 11563 39083
rect 11563 39049 11572 39083
rect 11520 39040 11572 39049
rect 11888 39040 11940 39092
rect 12992 39083 13044 39092
rect 12992 39049 13001 39083
rect 13001 39049 13035 39083
rect 13035 39049 13044 39083
rect 12992 39040 13044 39049
rect 13820 39040 13872 39092
rect 14188 39083 14240 39092
rect 14188 39049 14197 39083
rect 14197 39049 14231 39083
rect 14231 39049 14240 39083
rect 14188 39040 14240 39049
rect 15108 39040 15160 39092
rect 16212 39040 16264 39092
rect 17592 39040 17644 39092
rect 2872 38904 2924 38956
rect 3148 38879 3200 38888
rect 3148 38845 3157 38879
rect 3157 38845 3191 38879
rect 3191 38845 3200 38879
rect 3148 38836 3200 38845
rect 3976 38879 4028 38888
rect 3976 38845 3985 38879
rect 3985 38845 4019 38879
rect 4019 38845 4028 38879
rect 3976 38836 4028 38845
rect 4528 38947 4580 38956
rect 4528 38913 4537 38947
rect 4537 38913 4571 38947
rect 4571 38913 4580 38947
rect 4528 38904 4580 38913
rect 6092 38972 6144 39024
rect 8208 38972 8260 39024
rect 12348 38972 12400 39024
rect 8392 38904 8444 38956
rect 10048 38947 10100 38956
rect 10048 38913 10057 38947
rect 10057 38913 10091 38947
rect 10091 38913 10100 38947
rect 10048 38904 10100 38913
rect 4988 38836 5040 38888
rect 4712 38768 4764 38820
rect 5908 38768 5960 38820
rect 9404 38879 9456 38888
rect 9404 38845 9413 38879
rect 9413 38845 9447 38879
rect 9447 38845 9456 38879
rect 9404 38836 9456 38845
rect 12164 38836 12216 38888
rect 16396 38904 16448 38956
rect 17040 38947 17092 38956
rect 17040 38913 17049 38947
rect 17049 38913 17083 38947
rect 17083 38913 17092 38947
rect 17040 38904 17092 38913
rect 5264 38700 5316 38752
rect 8208 38743 8260 38752
rect 8208 38709 8217 38743
rect 8217 38709 8251 38743
rect 8251 38709 8260 38743
rect 8208 38700 8260 38709
rect 17408 38836 17460 38888
rect 16580 38700 16632 38752
rect 17868 38972 17920 39024
rect 18788 38972 18840 39024
rect 19984 39040 20036 39092
rect 20168 39083 20220 39092
rect 20168 39049 20177 39083
rect 20177 39049 20211 39083
rect 20211 39049 20220 39083
rect 20168 39040 20220 39049
rect 20260 39040 20312 39092
rect 20352 39040 20404 39092
rect 17592 38768 17644 38820
rect 18604 38904 18656 38956
rect 19432 38904 19484 38956
rect 20904 39040 20956 39092
rect 21088 39040 21140 39092
rect 21548 39040 21600 39092
rect 21640 39040 21692 39092
rect 22008 39040 22060 39092
rect 24676 39040 24728 39092
rect 26332 39040 26384 39092
rect 26424 39040 26476 39092
rect 27620 39040 27672 39092
rect 28264 39083 28316 39092
rect 28264 39049 28273 39083
rect 28273 39049 28307 39083
rect 28307 39049 28316 39083
rect 28264 39040 28316 39049
rect 29828 39040 29880 39092
rect 30012 39040 30064 39092
rect 30472 39040 30524 39092
rect 30564 39040 30616 39092
rect 32404 39083 32456 39092
rect 32404 39049 32413 39083
rect 32413 39049 32447 39083
rect 32447 39049 32456 39083
rect 32404 39040 32456 39049
rect 20904 38947 20956 38956
rect 20904 38913 20908 38947
rect 20908 38913 20942 38947
rect 20942 38913 20956 38947
rect 20904 38904 20956 38913
rect 20996 38947 21048 38956
rect 20996 38913 21005 38947
rect 21005 38913 21039 38947
rect 21039 38913 21048 38947
rect 20996 38904 21048 38913
rect 24584 38972 24636 39024
rect 20352 38768 20404 38820
rect 23480 38836 23532 38888
rect 23572 38879 23624 38888
rect 23572 38845 23581 38879
rect 23581 38845 23615 38879
rect 23615 38845 23624 38879
rect 23572 38836 23624 38845
rect 23756 38904 23808 38956
rect 24124 38836 24176 38888
rect 27528 38947 27580 38956
rect 27528 38913 27537 38947
rect 27537 38913 27571 38947
rect 27571 38913 27580 38947
rect 27528 38904 27580 38913
rect 21180 38768 21232 38820
rect 23388 38768 23440 38820
rect 24768 38768 24820 38820
rect 26516 38768 26568 38820
rect 29920 39015 29972 39024
rect 29920 38981 29929 39015
rect 29929 38981 29963 39015
rect 29963 38981 29972 39015
rect 29920 38972 29972 38981
rect 35440 39083 35492 39092
rect 35440 39049 35449 39083
rect 35449 39049 35483 39083
rect 35483 39049 35492 39083
rect 35440 39040 35492 39049
rect 35900 39040 35952 39092
rect 28172 38904 28224 38956
rect 28908 38904 28960 38956
rect 30104 38904 30156 38956
rect 31208 38904 31260 38956
rect 32864 38947 32916 38956
rect 32864 38913 32873 38947
rect 32873 38913 32907 38947
rect 32907 38913 32916 38947
rect 32864 38904 32916 38913
rect 33048 38904 33100 38956
rect 33600 39015 33652 39024
rect 33600 38981 33609 39015
rect 33609 38981 33643 39015
rect 33643 38981 33652 39015
rect 33600 38972 33652 38981
rect 33876 38972 33928 39024
rect 39396 38972 39448 39024
rect 40684 38972 40736 39024
rect 33416 38904 33468 38956
rect 34060 38947 34112 38956
rect 34060 38913 34069 38947
rect 34069 38913 34103 38947
rect 34103 38913 34112 38947
rect 34060 38904 34112 38913
rect 34336 38904 34388 38956
rect 20904 38700 20956 38752
rect 22836 38700 22888 38752
rect 26240 38700 26292 38752
rect 27804 38700 27856 38752
rect 29736 38700 29788 38752
rect 30564 38743 30616 38752
rect 30564 38709 30573 38743
rect 30573 38709 30607 38743
rect 30607 38709 30616 38743
rect 30564 38700 30616 38709
rect 33140 38768 33192 38820
rect 33324 38768 33376 38820
rect 33508 38700 33560 38752
rect 34152 38879 34204 38888
rect 34152 38845 34161 38879
rect 34161 38845 34195 38879
rect 34195 38845 34204 38879
rect 34152 38836 34204 38845
rect 35256 38904 35308 38956
rect 34704 38836 34756 38888
rect 35624 38904 35676 38956
rect 35716 38947 35768 38956
rect 35716 38913 35725 38947
rect 35725 38913 35759 38947
rect 35759 38913 35768 38947
rect 35716 38904 35768 38913
rect 36268 38904 36320 38956
rect 37004 38904 37056 38956
rect 38660 38904 38712 38956
rect 39856 38904 39908 38956
rect 35532 38836 35584 38888
rect 39764 38879 39816 38888
rect 39764 38845 39773 38879
rect 39773 38845 39807 38879
rect 39807 38845 39816 38879
rect 39764 38836 39816 38845
rect 40224 38879 40276 38888
rect 40224 38845 40233 38879
rect 40233 38845 40267 38879
rect 40267 38845 40276 38879
rect 40224 38836 40276 38845
rect 38292 38768 38344 38820
rect 34060 38743 34112 38752
rect 34060 38709 34069 38743
rect 34069 38709 34103 38743
rect 34103 38709 34112 38743
rect 34060 38700 34112 38709
rect 34796 38700 34848 38752
rect 37280 38700 37332 38752
rect 38016 38700 38068 38752
rect 38752 38700 38804 38752
rect 41788 38700 41840 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 3976 38496 4028 38548
rect 5080 38539 5132 38548
rect 5080 38505 5089 38539
rect 5089 38505 5123 38539
rect 5123 38505 5132 38539
rect 5080 38496 5132 38505
rect 9404 38496 9456 38548
rect 17684 38496 17736 38548
rect 18604 38539 18656 38548
rect 18604 38505 18613 38539
rect 18613 38505 18647 38539
rect 18647 38505 18656 38539
rect 18604 38496 18656 38505
rect 23480 38496 23532 38548
rect 5264 38360 5316 38412
rect 10784 38360 10836 38412
rect 15384 38360 15436 38412
rect 17408 38403 17460 38412
rect 17408 38369 17417 38403
rect 17417 38369 17451 38403
rect 17451 38369 17460 38403
rect 17408 38360 17460 38369
rect 1492 38292 1544 38344
rect 6920 38292 6972 38344
rect 8208 38292 8260 38344
rect 9220 38335 9272 38344
rect 9220 38301 9229 38335
rect 9229 38301 9263 38335
rect 9263 38301 9272 38335
rect 9220 38292 9272 38301
rect 17316 38292 17368 38344
rect 18236 38335 18288 38344
rect 18236 38301 18245 38335
rect 18245 38301 18279 38335
rect 18279 38301 18288 38335
rect 19156 38360 19208 38412
rect 18236 38292 18288 38301
rect 18788 38335 18840 38344
rect 18788 38301 18797 38335
rect 18797 38301 18831 38335
rect 18831 38301 18840 38335
rect 18788 38292 18840 38301
rect 19248 38292 19300 38344
rect 21456 38292 21508 38344
rect 22284 38360 22336 38412
rect 22836 38360 22888 38412
rect 30380 38496 30432 38548
rect 33140 38496 33192 38548
rect 33968 38496 34020 38548
rect 34704 38496 34756 38548
rect 35348 38496 35400 38548
rect 35716 38496 35768 38548
rect 35992 38496 36044 38548
rect 37004 38496 37056 38548
rect 39120 38539 39172 38548
rect 39120 38505 39129 38539
rect 39129 38505 39163 38539
rect 39163 38505 39172 38539
rect 39120 38496 39172 38505
rect 40224 38496 40276 38548
rect 2136 38224 2188 38276
rect 7012 38224 7064 38276
rect 4620 38156 4672 38208
rect 10232 38224 10284 38276
rect 15936 38267 15988 38276
rect 15936 38233 15970 38267
rect 15970 38233 15988 38267
rect 15936 38224 15988 38233
rect 25688 38360 25740 38412
rect 26056 38360 26108 38412
rect 25504 38335 25556 38344
rect 25504 38301 25513 38335
rect 25513 38301 25547 38335
rect 25547 38301 25556 38335
rect 25504 38292 25556 38301
rect 29736 38335 29788 38344
rect 29736 38301 29745 38335
rect 29745 38301 29779 38335
rect 29779 38301 29788 38335
rect 29736 38292 29788 38301
rect 33324 38360 33376 38412
rect 30012 38292 30064 38344
rect 30564 38292 30616 38344
rect 30840 38335 30892 38344
rect 30840 38301 30849 38335
rect 30849 38301 30883 38335
rect 30883 38301 30892 38335
rect 30840 38292 30892 38301
rect 30932 38292 30984 38344
rect 32404 38292 32456 38344
rect 11244 38199 11296 38208
rect 11244 38165 11253 38199
rect 11253 38165 11287 38199
rect 11287 38165 11296 38199
rect 11244 38156 11296 38165
rect 17776 38199 17828 38208
rect 17776 38165 17785 38199
rect 17785 38165 17819 38199
rect 17819 38165 17828 38199
rect 17776 38156 17828 38165
rect 18144 38199 18196 38208
rect 18144 38165 18153 38199
rect 18153 38165 18187 38199
rect 18187 38165 18196 38199
rect 18144 38156 18196 38165
rect 29368 38224 29420 38276
rect 29644 38224 29696 38276
rect 33416 38335 33468 38344
rect 33416 38301 33425 38335
rect 33425 38301 33459 38335
rect 33459 38301 33468 38335
rect 33416 38292 33468 38301
rect 33508 38292 33560 38344
rect 33692 38292 33744 38344
rect 34060 38292 34112 38344
rect 34428 38292 34480 38344
rect 34796 38292 34848 38344
rect 35348 38335 35400 38344
rect 35348 38301 35357 38335
rect 35357 38301 35391 38335
rect 35391 38301 35400 38335
rect 35348 38292 35400 38301
rect 39764 38428 39816 38480
rect 35532 38224 35584 38276
rect 36544 38292 36596 38344
rect 38292 38360 38344 38412
rect 37004 38335 37056 38344
rect 37004 38301 37037 38335
rect 37037 38301 37056 38335
rect 37004 38292 37056 38301
rect 37280 38335 37332 38344
rect 37280 38301 37289 38335
rect 37289 38301 37323 38335
rect 37323 38301 37332 38335
rect 37280 38292 37332 38301
rect 39212 38360 39264 38412
rect 40040 38403 40092 38412
rect 40040 38369 40049 38403
rect 40049 38369 40083 38403
rect 40083 38369 40092 38403
rect 40040 38360 40092 38369
rect 40684 38360 40736 38412
rect 39304 38335 39356 38344
rect 39304 38301 39313 38335
rect 39313 38301 39347 38335
rect 39347 38301 39356 38335
rect 39304 38292 39356 38301
rect 36360 38224 36412 38276
rect 24400 38199 24452 38208
rect 24400 38165 24409 38199
rect 24409 38165 24443 38199
rect 24443 38165 24452 38199
rect 24400 38156 24452 38165
rect 25504 38156 25556 38208
rect 26424 38156 26476 38208
rect 27528 38156 27580 38208
rect 29092 38156 29144 38208
rect 32772 38156 32824 38208
rect 33232 38156 33284 38208
rect 33508 38156 33560 38208
rect 34796 38156 34848 38208
rect 35348 38156 35400 38208
rect 36452 38199 36504 38208
rect 36452 38165 36461 38199
rect 36461 38165 36495 38199
rect 36495 38165 36504 38199
rect 36452 38156 36504 38165
rect 38936 38156 38988 38208
rect 39580 38224 39632 38276
rect 40316 38292 40368 38344
rect 40500 38292 40552 38344
rect 42064 38335 42116 38344
rect 42064 38301 42073 38335
rect 42073 38301 42107 38335
rect 42107 38301 42116 38335
rect 42064 38292 42116 38301
rect 40224 38224 40276 38276
rect 41328 38156 41380 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 2136 37995 2188 38004
rect 2136 37961 2145 37995
rect 2145 37961 2179 37995
rect 2179 37961 2188 37995
rect 2136 37952 2188 37961
rect 2504 37952 2556 38004
rect 5264 37952 5316 38004
rect 6736 37995 6788 38004
rect 6736 37961 6745 37995
rect 6745 37961 6779 37995
rect 6779 37961 6788 37995
rect 6736 37952 6788 37961
rect 8944 37952 8996 38004
rect 9036 37995 9088 38004
rect 9036 37961 9045 37995
rect 9045 37961 9079 37995
rect 9079 37961 9088 37995
rect 9036 37952 9088 37961
rect 9128 37952 9180 38004
rect 9220 37952 9272 38004
rect 10048 37995 10100 38004
rect 10048 37961 10057 37995
rect 10057 37961 10091 37995
rect 10091 37961 10100 37995
rect 10048 37952 10100 37961
rect 2780 37859 2832 37868
rect 2780 37825 2789 37859
rect 2789 37825 2823 37859
rect 2823 37825 2832 37859
rect 2780 37816 2832 37825
rect 1492 37748 1544 37800
rect 3608 37816 3660 37868
rect 4896 37859 4948 37868
rect 4896 37825 4930 37859
rect 4930 37825 4948 37859
rect 4896 37816 4948 37825
rect 5448 37816 5500 37868
rect 7472 37859 7524 37868
rect 7472 37825 7506 37859
rect 7506 37825 7524 37859
rect 7472 37816 7524 37825
rect 11244 37884 11296 37936
rect 12532 37884 12584 37936
rect 15200 37952 15252 38004
rect 15844 37952 15896 38004
rect 15936 37995 15988 38004
rect 15936 37961 15945 37995
rect 15945 37961 15979 37995
rect 15979 37961 15988 37995
rect 15936 37952 15988 37961
rect 17960 37952 18012 38004
rect 19248 37952 19300 38004
rect 21456 37952 21508 38004
rect 23572 37952 23624 38004
rect 24400 37952 24452 38004
rect 15476 37884 15528 37936
rect 20812 37884 20864 37936
rect 29092 37952 29144 38004
rect 6828 37748 6880 37800
rect 6920 37680 6972 37732
rect 9128 37791 9180 37800
rect 9128 37757 9137 37791
rect 9137 37757 9171 37791
rect 9171 37757 9180 37791
rect 9128 37748 9180 37757
rect 9404 37748 9456 37800
rect 12808 37748 12860 37800
rect 6000 37655 6052 37664
rect 6000 37621 6009 37655
rect 6009 37621 6043 37655
rect 6043 37621 6052 37655
rect 6000 37612 6052 37621
rect 6184 37612 6236 37664
rect 7104 37655 7156 37664
rect 7104 37621 7113 37655
rect 7113 37621 7147 37655
rect 7147 37621 7156 37655
rect 7104 37612 7156 37621
rect 8668 37655 8720 37664
rect 8668 37621 8677 37655
rect 8677 37621 8711 37655
rect 8711 37621 8720 37655
rect 8668 37612 8720 37621
rect 13360 37612 13412 37664
rect 15200 37816 15252 37868
rect 15660 37816 15712 37868
rect 16580 37816 16632 37868
rect 17684 37859 17736 37868
rect 17684 37825 17718 37859
rect 17718 37825 17736 37859
rect 14188 37791 14240 37800
rect 14188 37757 14197 37791
rect 14197 37757 14231 37791
rect 14231 37757 14240 37791
rect 14188 37748 14240 37757
rect 14556 37748 14608 37800
rect 15200 37680 15252 37732
rect 17684 37816 17736 37825
rect 23388 37859 23440 37868
rect 23388 37825 23392 37859
rect 23392 37825 23426 37859
rect 23426 37825 23440 37859
rect 23388 37816 23440 37825
rect 23480 37859 23532 37868
rect 23480 37825 23489 37859
rect 23489 37825 23523 37859
rect 23523 37825 23532 37859
rect 23480 37816 23532 37825
rect 23664 37816 23716 37868
rect 30840 37952 30892 38004
rect 33692 37952 33744 38004
rect 24124 37859 24176 37868
rect 24124 37825 24133 37859
rect 24133 37825 24167 37859
rect 24167 37825 24176 37859
rect 24124 37816 24176 37825
rect 25504 37816 25556 37868
rect 25044 37748 25096 37800
rect 25136 37791 25188 37800
rect 25136 37757 25145 37791
rect 25145 37757 25179 37791
rect 25179 37757 25188 37791
rect 25136 37748 25188 37757
rect 27804 37748 27856 37800
rect 29092 37748 29144 37800
rect 30380 37859 30432 37868
rect 30380 37825 30389 37859
rect 30389 37825 30423 37859
rect 30423 37825 30432 37859
rect 30380 37816 30432 37825
rect 40040 37952 40092 38004
rect 41880 37952 41932 38004
rect 39580 37884 39632 37936
rect 32404 37816 32456 37868
rect 32772 37816 32824 37868
rect 38292 37816 38344 37868
rect 35532 37748 35584 37800
rect 37280 37748 37332 37800
rect 37372 37748 37424 37800
rect 38568 37791 38620 37800
rect 38568 37757 38577 37791
rect 38577 37757 38611 37791
rect 38611 37757 38620 37791
rect 38568 37748 38620 37757
rect 38936 37816 38988 37868
rect 39120 37859 39172 37868
rect 39120 37825 39129 37859
rect 39129 37825 39163 37859
rect 39163 37825 39172 37859
rect 39120 37816 39172 37825
rect 39304 37816 39356 37868
rect 40132 37859 40184 37868
rect 40132 37825 40141 37859
rect 40141 37825 40175 37859
rect 40175 37825 40184 37859
rect 40132 37816 40184 37825
rect 40316 37748 40368 37800
rect 41696 37816 41748 37868
rect 41788 37816 41840 37868
rect 43260 37816 43312 37868
rect 44180 37748 44232 37800
rect 44456 37791 44508 37800
rect 44456 37757 44465 37791
rect 44465 37757 44499 37791
rect 44499 37757 44508 37791
rect 44456 37748 44508 37757
rect 42064 37680 42116 37732
rect 42800 37680 42852 37732
rect 17592 37612 17644 37664
rect 25688 37612 25740 37664
rect 30012 37655 30064 37664
rect 30012 37621 30021 37655
rect 30021 37621 30055 37655
rect 30055 37621 30064 37655
rect 30012 37612 30064 37621
rect 30564 37655 30616 37664
rect 30564 37621 30573 37655
rect 30573 37621 30607 37655
rect 30607 37621 30616 37655
rect 30564 37612 30616 37621
rect 33232 37612 33284 37664
rect 36544 37612 36596 37664
rect 37648 37612 37700 37664
rect 38752 37655 38804 37664
rect 38752 37621 38761 37655
rect 38761 37621 38795 37655
rect 38795 37621 38804 37655
rect 38752 37612 38804 37621
rect 39672 37612 39724 37664
rect 41512 37612 41564 37664
rect 43076 37655 43128 37664
rect 43076 37621 43085 37655
rect 43085 37621 43119 37655
rect 43119 37621 43128 37655
rect 43076 37612 43128 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2780 37408 2832 37460
rect 4896 37408 4948 37460
rect 6276 37408 6328 37460
rect 6736 37408 6788 37460
rect 7012 37408 7064 37460
rect 7472 37408 7524 37460
rect 12532 37408 12584 37460
rect 17684 37451 17736 37460
rect 17684 37417 17693 37451
rect 17693 37417 17727 37451
rect 17727 37417 17736 37451
rect 17684 37408 17736 37417
rect 18788 37408 18840 37460
rect 2872 37315 2924 37324
rect 2872 37281 2881 37315
rect 2881 37281 2915 37315
rect 2915 37281 2924 37315
rect 2872 37272 2924 37281
rect 4804 37272 4856 37324
rect 5448 37272 5500 37324
rect 5908 37315 5960 37324
rect 5908 37281 5917 37315
rect 5917 37281 5951 37315
rect 5951 37281 5960 37315
rect 5908 37272 5960 37281
rect 6000 37272 6052 37324
rect 20444 37408 20496 37460
rect 27528 37408 27580 37460
rect 28908 37451 28960 37460
rect 28908 37417 28917 37451
rect 28917 37417 28951 37451
rect 28951 37417 28960 37451
rect 28908 37408 28960 37417
rect 33232 37451 33284 37460
rect 33232 37417 33241 37451
rect 33241 37417 33275 37451
rect 33275 37417 33284 37451
rect 33232 37408 33284 37417
rect 36360 37408 36412 37460
rect 36820 37408 36872 37460
rect 38292 37408 38344 37460
rect 21456 37315 21508 37324
rect 21456 37281 21465 37315
rect 21465 37281 21499 37315
rect 21499 37281 21508 37315
rect 21456 37272 21508 37281
rect 25688 37272 25740 37324
rect 26056 37272 26108 37324
rect 27068 37315 27120 37324
rect 27068 37281 27077 37315
rect 27077 37281 27111 37315
rect 27111 37281 27120 37315
rect 27068 37272 27120 37281
rect 940 37204 992 37256
rect 1584 37111 1636 37120
rect 1584 37077 1593 37111
rect 1593 37077 1627 37111
rect 1627 37077 1636 37111
rect 1584 37068 1636 37077
rect 1952 37111 2004 37120
rect 1952 37077 1961 37111
rect 1961 37077 1995 37111
rect 1995 37077 2004 37111
rect 1952 37068 2004 37077
rect 4620 37204 4672 37256
rect 2780 37111 2832 37120
rect 2780 37077 2789 37111
rect 2789 37077 2823 37111
rect 2823 37077 2832 37111
rect 2780 37068 2832 37077
rect 4988 37068 5040 37120
rect 7104 37247 7156 37256
rect 7104 37213 7113 37247
rect 7113 37213 7147 37247
rect 7147 37213 7156 37247
rect 7104 37204 7156 37213
rect 8668 37204 8720 37256
rect 12808 37204 12860 37256
rect 15844 37204 15896 37256
rect 17776 37204 17828 37256
rect 18512 37204 18564 37256
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 23480 37247 23532 37256
rect 5908 37136 5960 37188
rect 13728 37068 13780 37120
rect 18236 37068 18288 37120
rect 20812 37136 20864 37188
rect 20996 37068 21048 37120
rect 22284 37068 22336 37120
rect 22468 37068 22520 37120
rect 23480 37213 23489 37247
rect 23489 37213 23523 37247
rect 23523 37213 23532 37247
rect 23480 37204 23532 37213
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 25228 37204 25280 37256
rect 22928 37111 22980 37120
rect 22928 37077 22937 37111
rect 22937 37077 22971 37111
rect 22971 37077 22980 37111
rect 22928 37068 22980 37077
rect 24860 37068 24912 37120
rect 26056 37136 26108 37188
rect 30564 37272 30616 37324
rect 27436 37179 27488 37188
rect 27436 37145 27445 37179
rect 27445 37145 27479 37179
rect 27479 37145 27488 37179
rect 27436 37136 27488 37145
rect 30012 37247 30064 37256
rect 30012 37213 30021 37247
rect 30021 37213 30055 37247
rect 30055 37213 30064 37247
rect 30012 37204 30064 37213
rect 35532 37315 35584 37324
rect 35532 37281 35541 37315
rect 35541 37281 35575 37315
rect 35575 37281 35584 37315
rect 35532 37272 35584 37281
rect 35900 37272 35952 37324
rect 36452 37272 36504 37324
rect 37004 37272 37056 37324
rect 32404 37204 32456 37256
rect 32772 37247 32824 37256
rect 32772 37213 32781 37247
rect 32781 37213 32815 37247
rect 32815 37213 32824 37247
rect 32772 37204 32824 37213
rect 33140 37204 33192 37256
rect 38016 37204 38068 37256
rect 39120 37408 39172 37460
rect 39304 37408 39356 37460
rect 44456 37408 44508 37460
rect 43076 37272 43128 37324
rect 42432 37247 42484 37256
rect 29092 37068 29144 37120
rect 29920 37111 29972 37120
rect 29920 37077 29929 37111
rect 29929 37077 29963 37111
rect 29963 37077 29972 37111
rect 29920 37068 29972 37077
rect 30288 37068 30340 37120
rect 30840 37068 30892 37120
rect 37280 37111 37332 37120
rect 37280 37077 37289 37111
rect 37289 37077 37323 37111
rect 37323 37077 37332 37111
rect 37280 37068 37332 37077
rect 38292 37179 38344 37188
rect 38292 37145 38301 37179
rect 38301 37145 38335 37179
rect 38335 37145 38344 37179
rect 38292 37136 38344 37145
rect 38384 37179 38436 37188
rect 38384 37145 38393 37179
rect 38393 37145 38427 37179
rect 38427 37145 38436 37179
rect 38384 37136 38436 37145
rect 39212 37136 39264 37188
rect 39580 37136 39632 37188
rect 39948 37136 40000 37188
rect 38660 37111 38712 37120
rect 38660 37077 38669 37111
rect 38669 37077 38703 37111
rect 38703 37077 38712 37111
rect 38660 37068 38712 37077
rect 39488 37068 39540 37120
rect 39856 37068 39908 37120
rect 42432 37213 42441 37247
rect 42441 37213 42475 37247
rect 42475 37213 42484 37247
rect 42432 37204 42484 37213
rect 43720 37068 43772 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1952 36864 2004 36916
rect 2780 36864 2832 36916
rect 12808 36907 12860 36916
rect 12808 36873 12817 36907
rect 12817 36873 12851 36907
rect 12851 36873 12860 36907
rect 12808 36864 12860 36873
rect 14188 36864 14240 36916
rect 17040 36864 17092 36916
rect 19248 36864 19300 36916
rect 20812 36907 20864 36916
rect 20812 36873 20821 36907
rect 20821 36873 20855 36907
rect 20855 36873 20864 36907
rect 20812 36864 20864 36873
rect 22928 36864 22980 36916
rect 24400 36864 24452 36916
rect 25136 36864 25188 36916
rect 27436 36864 27488 36916
rect 29276 36864 29328 36916
rect 29828 36864 29880 36916
rect 29920 36864 29972 36916
rect 5540 36796 5592 36848
rect 6368 36839 6420 36848
rect 6368 36805 6377 36839
rect 6377 36805 6411 36839
rect 6411 36805 6420 36839
rect 6368 36796 6420 36805
rect 1492 36771 1544 36780
rect 1492 36737 1501 36771
rect 1501 36737 1535 36771
rect 1535 36737 1544 36771
rect 1492 36728 1544 36737
rect 9496 36728 9548 36780
rect 10692 36771 10744 36780
rect 10692 36737 10701 36771
rect 10701 36737 10735 36771
rect 10735 36737 10744 36771
rect 10692 36728 10744 36737
rect 3792 36660 3844 36712
rect 11152 36728 11204 36780
rect 12440 36839 12492 36848
rect 12440 36805 12449 36839
rect 12449 36805 12483 36839
rect 12483 36805 12492 36839
rect 12440 36796 12492 36805
rect 12900 36771 12952 36780
rect 12900 36737 12909 36771
rect 12909 36737 12943 36771
rect 12943 36737 12952 36771
rect 12900 36728 12952 36737
rect 13084 36771 13136 36780
rect 13084 36737 13093 36771
rect 13093 36737 13127 36771
rect 13127 36737 13136 36771
rect 13084 36728 13136 36737
rect 13360 36728 13412 36780
rect 6184 36524 6236 36576
rect 8300 36524 8352 36576
rect 11060 36524 11112 36576
rect 13544 36660 13596 36712
rect 13820 36771 13872 36780
rect 13820 36737 13829 36771
rect 13829 36737 13863 36771
rect 13863 36737 13872 36771
rect 13820 36728 13872 36737
rect 20076 36796 20128 36848
rect 21456 36796 21508 36848
rect 23664 36796 23716 36848
rect 13728 36592 13780 36644
rect 16028 36728 16080 36780
rect 20352 36728 20404 36780
rect 18420 36660 18472 36712
rect 20444 36660 20496 36712
rect 13636 36524 13688 36576
rect 16672 36567 16724 36576
rect 16672 36533 16681 36567
rect 16681 36533 16715 36567
rect 16715 36533 16724 36567
rect 16672 36524 16724 36533
rect 23020 36728 23072 36780
rect 24768 36771 24820 36780
rect 24768 36737 24772 36771
rect 24772 36737 24806 36771
rect 24806 36737 24820 36771
rect 24768 36728 24820 36737
rect 24860 36771 24912 36780
rect 24860 36737 24869 36771
rect 24869 36737 24903 36771
rect 24903 36737 24912 36771
rect 24860 36728 24912 36737
rect 25044 36796 25096 36848
rect 27068 36796 27120 36848
rect 27988 36796 28040 36848
rect 21364 36703 21416 36712
rect 21364 36669 21373 36703
rect 21373 36669 21407 36703
rect 21407 36669 21416 36703
rect 21364 36660 21416 36669
rect 25504 36771 25556 36780
rect 25504 36737 25513 36771
rect 25513 36737 25547 36771
rect 25547 36737 25556 36771
rect 25504 36728 25556 36737
rect 27344 36728 27396 36780
rect 30840 36907 30892 36916
rect 30840 36873 30849 36907
rect 30849 36873 30883 36907
rect 30883 36873 30892 36907
rect 30840 36864 30892 36873
rect 31024 36864 31076 36916
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 29368 36771 29420 36780
rect 29368 36737 29377 36771
rect 29377 36737 29411 36771
rect 29411 36737 29420 36771
rect 29368 36728 29420 36737
rect 26148 36660 26200 36712
rect 30104 36728 30156 36780
rect 30380 36728 30432 36780
rect 30748 36728 30800 36780
rect 31024 36771 31076 36780
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 29920 36660 29972 36712
rect 32772 36728 32824 36780
rect 31668 36703 31720 36712
rect 31668 36669 31677 36703
rect 31677 36669 31711 36703
rect 31711 36669 31720 36703
rect 31668 36660 31720 36669
rect 32404 36660 32456 36712
rect 33784 36728 33836 36780
rect 33968 36771 34020 36780
rect 33968 36737 33977 36771
rect 33977 36737 34011 36771
rect 34011 36737 34020 36771
rect 33968 36728 34020 36737
rect 34612 36796 34664 36848
rect 34336 36771 34388 36780
rect 34336 36737 34345 36771
rect 34345 36737 34379 36771
rect 34379 36737 34388 36771
rect 34336 36728 34388 36737
rect 35900 36864 35952 36916
rect 36544 36796 36596 36848
rect 37648 36796 37700 36848
rect 35992 36728 36044 36780
rect 36176 36771 36228 36780
rect 36176 36737 36185 36771
rect 36185 36737 36219 36771
rect 36219 36737 36228 36771
rect 36176 36728 36228 36737
rect 38016 36864 38068 36916
rect 38476 36864 38528 36916
rect 39856 36864 39908 36916
rect 44180 36907 44232 36916
rect 44180 36873 44189 36907
rect 44189 36873 44223 36907
rect 44223 36873 44232 36907
rect 44180 36864 44232 36873
rect 39212 36796 39264 36848
rect 39488 36796 39540 36848
rect 39672 36796 39724 36848
rect 35716 36660 35768 36712
rect 29828 36592 29880 36644
rect 32864 36592 32916 36644
rect 33416 36592 33468 36644
rect 21548 36524 21600 36576
rect 27804 36524 27856 36576
rect 29000 36567 29052 36576
rect 29000 36533 29009 36567
rect 29009 36533 29043 36567
rect 29043 36533 29052 36567
rect 29000 36524 29052 36533
rect 29736 36524 29788 36576
rect 30288 36524 30340 36576
rect 30380 36524 30432 36576
rect 33048 36524 33100 36576
rect 34520 36567 34572 36576
rect 34520 36533 34529 36567
rect 34529 36533 34563 36567
rect 34563 36533 34572 36567
rect 34520 36524 34572 36533
rect 36176 36524 36228 36576
rect 39764 36660 39816 36712
rect 41328 36771 41380 36780
rect 41328 36737 41337 36771
rect 41337 36737 41371 36771
rect 41371 36737 41380 36771
rect 41328 36728 41380 36737
rect 41420 36728 41472 36780
rect 41604 36771 41656 36780
rect 41604 36737 41613 36771
rect 41613 36737 41647 36771
rect 41647 36737 41656 36771
rect 41604 36728 41656 36737
rect 41880 36771 41932 36780
rect 41880 36737 41889 36771
rect 41889 36737 41923 36771
rect 41923 36737 41932 36771
rect 41880 36728 41932 36737
rect 42064 36728 42116 36780
rect 42800 36796 42852 36848
rect 43720 36796 43772 36848
rect 42432 36771 42484 36780
rect 42432 36737 42441 36771
rect 42441 36737 42475 36771
rect 42475 36737 42484 36771
rect 42432 36728 42484 36737
rect 42708 36703 42760 36712
rect 42708 36669 42717 36703
rect 42717 36669 42751 36703
rect 42751 36669 42760 36703
rect 42708 36660 42760 36669
rect 37280 36567 37332 36576
rect 37280 36533 37289 36567
rect 37289 36533 37323 36567
rect 37323 36533 37332 36567
rect 37280 36524 37332 36533
rect 37740 36524 37792 36576
rect 38292 36524 38344 36576
rect 40316 36567 40368 36576
rect 40316 36533 40325 36567
rect 40325 36533 40359 36567
rect 40359 36533 40368 36567
rect 40316 36524 40368 36533
rect 41328 36524 41380 36576
rect 41512 36567 41564 36576
rect 41512 36533 41521 36567
rect 41521 36533 41555 36567
rect 41555 36533 41564 36567
rect 41512 36524 41564 36533
rect 41696 36567 41748 36576
rect 41696 36533 41705 36567
rect 41705 36533 41739 36567
rect 41739 36533 41748 36567
rect 41696 36524 41748 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3792 36320 3844 36372
rect 10692 36320 10744 36372
rect 11980 36320 12032 36372
rect 7012 36184 7064 36236
rect 7748 36184 7800 36236
rect 9772 36252 9824 36304
rect 8944 36184 8996 36236
rect 11060 36184 11112 36236
rect 5356 36159 5408 36168
rect 5356 36125 5365 36159
rect 5365 36125 5399 36159
rect 5399 36125 5408 36159
rect 5356 36116 5408 36125
rect 6184 36116 6236 36168
rect 6552 36091 6604 36100
rect 6552 36057 6561 36091
rect 6561 36057 6595 36091
rect 6595 36057 6604 36091
rect 6552 36048 6604 36057
rect 4068 35980 4120 36032
rect 5080 35980 5132 36032
rect 5540 35980 5592 36032
rect 7012 36048 7064 36100
rect 8392 36048 8444 36100
rect 9588 36159 9640 36168
rect 9588 36125 9597 36159
rect 9597 36125 9631 36159
rect 9631 36125 9640 36159
rect 9588 36116 9640 36125
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 12900 36184 12952 36236
rect 12808 36159 12860 36168
rect 12808 36125 12817 36159
rect 12817 36125 12851 36159
rect 12851 36125 12860 36159
rect 12808 36116 12860 36125
rect 12992 36116 13044 36168
rect 13728 36320 13780 36372
rect 14556 36320 14608 36372
rect 16028 36363 16080 36372
rect 16028 36329 16037 36363
rect 16037 36329 16071 36363
rect 16071 36329 16080 36363
rect 16028 36320 16080 36329
rect 20444 36320 20496 36372
rect 23020 36363 23072 36372
rect 23020 36329 23029 36363
rect 23029 36329 23063 36363
rect 23063 36329 23072 36363
rect 23020 36320 23072 36329
rect 29000 36320 29052 36372
rect 31668 36320 31720 36372
rect 32864 36320 32916 36372
rect 34520 36320 34572 36372
rect 35532 36320 35584 36372
rect 13820 36295 13872 36304
rect 13820 36261 13829 36295
rect 13829 36261 13863 36295
rect 13863 36261 13872 36295
rect 13820 36252 13872 36261
rect 21548 36252 21600 36304
rect 13636 36227 13688 36236
rect 13636 36193 13645 36227
rect 13645 36193 13679 36227
rect 13679 36193 13688 36227
rect 13636 36184 13688 36193
rect 16764 36184 16816 36236
rect 16948 36184 17000 36236
rect 17776 36227 17828 36236
rect 17776 36193 17785 36227
rect 17785 36193 17819 36227
rect 17819 36193 17828 36227
rect 17776 36184 17828 36193
rect 13544 36159 13596 36168
rect 13544 36125 13553 36159
rect 13553 36125 13587 36159
rect 13587 36125 13596 36159
rect 13544 36116 13596 36125
rect 13912 36159 13964 36168
rect 13912 36125 13921 36159
rect 13921 36125 13955 36159
rect 13955 36125 13964 36159
rect 13912 36116 13964 36125
rect 18052 36159 18104 36168
rect 18052 36125 18061 36159
rect 18061 36125 18095 36159
rect 18095 36125 18104 36159
rect 18052 36116 18104 36125
rect 19432 36116 19484 36168
rect 21456 36184 21508 36236
rect 22284 36184 22336 36236
rect 27344 36252 27396 36304
rect 29184 36252 29236 36304
rect 29920 36295 29972 36304
rect 29920 36261 29929 36295
rect 29929 36261 29963 36295
rect 29963 36261 29972 36295
rect 29920 36252 29972 36261
rect 23296 36184 23348 36236
rect 25228 36184 25280 36236
rect 27804 36184 27856 36236
rect 24860 36159 24912 36168
rect 6920 35980 6972 36032
rect 7840 35980 7892 36032
rect 9312 36023 9364 36032
rect 9312 35989 9321 36023
rect 9321 35989 9355 36023
rect 9355 35989 9364 36023
rect 9312 35980 9364 35989
rect 9496 36023 9548 36032
rect 9496 35989 9505 36023
rect 9505 35989 9539 36023
rect 9539 35989 9548 36023
rect 11060 36048 11112 36100
rect 9496 35980 9548 35989
rect 9680 36023 9732 36032
rect 9680 35989 9689 36023
rect 9689 35989 9723 36023
rect 9723 35989 9732 36023
rect 9680 35980 9732 35989
rect 9772 35980 9824 36032
rect 10232 35980 10284 36032
rect 15200 36048 15252 36100
rect 12808 35980 12860 36032
rect 13084 35980 13136 36032
rect 14004 35980 14056 36032
rect 15660 36091 15712 36100
rect 15660 36057 15669 36091
rect 15669 36057 15703 36091
rect 15703 36057 15712 36091
rect 15660 36048 15712 36057
rect 17960 36048 18012 36100
rect 17868 36023 17920 36032
rect 17868 35989 17877 36023
rect 17877 35989 17911 36023
rect 17911 35989 17920 36023
rect 17868 35980 17920 35989
rect 24860 36125 24869 36159
rect 24869 36125 24903 36159
rect 24903 36125 24912 36159
rect 24860 36116 24912 36125
rect 25780 36159 25832 36168
rect 25780 36125 25789 36159
rect 25789 36125 25823 36159
rect 25823 36125 25832 36159
rect 25780 36116 25832 36125
rect 26332 36116 26384 36168
rect 27620 36048 27672 36100
rect 29092 36048 29144 36100
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 29828 36159 29880 36168
rect 29828 36125 29837 36159
rect 29837 36125 29871 36159
rect 29871 36125 29880 36159
rect 29828 36116 29880 36125
rect 30012 36159 30064 36168
rect 30012 36125 30021 36159
rect 30021 36125 30055 36159
rect 30055 36125 30064 36159
rect 30012 36116 30064 36125
rect 30564 36116 30616 36168
rect 32680 36116 32732 36168
rect 32772 36159 32824 36168
rect 32772 36125 32781 36159
rect 32781 36125 32815 36159
rect 32815 36125 32824 36159
rect 32772 36116 32824 36125
rect 33048 36159 33100 36168
rect 33048 36125 33083 36159
rect 33083 36125 33100 36159
rect 33048 36116 33100 36125
rect 20904 36023 20956 36032
rect 20904 35989 20913 36023
rect 20913 35989 20947 36023
rect 20947 35989 20956 36023
rect 20904 35980 20956 35989
rect 21456 35980 21508 36032
rect 24400 36023 24452 36032
rect 24400 35989 24409 36023
rect 24409 35989 24443 36023
rect 24443 35989 24452 36023
rect 24400 35980 24452 35989
rect 24768 36023 24820 36032
rect 24768 35989 24777 36023
rect 24777 35989 24811 36023
rect 24811 35989 24820 36023
rect 24768 35980 24820 35989
rect 29184 36023 29236 36032
rect 29184 35989 29193 36023
rect 29193 35989 29227 36023
rect 29227 35989 29236 36023
rect 29184 35980 29236 35989
rect 32864 36091 32916 36100
rect 32864 36057 32873 36091
rect 32873 36057 32907 36091
rect 32907 36057 32916 36091
rect 32864 36048 32916 36057
rect 35716 36048 35768 36100
rect 39212 36320 39264 36372
rect 40316 36320 40368 36372
rect 41696 36320 41748 36372
rect 42708 36320 42760 36372
rect 43720 36320 43772 36372
rect 38752 36184 38804 36236
rect 39856 36184 39908 36236
rect 40224 36184 40276 36236
rect 37188 36048 37240 36100
rect 34704 36023 34756 36032
rect 34704 35989 34713 36023
rect 34713 35989 34747 36023
rect 34747 35989 34756 36023
rect 34704 35980 34756 35989
rect 37740 36023 37792 36032
rect 37740 35989 37749 36023
rect 37749 35989 37783 36023
rect 37783 35989 37792 36023
rect 37740 35980 37792 35989
rect 39212 36048 39264 36100
rect 41604 35980 41656 36032
rect 42064 35980 42116 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4712 35776 4764 35828
rect 3332 35683 3384 35692
rect 3332 35649 3366 35683
rect 3366 35649 3384 35683
rect 3332 35640 3384 35649
rect 5356 35776 5408 35828
rect 5908 35819 5960 35828
rect 5908 35785 5917 35819
rect 5917 35785 5951 35819
rect 5951 35785 5960 35819
rect 5908 35776 5960 35785
rect 6000 35776 6052 35828
rect 6276 35776 6328 35828
rect 9404 35776 9456 35828
rect 2964 35436 3016 35488
rect 4620 35436 4672 35488
rect 9496 35708 9548 35760
rect 9772 35708 9824 35760
rect 7012 35640 7064 35692
rect 7104 35683 7156 35692
rect 7104 35649 7113 35683
rect 7113 35649 7147 35683
rect 7147 35649 7156 35683
rect 7104 35640 7156 35649
rect 7840 35640 7892 35692
rect 6000 35615 6052 35624
rect 6000 35581 6009 35615
rect 6009 35581 6043 35615
rect 6043 35581 6052 35615
rect 6000 35572 6052 35581
rect 6920 35615 6972 35624
rect 6920 35581 6929 35615
rect 6929 35581 6963 35615
rect 6963 35581 6972 35615
rect 6920 35572 6972 35581
rect 8300 35640 8352 35692
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 12900 35776 12952 35828
rect 13820 35776 13872 35828
rect 13912 35819 13964 35828
rect 13912 35785 13921 35819
rect 13921 35785 13955 35819
rect 13955 35785 13964 35819
rect 13912 35776 13964 35785
rect 16672 35776 16724 35828
rect 14004 35708 14056 35760
rect 8392 35572 8444 35624
rect 9680 35572 9732 35624
rect 11060 35572 11112 35624
rect 14556 35640 14608 35692
rect 14740 35683 14792 35692
rect 14740 35649 14749 35683
rect 14749 35649 14783 35683
rect 14783 35649 14792 35683
rect 14740 35640 14792 35649
rect 17868 35776 17920 35828
rect 19432 35776 19484 35828
rect 20352 35776 20404 35828
rect 20444 35819 20496 35828
rect 20444 35785 20453 35819
rect 20453 35785 20487 35819
rect 20487 35785 20496 35819
rect 20444 35776 20496 35785
rect 17960 35708 18012 35760
rect 24400 35776 24452 35828
rect 25780 35776 25832 35828
rect 30932 35776 30984 35828
rect 32404 35776 32456 35828
rect 32772 35776 32824 35828
rect 32864 35776 32916 35828
rect 33968 35776 34020 35828
rect 34060 35776 34112 35828
rect 34612 35776 34664 35828
rect 35716 35819 35768 35828
rect 35716 35785 35725 35819
rect 35725 35785 35759 35819
rect 35759 35785 35768 35819
rect 35716 35776 35768 35785
rect 37924 35819 37976 35828
rect 37924 35785 37933 35819
rect 37933 35785 37967 35819
rect 37967 35785 37976 35819
rect 37924 35776 37976 35785
rect 38384 35776 38436 35828
rect 11980 35572 12032 35624
rect 12532 35572 12584 35624
rect 15660 35572 15712 35624
rect 16948 35572 17000 35624
rect 20904 35640 20956 35692
rect 27620 35640 27672 35692
rect 29552 35640 29604 35692
rect 30012 35640 30064 35692
rect 37188 35708 37240 35760
rect 17776 35572 17828 35624
rect 5816 35436 5868 35488
rect 22376 35615 22428 35624
rect 22376 35581 22385 35615
rect 22385 35581 22419 35615
rect 22419 35581 22428 35615
rect 22376 35572 22428 35581
rect 23296 35572 23348 35624
rect 6920 35436 6972 35488
rect 9588 35436 9640 35488
rect 10692 35479 10744 35488
rect 10692 35445 10701 35479
rect 10701 35445 10735 35479
rect 10735 35445 10744 35479
rect 10692 35436 10744 35445
rect 19156 35479 19208 35488
rect 19156 35445 19165 35479
rect 19165 35445 19199 35479
rect 19199 35445 19208 35479
rect 19156 35436 19208 35445
rect 21548 35436 21600 35488
rect 27620 35504 27672 35556
rect 29920 35572 29972 35624
rect 30288 35615 30340 35624
rect 30288 35581 30297 35615
rect 30297 35581 30331 35615
rect 30331 35581 30340 35615
rect 30288 35572 30340 35581
rect 33416 35640 33468 35692
rect 34152 35683 34204 35692
rect 34152 35649 34161 35683
rect 34161 35649 34195 35683
rect 34195 35649 34204 35683
rect 34152 35640 34204 35649
rect 34704 35640 34756 35692
rect 33600 35615 33652 35624
rect 33600 35581 33609 35615
rect 33609 35581 33643 35615
rect 33643 35581 33652 35615
rect 33600 35572 33652 35581
rect 37740 35572 37792 35624
rect 38476 35572 38528 35624
rect 41512 35615 41564 35624
rect 41512 35581 41521 35615
rect 41521 35581 41555 35615
rect 41555 35581 41564 35615
rect 41512 35572 41564 35581
rect 29828 35504 29880 35556
rect 30104 35504 30156 35556
rect 33508 35504 33560 35556
rect 25228 35436 25280 35488
rect 25872 35436 25924 35488
rect 40960 35479 41012 35488
rect 40960 35445 40969 35479
rect 40969 35445 41003 35479
rect 41003 35445 41012 35479
rect 40960 35436 41012 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3332 35232 3384 35284
rect 2964 35028 3016 35080
rect 4620 35232 4672 35284
rect 4804 35232 4856 35284
rect 6552 35232 6604 35284
rect 6920 35232 6972 35284
rect 9312 35232 9364 35284
rect 9864 35232 9916 35284
rect 10692 35232 10744 35284
rect 18052 35232 18104 35284
rect 19156 35232 19208 35284
rect 22376 35232 22428 35284
rect 26148 35232 26200 35284
rect 4620 35096 4672 35148
rect 4252 35071 4304 35080
rect 4252 35037 4261 35071
rect 4261 35037 4295 35071
rect 4295 35037 4304 35071
rect 4252 35028 4304 35037
rect 6184 35096 6236 35148
rect 12440 35164 12492 35216
rect 13176 35164 13228 35216
rect 2136 34960 2188 35012
rect 5080 34960 5132 35012
rect 5540 34960 5592 35012
rect 3056 34935 3108 34944
rect 3056 34901 3065 34935
rect 3065 34901 3099 34935
rect 3099 34901 3108 34935
rect 3056 34892 3108 34901
rect 5356 34892 5408 34944
rect 5816 34892 5868 34944
rect 6920 34892 6972 34944
rect 9496 34960 9548 35012
rect 18144 35096 18196 35148
rect 18420 35139 18472 35148
rect 18420 35105 18429 35139
rect 18429 35105 18463 35139
rect 18463 35105 18472 35139
rect 18420 35096 18472 35105
rect 18236 35071 18288 35080
rect 18236 35037 18245 35071
rect 18245 35037 18279 35071
rect 18279 35037 18288 35071
rect 30288 35275 30340 35284
rect 30288 35241 30297 35275
rect 30297 35241 30331 35275
rect 30331 35241 30340 35275
rect 30288 35232 30340 35241
rect 33600 35232 33652 35284
rect 34152 35232 34204 35284
rect 35716 35232 35768 35284
rect 22468 35139 22520 35148
rect 22468 35105 22477 35139
rect 22477 35105 22511 35139
rect 22511 35105 22520 35139
rect 22468 35096 22520 35105
rect 23296 35096 23348 35148
rect 25872 35096 25924 35148
rect 27804 35096 27856 35148
rect 18236 35028 18288 35037
rect 19432 35028 19484 35080
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 24032 35071 24084 35080
rect 24032 35037 24041 35071
rect 24041 35037 24075 35071
rect 24075 35037 24084 35071
rect 24032 35028 24084 35037
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30104 35071 30156 35080
rect 30104 35037 30113 35071
rect 30113 35037 30147 35071
rect 30147 35037 30156 35071
rect 30104 35028 30156 35037
rect 22100 34960 22152 35012
rect 27896 35003 27948 35012
rect 27896 34969 27905 35003
rect 27905 34969 27939 35003
rect 27939 34969 27948 35003
rect 27896 34960 27948 34969
rect 12256 34892 12308 34944
rect 19984 34892 20036 34944
rect 24584 34892 24636 34944
rect 26056 34892 26108 34944
rect 26516 34892 26568 34944
rect 26608 34892 26660 34944
rect 28080 34892 28132 34944
rect 30288 34892 30340 34944
rect 33140 35071 33192 35080
rect 33140 35037 33149 35071
rect 33149 35037 33183 35071
rect 33183 35037 33192 35071
rect 33140 35028 33192 35037
rect 33324 35071 33376 35080
rect 33324 35037 33333 35071
rect 33333 35037 33367 35071
rect 33367 35037 33376 35071
rect 33324 35028 33376 35037
rect 33508 35028 33560 35080
rect 40224 35096 40276 35148
rect 40960 35139 41012 35148
rect 40960 35105 40969 35139
rect 40969 35105 41003 35139
rect 41003 35105 41012 35139
rect 40960 35096 41012 35105
rect 37188 35071 37240 35080
rect 37188 35037 37197 35071
rect 37197 35037 37231 35071
rect 37231 35037 37240 35071
rect 37188 35028 37240 35037
rect 38660 35071 38712 35080
rect 38660 35037 38669 35071
rect 38669 35037 38703 35071
rect 38703 35037 38712 35071
rect 38660 35028 38712 35037
rect 40040 35028 40092 35080
rect 36176 34892 36228 34944
rect 36268 34892 36320 34944
rect 39304 34960 39356 35012
rect 38016 34892 38068 34944
rect 38752 34892 38804 34944
rect 41972 34892 42024 34944
rect 44088 34892 44140 34944
rect 45284 34892 45336 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2136 34731 2188 34740
rect 2136 34697 2145 34731
rect 2145 34697 2179 34731
rect 2179 34697 2188 34731
rect 2136 34688 2188 34697
rect 4252 34688 4304 34740
rect 13268 34688 13320 34740
rect 3792 34552 3844 34604
rect 5172 34552 5224 34604
rect 7564 34595 7616 34604
rect 7564 34561 7573 34595
rect 7573 34561 7607 34595
rect 7607 34561 7616 34595
rect 7564 34552 7616 34561
rect 8576 34595 8628 34604
rect 8576 34561 8585 34595
rect 8585 34561 8619 34595
rect 8619 34561 8628 34595
rect 8576 34552 8628 34561
rect 10232 34552 10284 34604
rect 13728 34620 13780 34672
rect 13268 34552 13320 34604
rect 13360 34552 13412 34604
rect 14556 34688 14608 34740
rect 16856 34688 16908 34740
rect 18052 34688 18104 34740
rect 18236 34688 18288 34740
rect 19432 34688 19484 34740
rect 19984 34688 20036 34740
rect 20444 34688 20496 34740
rect 21548 34688 21600 34740
rect 2872 34416 2924 34468
rect 8852 34527 8904 34536
rect 8852 34493 8861 34527
rect 8861 34493 8895 34527
rect 8895 34493 8904 34527
rect 8852 34484 8904 34493
rect 14188 34552 14240 34604
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 20260 34552 20312 34561
rect 23388 34688 23440 34740
rect 24032 34688 24084 34740
rect 24768 34731 24820 34740
rect 24768 34697 24777 34731
rect 24777 34697 24811 34731
rect 24811 34697 24820 34731
rect 24768 34688 24820 34697
rect 27896 34688 27948 34740
rect 33140 34731 33192 34740
rect 33140 34697 33149 34731
rect 33149 34697 33183 34731
rect 33183 34697 33192 34731
rect 33140 34688 33192 34697
rect 33324 34688 33376 34740
rect 36268 34688 36320 34740
rect 26424 34663 26476 34672
rect 26424 34629 26433 34663
rect 26433 34629 26467 34663
rect 26467 34629 26476 34663
rect 26424 34620 26476 34629
rect 22652 34552 22704 34604
rect 24676 34595 24728 34604
rect 24676 34561 24685 34595
rect 24685 34561 24719 34595
rect 24719 34561 24728 34595
rect 24676 34552 24728 34561
rect 26240 34595 26292 34604
rect 26240 34561 26249 34595
rect 26249 34561 26283 34595
rect 26283 34561 26292 34595
rect 26240 34552 26292 34561
rect 26516 34595 26568 34604
rect 26516 34561 26525 34595
rect 26525 34561 26559 34595
rect 26559 34561 26568 34595
rect 26516 34552 26568 34561
rect 28540 34620 28592 34672
rect 31668 34620 31720 34672
rect 17868 34527 17920 34536
rect 17868 34493 17877 34527
rect 17877 34493 17911 34527
rect 17911 34493 17920 34527
rect 17868 34484 17920 34493
rect 18420 34484 18472 34536
rect 5724 34416 5776 34468
rect 12440 34416 12492 34468
rect 20996 34484 21048 34536
rect 4804 34391 4856 34400
rect 4804 34357 4813 34391
rect 4813 34357 4847 34391
rect 4847 34357 4856 34391
rect 4804 34348 4856 34357
rect 7380 34391 7432 34400
rect 7380 34357 7389 34391
rect 7389 34357 7423 34391
rect 7423 34357 7432 34391
rect 7380 34348 7432 34357
rect 8760 34391 8812 34400
rect 8760 34357 8769 34391
rect 8769 34357 8803 34391
rect 8803 34357 8812 34391
rect 8760 34348 8812 34357
rect 9496 34391 9548 34400
rect 9496 34357 9505 34391
rect 9505 34357 9539 34391
rect 9539 34357 9548 34391
rect 9496 34348 9548 34357
rect 9956 34348 10008 34400
rect 12900 34391 12952 34400
rect 12900 34357 12909 34391
rect 12909 34357 12943 34391
rect 12943 34357 12952 34391
rect 12900 34348 12952 34357
rect 13820 34348 13872 34400
rect 14280 34348 14332 34400
rect 15752 34348 15804 34400
rect 16120 34348 16172 34400
rect 17040 34348 17092 34400
rect 19616 34391 19668 34400
rect 19616 34357 19625 34391
rect 19625 34357 19659 34391
rect 19659 34357 19668 34391
rect 19616 34348 19668 34357
rect 21088 34348 21140 34400
rect 22008 34348 22060 34400
rect 24492 34484 24544 34536
rect 27620 34552 27672 34604
rect 28172 34552 28224 34604
rect 32588 34620 32640 34672
rect 33232 34552 33284 34604
rect 33600 34595 33652 34604
rect 31484 34484 31536 34536
rect 33600 34561 33609 34595
rect 33609 34561 33643 34595
rect 33643 34561 33652 34595
rect 33600 34552 33652 34561
rect 34060 34552 34112 34604
rect 38660 34688 38712 34740
rect 39764 34688 39816 34740
rect 37372 34620 37424 34672
rect 36544 34552 36596 34604
rect 34520 34484 34572 34536
rect 36820 34595 36872 34604
rect 36820 34561 36829 34595
rect 36829 34561 36863 34595
rect 36863 34561 36872 34595
rect 36820 34552 36872 34561
rect 37924 34552 37976 34604
rect 38292 34552 38344 34604
rect 38476 34595 38528 34604
rect 38476 34561 38485 34595
rect 38485 34561 38519 34595
rect 38519 34561 38528 34595
rect 38476 34552 38528 34561
rect 37096 34484 37148 34536
rect 38844 34620 38896 34672
rect 40592 34620 40644 34672
rect 41512 34688 41564 34740
rect 41696 34688 41748 34740
rect 38752 34595 38804 34604
rect 38752 34561 38761 34595
rect 38761 34561 38795 34595
rect 38795 34561 38804 34595
rect 38752 34552 38804 34561
rect 37004 34416 37056 34468
rect 38384 34416 38436 34468
rect 39120 34527 39172 34536
rect 39120 34493 39129 34527
rect 39129 34493 39163 34527
rect 39163 34493 39172 34527
rect 39120 34484 39172 34493
rect 39580 34484 39632 34536
rect 41604 34595 41656 34604
rect 41604 34561 41613 34595
rect 41613 34561 41647 34595
rect 41647 34561 41656 34595
rect 41604 34552 41656 34561
rect 43536 34620 43588 34672
rect 41972 34595 42024 34604
rect 41972 34561 41981 34595
rect 41981 34561 42015 34595
rect 42015 34561 42024 34595
rect 41972 34552 42024 34561
rect 42524 34595 42576 34604
rect 42524 34561 42533 34595
rect 42533 34561 42567 34595
rect 42567 34561 42576 34595
rect 42524 34552 42576 34561
rect 42800 34527 42852 34536
rect 42800 34493 42809 34527
rect 42809 34493 42843 34527
rect 42843 34493 42852 34527
rect 42800 34484 42852 34493
rect 43076 34484 43128 34536
rect 32588 34348 32640 34400
rect 33324 34348 33376 34400
rect 38108 34391 38160 34400
rect 38108 34357 38117 34391
rect 38117 34357 38151 34391
rect 38151 34357 38160 34391
rect 38108 34348 38160 34357
rect 40408 34348 40460 34400
rect 40684 34391 40736 34400
rect 40684 34357 40693 34391
rect 40693 34357 40727 34391
rect 40727 34357 40736 34391
rect 40684 34348 40736 34357
rect 40776 34348 40828 34400
rect 43536 34348 43588 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5172 34187 5224 34196
rect 5172 34153 5181 34187
rect 5181 34153 5215 34187
rect 5215 34153 5224 34187
rect 5172 34144 5224 34153
rect 8852 34144 8904 34196
rect 8944 34051 8996 34060
rect 8944 34017 8953 34051
rect 8953 34017 8987 34051
rect 8987 34017 8996 34051
rect 8944 34008 8996 34017
rect 12440 34051 12492 34060
rect 12440 34017 12449 34051
rect 12449 34017 12483 34051
rect 12483 34017 12492 34051
rect 12440 34008 12492 34017
rect 13728 34144 13780 34196
rect 14556 34144 14608 34196
rect 14648 34187 14700 34196
rect 14648 34153 14657 34187
rect 14657 34153 14691 34187
rect 14691 34153 14700 34187
rect 14648 34144 14700 34153
rect 15660 34144 15712 34196
rect 15752 34187 15804 34196
rect 15752 34153 15761 34187
rect 15761 34153 15795 34187
rect 15795 34153 15804 34187
rect 15752 34144 15804 34153
rect 16028 34144 16080 34196
rect 16672 34144 16724 34196
rect 20260 34144 20312 34196
rect 22008 34144 22060 34196
rect 3240 33983 3292 33992
rect 3240 33949 3249 33983
rect 3249 33949 3283 33983
rect 3283 33949 3292 33983
rect 3240 33940 3292 33949
rect 5172 33940 5224 33992
rect 5724 33983 5776 33992
rect 5724 33949 5733 33983
rect 5733 33949 5767 33983
rect 5767 33949 5776 33983
rect 5724 33940 5776 33949
rect 7104 33983 7156 33992
rect 7104 33949 7113 33983
rect 7113 33949 7147 33983
rect 7147 33949 7156 33983
rect 7104 33940 7156 33949
rect 7380 33983 7432 33992
rect 7380 33949 7414 33983
rect 7414 33949 7432 33983
rect 7380 33940 7432 33949
rect 8760 33940 8812 33992
rect 3884 33872 3936 33924
rect 4160 33872 4212 33924
rect 9956 33872 10008 33924
rect 2412 33804 2464 33856
rect 6092 33804 6144 33856
rect 9128 33804 9180 33856
rect 10876 33915 10928 33924
rect 10876 33881 10885 33915
rect 10885 33881 10919 33915
rect 10919 33881 10928 33915
rect 10876 33872 10928 33881
rect 12900 33983 12952 33992
rect 12900 33949 12942 33983
rect 12942 33949 12952 33983
rect 12900 33940 12952 33949
rect 13360 33940 13412 33992
rect 13544 33940 13596 33992
rect 13728 33983 13780 33992
rect 13728 33949 13737 33983
rect 13737 33949 13771 33983
rect 13771 33949 13780 33983
rect 13728 33940 13780 33949
rect 14372 33940 14424 33992
rect 14464 33940 14516 33992
rect 16028 33983 16080 33992
rect 16028 33949 16037 33983
rect 16037 33949 16071 33983
rect 16071 33949 16080 33983
rect 16028 33940 16080 33949
rect 16120 33983 16172 33992
rect 16120 33949 16129 33983
rect 16129 33949 16163 33983
rect 16163 33949 16172 33983
rect 16120 33940 16172 33949
rect 16212 33940 16264 33992
rect 17132 33983 17184 33992
rect 17132 33949 17141 33983
rect 17141 33949 17175 33983
rect 17175 33949 17184 33983
rect 17132 33940 17184 33949
rect 17316 33983 17368 33992
rect 17316 33949 17325 33983
rect 17325 33949 17359 33983
rect 17359 33949 17368 33983
rect 17316 33940 17368 33949
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 22284 34076 22336 34128
rect 22100 34051 22152 34060
rect 22100 34017 22109 34051
rect 22109 34017 22143 34051
rect 22143 34017 22152 34051
rect 22100 34008 22152 34017
rect 29368 34144 29420 34196
rect 33048 34144 33100 34196
rect 33324 34144 33376 34196
rect 33692 34144 33744 34196
rect 33876 34144 33928 34196
rect 34060 34187 34112 34196
rect 34060 34153 34069 34187
rect 34069 34153 34103 34187
rect 34103 34153 34112 34187
rect 34060 34144 34112 34153
rect 37004 34144 37056 34196
rect 40040 34144 40092 34196
rect 42524 34144 42576 34196
rect 42800 34144 42852 34196
rect 10968 33804 11020 33856
rect 11612 33847 11664 33856
rect 11612 33813 11621 33847
rect 11621 33813 11655 33847
rect 11655 33813 11664 33847
rect 11612 33804 11664 33813
rect 11888 33804 11940 33856
rect 12808 33847 12860 33856
rect 12808 33813 12817 33847
rect 12817 33813 12851 33847
rect 12851 33813 12860 33847
rect 12808 33804 12860 33813
rect 13820 33872 13872 33924
rect 15752 33872 15804 33924
rect 17224 33872 17276 33924
rect 15016 33804 15068 33856
rect 16856 33804 16908 33856
rect 17592 33915 17644 33924
rect 17592 33881 17601 33915
rect 17601 33881 17635 33915
rect 17635 33881 17644 33915
rect 17592 33872 17644 33881
rect 17684 33872 17736 33924
rect 18144 33847 18196 33856
rect 18144 33813 18153 33847
rect 18153 33813 18187 33847
rect 18187 33813 18196 33847
rect 18144 33804 18196 33813
rect 19616 33872 19668 33924
rect 23480 33940 23532 33992
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 27988 33940 28040 33992
rect 28724 33940 28776 33992
rect 33048 34051 33100 34060
rect 33048 34017 33057 34051
rect 33057 34017 33091 34051
rect 33091 34017 33100 34051
rect 33048 34008 33100 34017
rect 33232 34008 33284 34060
rect 33140 33940 33192 33992
rect 33416 33983 33468 33992
rect 33416 33949 33425 33983
rect 33425 33949 33459 33983
rect 33459 33949 33468 33983
rect 33416 33940 33468 33949
rect 33600 33983 33652 33992
rect 33600 33949 33609 33983
rect 33609 33949 33643 33983
rect 33643 33949 33652 33983
rect 33600 33940 33652 33949
rect 33968 33983 34020 33992
rect 33968 33949 33977 33983
rect 33977 33949 34011 33983
rect 34011 33949 34020 33983
rect 33968 33940 34020 33949
rect 37280 34008 37332 34060
rect 37648 34051 37700 34060
rect 37648 34017 37657 34051
rect 37657 34017 37691 34051
rect 37691 34017 37700 34051
rect 37648 34008 37700 34017
rect 38384 34008 38436 34060
rect 40776 34008 40828 34060
rect 41328 34008 41380 34060
rect 21180 33915 21232 33924
rect 21180 33881 21189 33915
rect 21189 33881 21223 33915
rect 21223 33881 21232 33915
rect 21180 33872 21232 33881
rect 32864 33872 32916 33924
rect 21640 33847 21692 33856
rect 21640 33813 21649 33847
rect 21649 33813 21683 33847
rect 21683 33813 21692 33847
rect 21640 33804 21692 33813
rect 22008 33847 22060 33856
rect 22008 33813 22017 33847
rect 22017 33813 22051 33847
rect 22051 33813 22060 33847
rect 22008 33804 22060 33813
rect 25228 33804 25280 33856
rect 27528 33804 27580 33856
rect 33140 33804 33192 33856
rect 33416 33847 33468 33856
rect 33416 33813 33425 33847
rect 33425 33813 33459 33847
rect 33459 33813 33468 33847
rect 33416 33804 33468 33813
rect 35900 33804 35952 33856
rect 36636 33804 36688 33856
rect 37004 33940 37056 33992
rect 39028 33940 39080 33992
rect 40408 33940 40460 33992
rect 38016 33872 38068 33924
rect 39948 33872 40000 33924
rect 41972 33872 42024 33924
rect 42984 33915 43036 33924
rect 42984 33881 42993 33915
rect 42993 33881 43027 33915
rect 43027 33881 43036 33915
rect 42984 33872 43036 33881
rect 43076 33872 43128 33924
rect 43444 33872 43496 33924
rect 37280 33804 37332 33856
rect 38292 33804 38344 33856
rect 38844 33804 38896 33856
rect 39580 33804 39632 33856
rect 43628 33804 43680 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 3884 33643 3936 33652
rect 3884 33609 3893 33643
rect 3893 33609 3927 33643
rect 3927 33609 3936 33643
rect 3884 33600 3936 33609
rect 3516 33507 3568 33516
rect 3516 33473 3525 33507
rect 3525 33473 3559 33507
rect 3559 33473 3568 33507
rect 3516 33464 3568 33473
rect 4804 33600 4856 33652
rect 5080 33643 5132 33652
rect 5080 33609 5089 33643
rect 5089 33609 5123 33643
rect 5123 33609 5132 33643
rect 5080 33600 5132 33609
rect 5724 33600 5776 33652
rect 7564 33643 7616 33652
rect 7564 33609 7573 33643
rect 7573 33609 7607 33643
rect 7607 33609 7616 33643
rect 7564 33600 7616 33609
rect 8576 33600 8628 33652
rect 9128 33643 9180 33652
rect 9128 33609 9137 33643
rect 9137 33609 9171 33643
rect 9171 33609 9180 33643
rect 9128 33600 9180 33609
rect 4160 33464 4212 33516
rect 2504 33260 2556 33312
rect 2596 33260 2648 33312
rect 4620 33439 4672 33448
rect 4620 33405 4629 33439
rect 4629 33405 4663 33439
rect 4663 33405 4672 33439
rect 4620 33396 4672 33405
rect 5632 33532 5684 33584
rect 6092 33464 6144 33516
rect 6920 33464 6972 33516
rect 9496 33600 9548 33652
rect 10876 33600 10928 33652
rect 11244 33600 11296 33652
rect 12164 33643 12216 33652
rect 12164 33609 12173 33643
rect 12173 33609 12207 33643
rect 12207 33609 12216 33643
rect 12164 33600 12216 33609
rect 12808 33600 12860 33652
rect 5540 33328 5592 33380
rect 6368 33439 6420 33448
rect 6368 33405 6377 33439
rect 6377 33405 6411 33439
rect 6411 33405 6420 33439
rect 6368 33396 6420 33405
rect 8024 33439 8076 33448
rect 8024 33405 8033 33439
rect 8033 33405 8067 33439
rect 8067 33405 8076 33439
rect 8024 33396 8076 33405
rect 11060 33507 11112 33516
rect 11060 33473 11069 33507
rect 11069 33473 11103 33507
rect 11103 33473 11112 33507
rect 11060 33464 11112 33473
rect 11612 33464 11664 33516
rect 11704 33507 11756 33516
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 11888 33464 11940 33516
rect 14556 33600 14608 33652
rect 14464 33464 14516 33516
rect 14648 33575 14700 33584
rect 14648 33541 14657 33575
rect 14657 33541 14691 33575
rect 14691 33541 14700 33575
rect 14648 33532 14700 33541
rect 16028 33600 16080 33652
rect 16856 33600 16908 33652
rect 17224 33600 17276 33652
rect 17316 33575 17368 33584
rect 17316 33541 17325 33575
rect 17325 33541 17359 33575
rect 17359 33541 17368 33575
rect 17316 33532 17368 33541
rect 14924 33464 14976 33516
rect 9404 33439 9456 33448
rect 9404 33405 9413 33439
rect 9413 33405 9447 33439
rect 9447 33405 9456 33439
rect 9404 33396 9456 33405
rect 10600 33396 10652 33448
rect 10968 33396 11020 33448
rect 11244 33396 11296 33448
rect 6828 33328 6880 33380
rect 5632 33303 5684 33312
rect 5632 33269 5641 33303
rect 5641 33269 5675 33303
rect 5675 33269 5684 33303
rect 5632 33260 5684 33269
rect 9588 33260 9640 33312
rect 11980 33303 12032 33312
rect 11980 33269 11989 33303
rect 11989 33269 12023 33303
rect 12023 33269 12032 33303
rect 11980 33260 12032 33269
rect 14280 33371 14332 33380
rect 14280 33337 14289 33371
rect 14289 33337 14323 33371
rect 14323 33337 14332 33371
rect 14280 33328 14332 33337
rect 14096 33260 14148 33312
rect 15200 33439 15252 33448
rect 15200 33405 15209 33439
rect 15209 33405 15243 33439
rect 15243 33405 15252 33439
rect 15200 33396 15252 33405
rect 15292 33439 15344 33448
rect 15292 33405 15301 33439
rect 15301 33405 15335 33439
rect 15335 33405 15344 33439
rect 15292 33396 15344 33405
rect 16212 33464 16264 33516
rect 16396 33507 16448 33516
rect 16396 33473 16405 33507
rect 16405 33473 16439 33507
rect 16439 33473 16448 33507
rect 16396 33464 16448 33473
rect 16488 33464 16540 33516
rect 16304 33396 16356 33448
rect 17776 33507 17828 33516
rect 17776 33473 17785 33507
rect 17785 33473 17819 33507
rect 17819 33473 17828 33507
rect 17776 33464 17828 33473
rect 17684 33328 17736 33380
rect 15844 33303 15896 33312
rect 15844 33269 15853 33303
rect 15853 33269 15887 33303
rect 15887 33269 15896 33303
rect 15844 33260 15896 33269
rect 15936 33260 15988 33312
rect 18052 33600 18104 33652
rect 20076 33600 20128 33652
rect 21640 33600 21692 33652
rect 24400 33643 24452 33652
rect 24400 33609 24409 33643
rect 24409 33609 24443 33643
rect 24443 33609 24452 33643
rect 24400 33600 24452 33609
rect 25044 33600 25096 33652
rect 25228 33600 25280 33652
rect 21548 33532 21600 33584
rect 18144 33464 18196 33516
rect 19156 33396 19208 33448
rect 20260 33464 20312 33516
rect 23940 33532 23992 33584
rect 27528 33600 27580 33652
rect 24768 33464 24820 33516
rect 26332 33464 26384 33516
rect 27712 33464 27764 33516
rect 24676 33396 24728 33448
rect 23940 33328 23992 33380
rect 29460 33396 29512 33448
rect 18788 33303 18840 33312
rect 18788 33269 18797 33303
rect 18797 33269 18831 33303
rect 18831 33269 18840 33303
rect 18788 33260 18840 33269
rect 18880 33260 18932 33312
rect 21272 33303 21324 33312
rect 21272 33269 21281 33303
rect 21281 33269 21315 33303
rect 21315 33269 21324 33303
rect 21272 33260 21324 33269
rect 29368 33260 29420 33312
rect 29552 33260 29604 33312
rect 30748 33396 30800 33448
rect 33968 33600 34020 33652
rect 35532 33600 35584 33652
rect 37188 33532 37240 33584
rect 35900 33464 35952 33516
rect 36820 33464 36872 33516
rect 37648 33532 37700 33584
rect 39028 33532 39080 33584
rect 38844 33464 38896 33516
rect 40684 33600 40736 33652
rect 42892 33643 42944 33652
rect 42892 33609 42901 33643
rect 42901 33609 42935 33643
rect 42935 33609 42944 33643
rect 42892 33600 42944 33609
rect 42984 33600 43036 33652
rect 43628 33600 43680 33652
rect 31760 33439 31812 33448
rect 31760 33405 31769 33439
rect 31769 33405 31803 33439
rect 31803 33405 31812 33439
rect 31760 33396 31812 33405
rect 34796 33396 34848 33448
rect 35992 33396 36044 33448
rect 38108 33396 38160 33448
rect 38292 33396 38344 33448
rect 39488 33507 39540 33516
rect 39488 33473 39497 33507
rect 39497 33473 39531 33507
rect 39531 33473 39540 33507
rect 39488 33464 39540 33473
rect 34060 33328 34112 33380
rect 40224 33507 40276 33516
rect 40224 33473 40233 33507
rect 40233 33473 40267 33507
rect 40267 33473 40276 33507
rect 40224 33464 40276 33473
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 36544 33260 36596 33312
rect 37004 33260 37056 33312
rect 39028 33303 39080 33312
rect 39028 33269 39037 33303
rect 39037 33269 39071 33303
rect 39071 33269 39080 33303
rect 39028 33260 39080 33269
rect 39212 33260 39264 33312
rect 40500 33439 40552 33448
rect 40500 33405 40509 33439
rect 40509 33405 40543 33439
rect 40543 33405 40552 33439
rect 41328 33464 41380 33516
rect 42064 33507 42116 33516
rect 42064 33473 42073 33507
rect 42073 33473 42107 33507
rect 42107 33473 42116 33507
rect 42064 33464 42116 33473
rect 43168 33532 43220 33584
rect 40500 33396 40552 33405
rect 42892 33396 42944 33448
rect 44272 33396 44324 33448
rect 44088 33371 44140 33380
rect 44088 33337 44097 33371
rect 44097 33337 44131 33371
rect 44131 33337 44140 33371
rect 44088 33328 44140 33337
rect 39856 33303 39908 33312
rect 39856 33269 39865 33303
rect 39865 33269 39899 33303
rect 39899 33269 39908 33303
rect 39856 33260 39908 33269
rect 41512 33303 41564 33312
rect 41512 33269 41521 33303
rect 41521 33269 41555 33303
rect 41555 33269 41564 33303
rect 41512 33260 41564 33269
rect 43904 33303 43956 33312
rect 43904 33269 43913 33303
rect 43913 33269 43947 33303
rect 43947 33269 43956 33303
rect 43904 33260 43956 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3516 33056 3568 33108
rect 2504 32963 2556 32972
rect 2504 32929 2513 32963
rect 2513 32929 2547 32963
rect 2547 32929 2556 32963
rect 2504 32920 2556 32929
rect 2872 32920 2924 32972
rect 4620 33056 4672 33108
rect 6368 33056 6420 33108
rect 7104 33056 7156 33108
rect 8116 33099 8168 33108
rect 8116 33065 8125 33099
rect 8125 33065 8159 33099
rect 8159 33065 8168 33099
rect 8116 33056 8168 33065
rect 2412 32895 2464 32904
rect 2412 32861 2421 32895
rect 2421 32861 2455 32895
rect 2455 32861 2464 32895
rect 2412 32852 2464 32861
rect 3700 32852 3752 32904
rect 5172 32852 5224 32904
rect 5632 32852 5684 32904
rect 6092 32895 6144 32904
rect 6092 32861 6101 32895
rect 6101 32861 6135 32895
rect 6135 32861 6144 32895
rect 6092 32852 6144 32861
rect 9220 32988 9272 33040
rect 11060 32988 11112 33040
rect 11888 33056 11940 33108
rect 14280 33056 14332 33108
rect 14648 33056 14700 33108
rect 12900 32988 12952 33040
rect 7288 32852 7340 32904
rect 8024 32852 8076 32904
rect 10048 32852 10100 32904
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 7196 32784 7248 32836
rect 11704 32963 11756 32972
rect 11704 32929 11713 32963
rect 11713 32929 11747 32963
rect 11747 32929 11756 32963
rect 11704 32920 11756 32929
rect 11612 32895 11664 32904
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 13544 32920 13596 32972
rect 14096 32920 14148 32972
rect 12992 32895 13044 32904
rect 12992 32861 13001 32895
rect 13001 32861 13035 32895
rect 13035 32861 13044 32895
rect 12992 32852 13044 32861
rect 13728 32852 13780 32904
rect 14464 32852 14516 32904
rect 15200 32988 15252 33040
rect 15108 32963 15160 32972
rect 15108 32929 15117 32963
rect 15117 32929 15151 32963
rect 15151 32929 15160 32963
rect 15108 32920 15160 32929
rect 16488 33056 16540 33108
rect 16764 33099 16816 33108
rect 16764 33065 16773 33099
rect 16773 33065 16807 33099
rect 16807 33065 16816 33099
rect 16764 33056 16816 33065
rect 17684 33056 17736 33108
rect 18420 33099 18472 33108
rect 18420 33065 18429 33099
rect 18429 33065 18463 33099
rect 18463 33065 18472 33099
rect 18420 33056 18472 33065
rect 24584 33056 24636 33108
rect 24768 33056 24820 33108
rect 27712 33056 27764 33108
rect 28908 33056 28960 33108
rect 30288 33056 30340 33108
rect 30748 33056 30800 33108
rect 31944 33056 31996 33108
rect 32680 33056 32732 33108
rect 34796 33056 34848 33108
rect 35992 33056 36044 33108
rect 36912 33056 36964 33108
rect 37096 33099 37148 33108
rect 37096 33065 37105 33099
rect 37105 33065 37139 33099
rect 37139 33065 37148 33099
rect 37096 33056 37148 33065
rect 15200 32895 15252 32904
rect 15200 32861 15209 32895
rect 15209 32861 15243 32895
rect 15243 32861 15252 32895
rect 15200 32852 15252 32861
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 5724 32716 5776 32768
rect 5908 32759 5960 32768
rect 5908 32725 5917 32759
rect 5917 32725 5951 32759
rect 5951 32725 5960 32759
rect 5908 32716 5960 32725
rect 10232 32716 10284 32768
rect 11244 32716 11296 32768
rect 15108 32784 15160 32836
rect 16212 32852 16264 32904
rect 17132 32784 17184 32836
rect 17868 32852 17920 32904
rect 18880 32852 18932 32904
rect 12716 32759 12768 32768
rect 12716 32725 12725 32759
rect 12725 32725 12759 32759
rect 12759 32725 12768 32759
rect 12716 32716 12768 32725
rect 13268 32716 13320 32768
rect 13636 32716 13688 32768
rect 17408 32716 17460 32768
rect 19248 32920 19300 32972
rect 20996 32920 21048 32972
rect 24492 32920 24544 32972
rect 23480 32852 23532 32904
rect 25044 32895 25096 32904
rect 25044 32861 25053 32895
rect 25053 32861 25087 32895
rect 25087 32861 25096 32895
rect 25044 32852 25096 32861
rect 26332 32963 26384 32972
rect 26332 32929 26341 32963
rect 26341 32929 26375 32963
rect 26375 32929 26384 32963
rect 26332 32920 26384 32929
rect 26608 32920 26660 32972
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 29460 32988 29512 33040
rect 30104 33031 30156 33040
rect 30104 32997 30113 33031
rect 30113 32997 30147 33031
rect 30147 32997 30156 33031
rect 30104 32988 30156 32997
rect 28816 32963 28868 32972
rect 28816 32929 28825 32963
rect 28825 32929 28859 32963
rect 28859 32929 28868 32963
rect 28816 32920 28868 32929
rect 29644 32963 29696 32972
rect 29644 32929 29653 32963
rect 29653 32929 29687 32963
rect 29687 32929 29696 32963
rect 29644 32920 29696 32929
rect 19064 32784 19116 32836
rect 21272 32784 21324 32836
rect 22284 32784 22336 32836
rect 24584 32784 24636 32836
rect 18236 32759 18288 32768
rect 18236 32725 18245 32759
rect 18245 32725 18279 32759
rect 18279 32725 18288 32759
rect 18236 32716 18288 32725
rect 18972 32716 19024 32768
rect 22008 32716 22060 32768
rect 27344 32716 27396 32768
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 30932 32895 30984 32904
rect 30932 32861 30941 32895
rect 30941 32861 30975 32895
rect 30975 32861 30984 32895
rect 30932 32852 30984 32861
rect 31760 32920 31812 32972
rect 32128 32920 32180 32972
rect 31392 32895 31444 32904
rect 31392 32861 31401 32895
rect 31401 32861 31435 32895
rect 31435 32861 31444 32895
rect 31392 32852 31444 32861
rect 31484 32895 31536 32904
rect 31484 32861 31493 32895
rect 31493 32861 31527 32895
rect 31527 32861 31536 32895
rect 31484 32852 31536 32861
rect 31944 32852 31996 32904
rect 32956 32988 33008 33040
rect 33048 33031 33100 33040
rect 33048 32997 33057 33031
rect 33057 32997 33091 33031
rect 33091 32997 33100 33031
rect 33048 32988 33100 32997
rect 32496 32963 32548 32972
rect 32496 32929 32505 32963
rect 32505 32929 32539 32963
rect 32539 32929 32548 32963
rect 32496 32920 32548 32929
rect 33692 32988 33744 33040
rect 35532 32988 35584 33040
rect 33324 32920 33376 32972
rect 29552 32784 29604 32836
rect 31668 32784 31720 32836
rect 33232 32895 33284 32904
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 33508 32895 33560 32904
rect 33508 32861 33517 32895
rect 33517 32861 33551 32895
rect 33551 32861 33560 32895
rect 33508 32852 33560 32861
rect 33784 32895 33836 32904
rect 33784 32861 33793 32895
rect 33793 32861 33827 32895
rect 33827 32861 33836 32895
rect 33784 32852 33836 32861
rect 34336 32852 34388 32904
rect 35716 32920 35768 32972
rect 39028 32920 39080 32972
rect 37280 32895 37332 32904
rect 37280 32861 37289 32895
rect 37289 32861 37323 32895
rect 37323 32861 37332 32895
rect 37280 32852 37332 32861
rect 37372 32895 37424 32904
rect 37372 32861 37381 32895
rect 37381 32861 37415 32895
rect 37415 32861 37424 32895
rect 37372 32852 37424 32861
rect 39856 33056 39908 33108
rect 40224 33056 40276 33108
rect 40684 32920 40736 32972
rect 28632 32759 28684 32768
rect 28632 32725 28641 32759
rect 28641 32725 28675 32759
rect 28675 32725 28684 32759
rect 28632 32716 28684 32725
rect 32220 32716 32272 32768
rect 33876 32784 33928 32836
rect 34060 32827 34112 32836
rect 34060 32793 34069 32827
rect 34069 32793 34103 32827
rect 34103 32793 34112 32827
rect 34060 32784 34112 32793
rect 34520 32784 34572 32836
rect 36636 32784 36688 32836
rect 33324 32716 33376 32768
rect 38016 32759 38068 32768
rect 38016 32725 38025 32759
rect 38025 32725 38059 32759
rect 38059 32725 38068 32759
rect 38016 32716 38068 32725
rect 40408 32784 40460 32836
rect 40592 32784 40644 32836
rect 41144 32716 41196 32768
rect 43444 32716 43496 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 3240 32512 3292 32564
rect 3792 32555 3844 32564
rect 3792 32521 3801 32555
rect 3801 32521 3835 32555
rect 3835 32521 3844 32555
rect 3792 32512 3844 32521
rect 1768 32487 1820 32496
rect 1768 32453 1802 32487
rect 1802 32453 1820 32487
rect 1768 32444 1820 32453
rect 6460 32512 6512 32564
rect 6736 32555 6788 32564
rect 6736 32521 6745 32555
rect 6745 32521 6779 32555
rect 6779 32521 6788 32555
rect 6736 32512 6788 32521
rect 6828 32555 6880 32564
rect 6828 32521 6837 32555
rect 6837 32521 6871 32555
rect 6871 32521 6880 32555
rect 6828 32512 6880 32521
rect 7104 32512 7156 32564
rect 7196 32555 7248 32564
rect 7196 32521 7205 32555
rect 7205 32521 7239 32555
rect 7239 32521 7248 32555
rect 7196 32512 7248 32521
rect 7288 32512 7340 32564
rect 8024 32512 8076 32564
rect 8392 32512 8444 32564
rect 10140 32512 10192 32564
rect 10232 32512 10284 32564
rect 5172 32444 5224 32496
rect 3056 32376 3108 32428
rect 6092 32376 6144 32428
rect 1492 32351 1544 32360
rect 1492 32317 1501 32351
rect 1501 32317 1535 32351
rect 1535 32317 1544 32351
rect 1492 32308 1544 32317
rect 6276 32376 6328 32428
rect 7380 32240 7432 32292
rect 7656 32308 7708 32360
rect 9588 32444 9640 32496
rect 12716 32512 12768 32564
rect 10048 32376 10100 32428
rect 10232 32419 10284 32428
rect 10232 32385 10241 32419
rect 10241 32385 10275 32419
rect 10275 32385 10284 32419
rect 10232 32376 10284 32385
rect 12164 32419 12216 32428
rect 12164 32385 12173 32419
rect 12173 32385 12207 32419
rect 12207 32385 12216 32419
rect 12164 32376 12216 32385
rect 12256 32351 12308 32360
rect 12256 32317 12265 32351
rect 12265 32317 12299 32351
rect 12299 32317 12308 32351
rect 12256 32308 12308 32317
rect 10140 32240 10192 32292
rect 12440 32419 12492 32428
rect 12440 32385 12449 32419
rect 12449 32385 12483 32419
rect 12483 32385 12492 32419
rect 12440 32376 12492 32385
rect 13176 32512 13228 32564
rect 15108 32512 15160 32564
rect 15200 32512 15252 32564
rect 15936 32512 15988 32564
rect 15292 32444 15344 32496
rect 13176 32376 13228 32428
rect 13636 32419 13688 32428
rect 13636 32385 13645 32419
rect 13645 32385 13679 32419
rect 13679 32385 13688 32419
rect 13636 32376 13688 32385
rect 12992 32308 13044 32360
rect 15660 32376 15712 32428
rect 15752 32376 15804 32428
rect 16304 32512 16356 32564
rect 17040 32512 17092 32564
rect 17224 32512 17276 32564
rect 17408 32512 17460 32564
rect 17868 32512 17920 32564
rect 18236 32512 18288 32564
rect 18972 32512 19024 32564
rect 19064 32512 19116 32564
rect 6828 32172 6880 32224
rect 9496 32172 9548 32224
rect 10324 32172 10376 32224
rect 12716 32215 12768 32224
rect 12716 32181 12725 32215
rect 12725 32181 12759 32215
rect 12759 32181 12768 32215
rect 12716 32172 12768 32181
rect 13912 32172 13964 32224
rect 16212 32376 16264 32428
rect 16672 32308 16724 32360
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 17132 32376 17184 32428
rect 18328 32376 18380 32428
rect 18420 32376 18472 32428
rect 18788 32376 18840 32428
rect 17592 32240 17644 32292
rect 17224 32172 17276 32224
rect 23112 32512 23164 32564
rect 24768 32444 24820 32496
rect 26056 32512 26108 32564
rect 27344 32555 27396 32564
rect 27344 32521 27353 32555
rect 27353 32521 27387 32555
rect 27387 32521 27396 32555
rect 27344 32512 27396 32521
rect 28632 32512 28684 32564
rect 29644 32512 29696 32564
rect 30932 32555 30984 32564
rect 30932 32521 30941 32555
rect 30941 32521 30975 32555
rect 30975 32521 30984 32555
rect 30932 32512 30984 32521
rect 31392 32512 31444 32564
rect 33784 32512 33836 32564
rect 31760 32487 31812 32496
rect 31760 32453 31769 32487
rect 31769 32453 31803 32487
rect 31803 32453 31812 32487
rect 31760 32444 31812 32453
rect 32220 32444 32272 32496
rect 33600 32444 33652 32496
rect 43904 32512 43956 32564
rect 41144 32444 41196 32496
rect 21272 32419 21324 32428
rect 21272 32385 21281 32419
rect 21281 32385 21315 32419
rect 21315 32385 21324 32419
rect 21272 32376 21324 32385
rect 22836 32376 22888 32428
rect 28908 32376 28960 32428
rect 29920 32376 29972 32428
rect 30196 32376 30248 32428
rect 30840 32419 30892 32428
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 32404 32376 32456 32428
rect 32588 32376 32640 32428
rect 33048 32376 33100 32428
rect 33416 32376 33468 32428
rect 40132 32419 40184 32428
rect 40132 32385 40141 32419
rect 40141 32385 40175 32419
rect 40175 32385 40184 32419
rect 40132 32376 40184 32385
rect 21088 32351 21140 32360
rect 21088 32317 21097 32351
rect 21097 32317 21131 32351
rect 21131 32317 21140 32351
rect 21088 32308 21140 32317
rect 21824 32308 21876 32360
rect 25964 32351 26016 32360
rect 25964 32317 25973 32351
rect 25973 32317 26007 32351
rect 26007 32317 26016 32351
rect 25964 32308 26016 32317
rect 27436 32351 27488 32360
rect 27436 32317 27445 32351
rect 27445 32317 27479 32351
rect 27479 32317 27488 32351
rect 27436 32308 27488 32317
rect 27528 32308 27580 32360
rect 29368 32351 29420 32360
rect 29368 32317 29377 32351
rect 29377 32317 29411 32351
rect 29411 32317 29420 32351
rect 29368 32308 29420 32317
rect 33140 32308 33192 32360
rect 40408 32351 40460 32360
rect 40408 32317 40417 32351
rect 40417 32317 40451 32351
rect 40451 32317 40460 32351
rect 40408 32308 40460 32317
rect 28816 32240 28868 32292
rect 20536 32215 20588 32224
rect 20536 32181 20545 32215
rect 20545 32181 20579 32215
rect 20579 32181 20588 32215
rect 20536 32172 20588 32181
rect 22744 32172 22796 32224
rect 23572 32172 23624 32224
rect 26516 32215 26568 32224
rect 26516 32181 26525 32215
rect 26525 32181 26559 32215
rect 26559 32181 26568 32215
rect 26516 32172 26568 32181
rect 32680 32172 32732 32224
rect 33784 32172 33836 32224
rect 36636 32172 36688 32224
rect 36820 32172 36872 32224
rect 40684 32172 40736 32224
rect 41236 32172 41288 32224
rect 43812 32215 43864 32224
rect 43812 32181 43821 32215
rect 43821 32181 43855 32215
rect 43855 32181 43864 32215
rect 43812 32172 43864 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4620 31968 4672 32020
rect 6184 31968 6236 32020
rect 6736 31968 6788 32020
rect 7104 31968 7156 32020
rect 2412 31832 2464 31884
rect 10140 31900 10192 31952
rect 10324 32011 10376 32020
rect 10324 31977 10333 32011
rect 10333 31977 10367 32011
rect 10367 31977 10376 32011
rect 10324 31968 10376 31977
rect 11612 31968 11664 32020
rect 12348 31968 12400 32020
rect 14096 31968 14148 32020
rect 14832 31968 14884 32020
rect 15660 31968 15712 32020
rect 12808 31900 12860 31952
rect 5908 31832 5960 31884
rect 6460 31832 6512 31884
rect 5172 31807 5224 31816
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 7012 31764 7064 31816
rect 8300 31764 8352 31816
rect 8392 31764 8444 31816
rect 9496 31764 9548 31816
rect 9680 31764 9732 31816
rect 6828 31696 6880 31748
rect 9312 31739 9364 31748
rect 9312 31705 9321 31739
rect 9321 31705 9355 31739
rect 9355 31705 9364 31739
rect 12256 31832 12308 31884
rect 10048 31807 10100 31816
rect 10048 31773 10057 31807
rect 10057 31773 10091 31807
rect 10091 31773 10100 31807
rect 10048 31764 10100 31773
rect 10232 31764 10284 31816
rect 9312 31696 9364 31705
rect 10324 31739 10376 31748
rect 10324 31705 10333 31739
rect 10333 31705 10367 31739
rect 10367 31705 10376 31739
rect 10324 31696 10376 31705
rect 2412 31671 2464 31680
rect 2412 31637 2421 31671
rect 2421 31637 2455 31671
rect 2455 31637 2464 31671
rect 2412 31628 2464 31637
rect 3240 31628 3292 31680
rect 9404 31628 9456 31680
rect 9864 31628 9916 31680
rect 10048 31628 10100 31680
rect 11980 31764 12032 31816
rect 12164 31764 12216 31816
rect 13176 31900 13228 31952
rect 17776 31968 17828 32020
rect 18052 31968 18104 32020
rect 14280 31875 14332 31884
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14740 31832 14792 31884
rect 12256 31696 12308 31748
rect 13544 31764 13596 31816
rect 13636 31696 13688 31748
rect 13820 31739 13872 31748
rect 13820 31705 13829 31739
rect 13829 31705 13863 31739
rect 13863 31705 13872 31739
rect 13820 31696 13872 31705
rect 14372 31764 14424 31816
rect 14648 31764 14700 31816
rect 18144 31900 18196 31952
rect 20536 31968 20588 32020
rect 21088 31968 21140 32020
rect 18236 31832 18288 31884
rect 19156 31832 19208 31884
rect 19984 31832 20036 31884
rect 18420 31764 18472 31816
rect 14188 31696 14240 31748
rect 22192 31900 22244 31952
rect 21180 31875 21232 31884
rect 21180 31841 21189 31875
rect 21189 31841 21223 31875
rect 21223 31841 21232 31875
rect 21180 31832 21232 31841
rect 22744 31968 22796 32020
rect 22836 31968 22888 32020
rect 21272 31764 21324 31816
rect 23112 31875 23164 31884
rect 23112 31841 23121 31875
rect 23121 31841 23155 31875
rect 23155 31841 23164 31875
rect 23112 31832 23164 31841
rect 23204 31875 23256 31884
rect 23204 31841 23213 31875
rect 23213 31841 23247 31875
rect 23247 31841 23256 31875
rect 23204 31832 23256 31841
rect 23388 31900 23440 31952
rect 24492 31900 24544 31952
rect 28632 31968 28684 32020
rect 28908 31968 28960 32020
rect 30840 31968 30892 32020
rect 32404 32011 32456 32020
rect 32404 31977 32413 32011
rect 32413 31977 32447 32011
rect 32447 31977 32456 32011
rect 32404 31968 32456 31977
rect 33232 31968 33284 32020
rect 40132 31968 40184 32020
rect 24216 31832 24268 31884
rect 23664 31764 23716 31816
rect 23572 31696 23624 31748
rect 26424 31900 26476 31952
rect 26332 31832 26384 31884
rect 28540 31900 28592 31952
rect 28816 31900 28868 31952
rect 27712 31832 27764 31884
rect 32496 31900 32548 31952
rect 35900 31900 35952 31952
rect 25504 31764 25556 31816
rect 26240 31807 26292 31816
rect 26240 31773 26249 31807
rect 26249 31773 26283 31807
rect 26283 31773 26292 31807
rect 26240 31764 26292 31773
rect 26516 31807 26568 31816
rect 26516 31773 26525 31807
rect 26525 31773 26559 31807
rect 26559 31773 26568 31807
rect 26516 31764 26568 31773
rect 26700 31807 26752 31816
rect 26700 31773 26709 31807
rect 26709 31773 26743 31807
rect 26743 31773 26752 31807
rect 26700 31764 26752 31773
rect 29276 31764 29328 31816
rect 29828 31875 29880 31884
rect 29828 31841 29837 31875
rect 29837 31841 29871 31875
rect 29871 31841 29880 31875
rect 29828 31832 29880 31841
rect 32312 31807 32364 31816
rect 32312 31773 32321 31807
rect 32321 31773 32355 31807
rect 32355 31773 32364 31807
rect 32312 31764 32364 31773
rect 32496 31807 32548 31816
rect 32496 31773 32505 31807
rect 32505 31773 32539 31807
rect 32539 31773 32548 31807
rect 32496 31764 32548 31773
rect 34796 31764 34848 31816
rect 36544 31875 36596 31884
rect 36544 31841 36553 31875
rect 36553 31841 36587 31875
rect 36587 31841 36596 31875
rect 36544 31832 36596 31841
rect 36636 31875 36688 31884
rect 36636 31841 36645 31875
rect 36645 31841 36679 31875
rect 36679 31841 36688 31875
rect 36636 31832 36688 31841
rect 38660 31832 38712 31884
rect 38752 31832 38804 31884
rect 40500 31832 40552 31884
rect 41512 31832 41564 31884
rect 41236 31807 41288 31816
rect 41236 31773 41245 31807
rect 41245 31773 41279 31807
rect 41279 31773 41288 31807
rect 41236 31764 41288 31773
rect 42524 31807 42576 31816
rect 42524 31773 42533 31807
rect 42533 31773 42567 31807
rect 42567 31773 42576 31807
rect 42524 31764 42576 31773
rect 42800 31807 42852 31816
rect 42800 31773 42809 31807
rect 42809 31773 42843 31807
rect 42843 31773 42852 31807
rect 42800 31764 42852 31773
rect 27712 31696 27764 31748
rect 43536 31696 43588 31748
rect 20076 31628 20128 31680
rect 22100 31628 22152 31680
rect 22560 31671 22612 31680
rect 22560 31637 22569 31671
rect 22569 31637 22603 31671
rect 22603 31637 22612 31671
rect 22560 31628 22612 31637
rect 24124 31628 24176 31680
rect 24768 31628 24820 31680
rect 26332 31671 26384 31680
rect 26332 31637 26341 31671
rect 26341 31637 26375 31671
rect 26375 31637 26384 31671
rect 26332 31628 26384 31637
rect 33968 31628 34020 31680
rect 36452 31671 36504 31680
rect 36452 31637 36461 31671
rect 36461 31637 36495 31671
rect 36495 31637 36504 31671
rect 36452 31628 36504 31637
rect 38016 31628 38068 31680
rect 39488 31628 39540 31680
rect 44548 31671 44600 31680
rect 44548 31637 44557 31671
rect 44557 31637 44591 31671
rect 44591 31637 44600 31671
rect 44548 31628 44600 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2412 31424 2464 31476
rect 4068 31424 4120 31476
rect 4896 31356 4948 31408
rect 1492 31220 1544 31272
rect 2504 31263 2556 31272
rect 2504 31229 2513 31263
rect 2513 31229 2547 31263
rect 2547 31229 2556 31263
rect 2504 31220 2556 31229
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 3424 31220 3476 31272
rect 6460 31220 6512 31272
rect 7840 31263 7892 31272
rect 7840 31229 7849 31263
rect 7849 31229 7883 31263
rect 7883 31229 7892 31263
rect 7840 31220 7892 31229
rect 8300 31288 8352 31340
rect 9312 31424 9364 31476
rect 9680 31424 9732 31476
rect 10232 31424 10284 31476
rect 10324 31424 10376 31476
rect 8668 31331 8720 31340
rect 8668 31297 8677 31331
rect 8677 31297 8711 31331
rect 8711 31297 8720 31331
rect 8668 31288 8720 31297
rect 8944 31331 8996 31340
rect 8944 31297 8953 31331
rect 8953 31297 8987 31331
rect 8987 31297 8996 31331
rect 8944 31288 8996 31297
rect 9036 31331 9088 31340
rect 9036 31297 9045 31331
rect 9045 31297 9079 31331
rect 9079 31297 9088 31331
rect 9036 31288 9088 31297
rect 9496 31331 9548 31340
rect 9496 31297 9505 31331
rect 9505 31297 9539 31331
rect 9539 31297 9548 31331
rect 9496 31288 9548 31297
rect 10048 31399 10100 31408
rect 10048 31365 10057 31399
rect 10057 31365 10091 31399
rect 10091 31365 10100 31399
rect 10048 31356 10100 31365
rect 13360 31424 13412 31476
rect 14648 31424 14700 31476
rect 17776 31424 17828 31476
rect 21272 31467 21324 31476
rect 21272 31433 21281 31467
rect 21281 31433 21315 31467
rect 21315 31433 21324 31467
rect 21272 31424 21324 31433
rect 21548 31467 21600 31476
rect 21548 31433 21557 31467
rect 21557 31433 21591 31467
rect 21591 31433 21600 31467
rect 21548 31424 21600 31433
rect 13820 31356 13872 31408
rect 20076 31356 20128 31408
rect 22284 31424 22336 31476
rect 9588 31220 9640 31272
rect 1860 31084 1912 31136
rect 4068 31084 4120 31136
rect 9404 31152 9456 31204
rect 10232 31288 10284 31340
rect 10508 31288 10560 31340
rect 9864 31220 9916 31272
rect 8300 31127 8352 31136
rect 8300 31093 8309 31127
rect 8309 31093 8343 31127
rect 8343 31093 8352 31127
rect 8300 31084 8352 31093
rect 10508 31084 10560 31136
rect 10876 31288 10928 31340
rect 12348 31331 12400 31340
rect 12348 31297 12355 31331
rect 12355 31297 12400 31331
rect 12348 31288 12400 31297
rect 12532 31331 12584 31340
rect 12532 31297 12541 31331
rect 12541 31297 12575 31331
rect 12575 31297 12584 31331
rect 12532 31288 12584 31297
rect 12440 31152 12492 31204
rect 13084 31288 13136 31340
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 12808 31220 12860 31272
rect 12992 31220 13044 31272
rect 15568 31288 15620 31340
rect 15476 31220 15528 31272
rect 12808 31127 12860 31136
rect 12808 31093 12817 31127
rect 12817 31093 12851 31127
rect 12851 31093 12860 31127
rect 12808 31084 12860 31093
rect 12900 31084 12952 31136
rect 13176 31084 13228 31136
rect 13820 31152 13872 31204
rect 14096 31152 14148 31204
rect 14740 31084 14792 31136
rect 16212 31288 16264 31340
rect 18328 31331 18380 31340
rect 18328 31297 18337 31331
rect 18337 31297 18371 31331
rect 18371 31297 18380 31331
rect 18328 31288 18380 31297
rect 20812 31288 20864 31340
rect 22100 31399 22152 31408
rect 22100 31365 22109 31399
rect 22109 31365 22143 31399
rect 22143 31365 22152 31399
rect 22100 31356 22152 31365
rect 23664 31467 23716 31476
rect 23664 31433 23673 31467
rect 23673 31433 23707 31467
rect 23707 31433 23716 31467
rect 23664 31424 23716 31433
rect 24124 31467 24176 31476
rect 24124 31433 24133 31467
rect 24133 31433 24167 31467
rect 24167 31433 24176 31467
rect 24124 31424 24176 31433
rect 25964 31467 26016 31476
rect 25964 31433 25973 31467
rect 25973 31433 26007 31467
rect 26007 31433 26016 31467
rect 25964 31424 26016 31433
rect 26700 31424 26752 31476
rect 28632 31424 28684 31476
rect 29828 31467 29880 31476
rect 29828 31433 29837 31467
rect 29837 31433 29871 31467
rect 29871 31433 29880 31467
rect 29828 31424 29880 31433
rect 32312 31467 32364 31476
rect 32312 31433 32321 31467
rect 32321 31433 32355 31467
rect 32355 31433 32364 31467
rect 32312 31424 32364 31433
rect 32496 31424 32548 31476
rect 24768 31399 24820 31408
rect 24768 31365 24802 31399
rect 24802 31365 24820 31399
rect 24768 31356 24820 31365
rect 29920 31356 29972 31408
rect 19156 31220 19208 31272
rect 15476 31127 15528 31136
rect 15476 31093 15485 31127
rect 15485 31093 15519 31127
rect 15519 31093 15528 31127
rect 15476 31084 15528 31093
rect 15660 31084 15712 31136
rect 21824 31263 21876 31272
rect 21824 31229 21833 31263
rect 21833 31229 21867 31263
rect 21867 31229 21876 31263
rect 21824 31220 21876 31229
rect 26792 31288 26844 31340
rect 29368 31288 29420 31340
rect 24216 31263 24268 31272
rect 24216 31229 24225 31263
rect 24225 31229 24259 31263
rect 24259 31229 24268 31263
rect 24216 31220 24268 31229
rect 26240 31220 26292 31272
rect 26424 31263 26476 31272
rect 26424 31229 26433 31263
rect 26433 31229 26467 31263
rect 26467 31229 26476 31263
rect 26424 31220 26476 31229
rect 26516 31263 26568 31272
rect 26516 31229 26525 31263
rect 26525 31229 26559 31263
rect 26559 31229 26568 31263
rect 26516 31220 26568 31229
rect 27068 31220 27120 31272
rect 27528 31152 27580 31204
rect 30104 31220 30156 31272
rect 24768 31084 24820 31136
rect 33508 31331 33560 31340
rect 33508 31297 33517 31331
rect 33517 31297 33551 31331
rect 33551 31297 33560 31331
rect 33508 31288 33560 31297
rect 33600 31288 33652 31340
rect 33876 31424 33928 31476
rect 33968 31424 34020 31476
rect 39488 31467 39540 31476
rect 39488 31433 39497 31467
rect 39497 31433 39531 31467
rect 39531 31433 39540 31467
rect 39488 31424 39540 31433
rect 42524 31424 42576 31476
rect 43260 31424 43312 31476
rect 38016 31399 38068 31408
rect 38016 31365 38025 31399
rect 38025 31365 38059 31399
rect 38059 31365 38068 31399
rect 38016 31356 38068 31365
rect 43352 31356 43404 31408
rect 34060 31288 34112 31340
rect 35532 31288 35584 31340
rect 36360 31288 36412 31340
rect 37740 31331 37792 31340
rect 37740 31297 37749 31331
rect 37749 31297 37783 31331
rect 37783 31297 37792 31331
rect 37740 31288 37792 31297
rect 39120 31288 39172 31340
rect 43904 31331 43956 31340
rect 43904 31297 43913 31331
rect 43913 31297 43947 31331
rect 43947 31297 43956 31331
rect 43904 31288 43956 31297
rect 44548 31288 44600 31340
rect 33048 31152 33100 31204
rect 42892 31220 42944 31272
rect 43536 31220 43588 31272
rect 33876 31084 33928 31136
rect 35440 31152 35492 31204
rect 43076 31152 43128 31204
rect 35624 31084 35676 31136
rect 43444 31127 43496 31136
rect 43444 31093 43453 31127
rect 43453 31093 43487 31127
rect 43487 31093 43496 31127
rect 43444 31084 43496 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2780 30880 2832 30932
rect 3240 30855 3292 30864
rect 3240 30821 3249 30855
rect 3249 30821 3283 30855
rect 3283 30821 3292 30855
rect 3240 30812 3292 30821
rect 1492 30787 1544 30796
rect 1492 30753 1501 30787
rect 1501 30753 1535 30787
rect 1535 30753 1544 30787
rect 1492 30744 1544 30753
rect 1860 30744 1912 30796
rect 3424 30676 3476 30728
rect 4620 30880 4672 30932
rect 8944 30880 8996 30932
rect 9312 30880 9364 30932
rect 9404 30923 9456 30932
rect 9404 30889 9413 30923
rect 9413 30889 9447 30923
rect 9447 30889 9456 30923
rect 9404 30880 9456 30889
rect 11888 30880 11940 30932
rect 12808 30880 12860 30932
rect 13452 30880 13504 30932
rect 8300 30812 8352 30864
rect 10876 30812 10928 30864
rect 11244 30812 11296 30864
rect 9036 30744 9088 30796
rect 5172 30719 5224 30728
rect 5172 30685 5181 30719
rect 5181 30685 5215 30719
rect 5215 30685 5224 30719
rect 5172 30676 5224 30685
rect 8944 30719 8996 30728
rect 9496 30744 9548 30796
rect 8944 30685 8959 30719
rect 8959 30685 8993 30719
rect 8993 30685 8996 30719
rect 8944 30676 8996 30685
rect 9588 30719 9640 30728
rect 9588 30685 9597 30719
rect 9597 30685 9631 30719
rect 9631 30685 9640 30719
rect 9588 30676 9640 30685
rect 9772 30676 9824 30728
rect 3792 30608 3844 30660
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 11060 30676 11112 30728
rect 11888 30676 11940 30728
rect 12256 30676 12308 30728
rect 13544 30812 13596 30864
rect 12808 30787 12860 30796
rect 12808 30753 12817 30787
rect 12817 30753 12851 30787
rect 12851 30753 12860 30787
rect 12808 30744 12860 30753
rect 13176 30787 13228 30796
rect 13176 30753 13185 30787
rect 13185 30753 13219 30787
rect 13219 30753 13228 30787
rect 13176 30744 13228 30753
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 4160 30583 4212 30592
rect 4160 30549 4169 30583
rect 4169 30549 4203 30583
rect 4203 30549 4212 30583
rect 4160 30540 4212 30549
rect 4804 30540 4856 30592
rect 9864 30540 9916 30592
rect 11152 30583 11204 30592
rect 11152 30549 11161 30583
rect 11161 30549 11195 30583
rect 11195 30549 11204 30583
rect 11152 30540 11204 30549
rect 11336 30540 11388 30592
rect 13636 30719 13688 30728
rect 13636 30685 13645 30719
rect 13645 30685 13679 30719
rect 13679 30685 13688 30719
rect 13636 30676 13688 30685
rect 13912 30880 13964 30932
rect 15476 30880 15528 30932
rect 16488 30880 16540 30932
rect 18236 30880 18288 30932
rect 19340 30880 19392 30932
rect 21548 30880 21600 30932
rect 21824 30880 21876 30932
rect 16672 30787 16724 30796
rect 16672 30753 16681 30787
rect 16681 30753 16715 30787
rect 16715 30753 16724 30787
rect 16672 30744 16724 30753
rect 15292 30676 15344 30728
rect 15844 30719 15896 30728
rect 15844 30685 15853 30719
rect 15853 30685 15887 30719
rect 15887 30685 15896 30719
rect 15844 30676 15896 30685
rect 16488 30676 16540 30728
rect 26792 30923 26844 30932
rect 26792 30889 26801 30923
rect 26801 30889 26835 30923
rect 26835 30889 26844 30923
rect 26792 30880 26844 30889
rect 30104 30880 30156 30932
rect 33508 30923 33560 30932
rect 33508 30889 33517 30923
rect 33517 30889 33551 30923
rect 33551 30889 33560 30923
rect 33508 30880 33560 30889
rect 33876 30923 33928 30932
rect 33876 30889 33885 30923
rect 33885 30889 33919 30923
rect 33919 30889 33928 30923
rect 33876 30880 33928 30889
rect 43444 30880 43496 30932
rect 27804 30787 27856 30796
rect 27804 30753 27813 30787
rect 27813 30753 27847 30787
rect 27847 30753 27856 30787
rect 27804 30744 27856 30753
rect 30196 30744 30248 30796
rect 33324 30787 33376 30796
rect 33324 30753 33333 30787
rect 33333 30753 33367 30787
rect 33367 30753 33376 30787
rect 33324 30744 33376 30753
rect 35900 30787 35952 30796
rect 35900 30753 35909 30787
rect 35909 30753 35943 30787
rect 35943 30753 35952 30787
rect 35900 30744 35952 30753
rect 36452 30744 36504 30796
rect 43352 30812 43404 30864
rect 40316 30787 40368 30796
rect 40316 30753 40325 30787
rect 40325 30753 40359 30787
rect 40359 30753 40368 30787
rect 40316 30744 40368 30753
rect 42156 30744 42208 30796
rect 13912 30608 13964 30660
rect 14096 30651 14148 30660
rect 14096 30617 14105 30651
rect 14105 30617 14139 30651
rect 14139 30617 14148 30651
rect 14096 30608 14148 30617
rect 14832 30608 14884 30660
rect 16672 30608 16724 30660
rect 18236 30608 18288 30660
rect 19340 30608 19392 30660
rect 22560 30608 22612 30660
rect 13544 30540 13596 30592
rect 16212 30540 16264 30592
rect 16488 30583 16540 30592
rect 16488 30549 16497 30583
rect 16497 30549 16531 30583
rect 16531 30549 16540 30583
rect 16488 30540 16540 30549
rect 19432 30540 19484 30592
rect 24216 30583 24268 30592
rect 24216 30549 24225 30583
rect 24225 30549 24259 30583
rect 24259 30549 24268 30583
rect 24216 30540 24268 30549
rect 24768 30676 24820 30728
rect 26332 30676 26384 30728
rect 27160 30719 27212 30728
rect 27160 30685 27169 30719
rect 27169 30685 27203 30719
rect 27203 30685 27212 30719
rect 27160 30676 27212 30685
rect 29000 30676 29052 30728
rect 32956 30676 33008 30728
rect 34796 30676 34848 30728
rect 35440 30676 35492 30728
rect 35624 30719 35676 30728
rect 35624 30685 35633 30719
rect 35633 30685 35667 30719
rect 35667 30685 35676 30719
rect 35624 30676 35676 30685
rect 40224 30719 40276 30728
rect 40224 30685 40233 30719
rect 40233 30685 40267 30719
rect 40267 30685 40276 30719
rect 40224 30676 40276 30685
rect 43168 30719 43220 30728
rect 43168 30685 43177 30719
rect 43177 30685 43211 30719
rect 43211 30685 43220 30719
rect 43168 30676 43220 30685
rect 36360 30608 36412 30660
rect 25044 30540 25096 30592
rect 27344 30583 27396 30592
rect 27344 30549 27353 30583
rect 27353 30549 27387 30583
rect 27387 30549 27396 30583
rect 27344 30540 27396 30549
rect 27896 30540 27948 30592
rect 40592 30583 40644 30592
rect 40592 30549 40601 30583
rect 40601 30549 40635 30583
rect 40635 30549 40644 30583
rect 40592 30540 40644 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 2504 30336 2556 30388
rect 4804 30336 4856 30388
rect 4896 30268 4948 30320
rect 8668 30336 8720 30388
rect 6552 30311 6604 30320
rect 6552 30277 6561 30311
rect 6561 30277 6595 30311
rect 6595 30277 6604 30311
rect 6552 30268 6604 30277
rect 6644 30268 6696 30320
rect 5540 30064 5592 30116
rect 6736 30243 6788 30252
rect 6736 30209 6745 30243
rect 6745 30209 6779 30243
rect 6779 30209 6788 30243
rect 6736 30200 6788 30209
rect 6920 30311 6972 30320
rect 6920 30277 6929 30311
rect 6929 30277 6963 30311
rect 6963 30277 6972 30311
rect 6920 30268 6972 30277
rect 9588 30336 9640 30388
rect 12532 30336 12584 30388
rect 15844 30336 15896 30388
rect 10876 30268 10928 30320
rect 11152 30268 11204 30320
rect 15292 30268 15344 30320
rect 16672 30336 16724 30388
rect 17684 30336 17736 30388
rect 24124 30336 24176 30388
rect 5908 30132 5960 30184
rect 11336 30200 11388 30252
rect 18144 30268 18196 30320
rect 19432 30268 19484 30320
rect 20812 30268 20864 30320
rect 22192 30311 22244 30320
rect 22192 30277 22201 30311
rect 22201 30277 22235 30311
rect 22235 30277 22244 30311
rect 22192 30268 22244 30277
rect 27344 30268 27396 30320
rect 27712 30268 27764 30320
rect 32588 30268 32640 30320
rect 16580 30200 16632 30252
rect 18788 30200 18840 30252
rect 24216 30243 24268 30252
rect 24216 30209 24225 30243
rect 24225 30209 24259 30243
rect 24259 30209 24268 30243
rect 24216 30200 24268 30209
rect 26608 30243 26660 30252
rect 26608 30209 26617 30243
rect 26617 30209 26651 30243
rect 26651 30209 26660 30243
rect 26608 30200 26660 30209
rect 29920 30200 29972 30252
rect 12532 30175 12584 30184
rect 12532 30141 12541 30175
rect 12541 30141 12575 30175
rect 12575 30141 12584 30175
rect 12532 30132 12584 30141
rect 14096 30132 14148 30184
rect 16304 30132 16356 30184
rect 4896 29996 4948 30048
rect 7104 30064 7156 30116
rect 19156 30132 19208 30184
rect 19984 30132 20036 30184
rect 22836 30175 22888 30184
rect 22836 30141 22845 30175
rect 22845 30141 22879 30175
rect 22879 30141 22888 30175
rect 22836 30132 22888 30141
rect 26148 30132 26200 30184
rect 28448 30132 28500 30184
rect 29000 30132 29052 30184
rect 24584 30064 24636 30116
rect 6368 30039 6420 30048
rect 6368 30005 6377 30039
rect 6377 30005 6411 30039
rect 6411 30005 6420 30039
rect 6368 29996 6420 30005
rect 12716 29996 12768 30048
rect 16212 29996 16264 30048
rect 26792 30039 26844 30048
rect 26792 30005 26801 30039
rect 26801 30005 26835 30039
rect 26835 30005 26844 30039
rect 26792 29996 26844 30005
rect 30288 30132 30340 30184
rect 29552 30107 29604 30116
rect 29552 30073 29561 30107
rect 29561 30073 29595 30107
rect 29595 30073 29604 30107
rect 29552 30064 29604 30073
rect 33324 30336 33376 30388
rect 39488 30336 39540 30388
rect 40316 30336 40368 30388
rect 33508 30311 33560 30320
rect 33508 30277 33517 30311
rect 33517 30277 33551 30311
rect 33551 30277 33560 30311
rect 33508 30268 33560 30277
rect 33324 30243 33376 30252
rect 33324 30209 33333 30243
rect 33333 30209 33367 30243
rect 33367 30209 33376 30243
rect 33324 30200 33376 30209
rect 38108 30268 38160 30320
rect 41236 30268 41288 30320
rect 43536 30268 43588 30320
rect 29920 30039 29972 30048
rect 29920 30005 29929 30039
rect 29929 30005 29963 30039
rect 29963 30005 29972 30039
rect 29920 29996 29972 30005
rect 30012 29996 30064 30048
rect 32220 29996 32272 30048
rect 32956 30064 33008 30116
rect 34152 30064 34204 30116
rect 39120 30200 39172 30252
rect 38108 30175 38160 30184
rect 38108 30141 38117 30175
rect 38117 30141 38151 30175
rect 38151 30141 38160 30175
rect 38108 30132 38160 30141
rect 38752 30132 38804 30184
rect 39212 30175 39264 30184
rect 39212 30141 39221 30175
rect 39221 30141 39255 30175
rect 39255 30141 39264 30175
rect 39580 30243 39632 30252
rect 39580 30209 39589 30243
rect 39589 30209 39623 30243
rect 39623 30209 39632 30243
rect 39580 30200 39632 30209
rect 40132 30200 40184 30252
rect 41512 30200 41564 30252
rect 43168 30200 43220 30252
rect 43352 30243 43404 30252
rect 43352 30209 43361 30243
rect 43361 30209 43395 30243
rect 43395 30209 43404 30243
rect 43352 30200 43404 30209
rect 39212 30132 39264 30141
rect 40040 30132 40092 30184
rect 41328 30064 41380 30116
rect 43076 30064 43128 30116
rect 33140 29996 33192 30048
rect 34336 29996 34388 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 39304 30039 39356 30048
rect 39304 30005 39313 30039
rect 39313 30005 39347 30039
rect 39347 30005 39356 30039
rect 39304 29996 39356 30005
rect 39672 30039 39724 30048
rect 39672 30005 39681 30039
rect 39681 30005 39715 30039
rect 39715 30005 39724 30039
rect 39672 29996 39724 30005
rect 40500 29996 40552 30048
rect 41420 29996 41472 30048
rect 41972 29996 42024 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5172 29835 5224 29844
rect 5172 29801 5181 29835
rect 5181 29801 5215 29835
rect 5215 29801 5224 29835
rect 5172 29792 5224 29801
rect 6368 29792 6420 29844
rect 11244 29835 11296 29844
rect 11244 29801 11253 29835
rect 11253 29801 11287 29835
rect 11287 29801 11296 29835
rect 11244 29792 11296 29801
rect 12624 29792 12676 29844
rect 19340 29792 19392 29844
rect 27068 29835 27120 29844
rect 27068 29801 27077 29835
rect 27077 29801 27111 29835
rect 27111 29801 27120 29835
rect 27068 29792 27120 29801
rect 27160 29835 27212 29844
rect 27160 29801 27169 29835
rect 27169 29801 27203 29835
rect 27203 29801 27212 29835
rect 27160 29792 27212 29801
rect 28632 29792 28684 29844
rect 29000 29792 29052 29844
rect 29368 29835 29420 29844
rect 29368 29801 29377 29835
rect 29377 29801 29411 29835
rect 29411 29801 29420 29835
rect 29368 29792 29420 29801
rect 29920 29792 29972 29844
rect 30196 29835 30248 29844
rect 30196 29801 30205 29835
rect 30205 29801 30239 29835
rect 30239 29801 30248 29835
rect 30196 29792 30248 29801
rect 30288 29792 30340 29844
rect 32312 29792 32364 29844
rect 4988 29588 5040 29640
rect 5816 29588 5868 29640
rect 5908 29631 5960 29640
rect 5908 29597 5917 29631
rect 5917 29597 5951 29631
rect 5951 29597 5960 29631
rect 5908 29588 5960 29597
rect 27528 29724 27580 29776
rect 6644 29656 6696 29708
rect 6092 29631 6144 29640
rect 6092 29597 6101 29631
rect 6101 29597 6135 29631
rect 6135 29597 6144 29631
rect 6092 29588 6144 29597
rect 6184 29588 6236 29640
rect 6276 29631 6328 29640
rect 6276 29597 6285 29631
rect 6285 29597 6319 29631
rect 6319 29597 6328 29631
rect 6276 29588 6328 29597
rect 12256 29656 12308 29708
rect 7104 29520 7156 29572
rect 14924 29588 14976 29640
rect 21180 29656 21232 29708
rect 28448 29656 28500 29708
rect 15568 29588 15620 29640
rect 16304 29588 16356 29640
rect 18512 29588 18564 29640
rect 19984 29588 20036 29640
rect 22928 29631 22980 29640
rect 22928 29597 22937 29631
rect 22937 29597 22971 29631
rect 22971 29597 22980 29631
rect 22928 29588 22980 29597
rect 24860 29588 24912 29640
rect 25780 29588 25832 29640
rect 30104 29724 30156 29776
rect 30012 29656 30064 29708
rect 29552 29588 29604 29640
rect 24400 29563 24452 29572
rect 24400 29529 24409 29563
rect 24409 29529 24443 29563
rect 24443 29529 24452 29563
rect 24400 29520 24452 29529
rect 28632 29520 28684 29572
rect 10784 29452 10836 29504
rect 11428 29452 11480 29504
rect 15200 29452 15252 29504
rect 15384 29495 15436 29504
rect 15384 29461 15393 29495
rect 15393 29461 15427 29495
rect 15427 29461 15436 29495
rect 15384 29452 15436 29461
rect 21732 29452 21784 29504
rect 22100 29495 22152 29504
rect 22100 29461 22109 29495
rect 22109 29461 22143 29495
rect 22143 29461 22152 29495
rect 22100 29452 22152 29461
rect 25504 29495 25556 29504
rect 25504 29461 25513 29495
rect 25513 29461 25547 29495
rect 25547 29461 25556 29495
rect 25504 29452 25556 29461
rect 30472 29631 30524 29640
rect 30472 29597 30481 29631
rect 30481 29597 30515 29631
rect 30515 29597 30524 29631
rect 30472 29588 30524 29597
rect 32220 29724 32272 29776
rect 32956 29835 33008 29844
rect 32956 29801 32965 29835
rect 32965 29801 32999 29835
rect 32999 29801 33008 29835
rect 32956 29792 33008 29801
rect 33324 29792 33376 29844
rect 33508 29835 33560 29844
rect 33508 29801 33517 29835
rect 33517 29801 33551 29835
rect 33551 29801 33560 29835
rect 33508 29792 33560 29801
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33600 29588 33652 29597
rect 35624 29656 35676 29708
rect 33324 29563 33376 29572
rect 33324 29529 33333 29563
rect 33333 29529 33367 29563
rect 33367 29529 33376 29563
rect 33324 29520 33376 29529
rect 32220 29452 32272 29504
rect 33232 29452 33284 29504
rect 34152 29452 34204 29504
rect 35624 29563 35676 29572
rect 35624 29529 35633 29563
rect 35633 29529 35667 29563
rect 35667 29529 35676 29563
rect 35624 29520 35676 29529
rect 36360 29520 36412 29572
rect 39304 29792 39356 29844
rect 39672 29792 39724 29844
rect 40132 29835 40184 29844
rect 40132 29801 40141 29835
rect 40141 29801 40175 29835
rect 40175 29801 40184 29835
rect 40132 29792 40184 29801
rect 41236 29792 41288 29844
rect 41328 29792 41380 29844
rect 40224 29656 40276 29708
rect 39856 29588 39908 29640
rect 40500 29631 40552 29640
rect 40500 29597 40509 29631
rect 40509 29597 40543 29631
rect 40543 29597 40552 29631
rect 40500 29588 40552 29597
rect 40776 29631 40828 29640
rect 40776 29597 40785 29631
rect 40785 29597 40819 29631
rect 40819 29597 40828 29631
rect 40776 29588 40828 29597
rect 41972 29724 42024 29776
rect 42984 29835 43036 29844
rect 42984 29801 42993 29835
rect 42993 29801 43027 29835
rect 43027 29801 43036 29835
rect 42984 29792 43036 29801
rect 43076 29792 43128 29844
rect 43996 29792 44048 29844
rect 41420 29699 41472 29708
rect 41420 29665 41429 29699
rect 41429 29665 41463 29699
rect 41463 29665 41472 29699
rect 41420 29656 41472 29665
rect 41512 29699 41564 29708
rect 41512 29665 41521 29699
rect 41521 29665 41555 29699
rect 41555 29665 41564 29699
rect 41512 29656 41564 29665
rect 41328 29631 41380 29640
rect 41328 29597 41337 29631
rect 41337 29597 41371 29631
rect 41371 29597 41380 29631
rect 41328 29588 41380 29597
rect 43536 29724 43588 29776
rect 43904 29724 43956 29776
rect 39948 29520 40000 29572
rect 37096 29495 37148 29504
rect 37096 29461 37105 29495
rect 37105 29461 37139 29495
rect 37139 29461 37148 29495
rect 37096 29452 37148 29461
rect 37280 29452 37332 29504
rect 39580 29452 39632 29504
rect 40960 29452 41012 29504
rect 41696 29452 41748 29504
rect 41788 29452 41840 29504
rect 42708 29631 42760 29640
rect 42708 29597 42717 29631
rect 42717 29597 42751 29631
rect 42751 29597 42760 29631
rect 42708 29588 42760 29597
rect 43444 29588 43496 29640
rect 44088 29656 44140 29708
rect 42892 29520 42944 29572
rect 43352 29520 43404 29572
rect 43904 29588 43956 29640
rect 41972 29452 42024 29504
rect 43812 29495 43864 29504
rect 43812 29461 43821 29495
rect 43821 29461 43855 29495
rect 43855 29461 43864 29495
rect 43812 29452 43864 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5540 29248 5592 29300
rect 5908 29248 5960 29300
rect 6092 29248 6144 29300
rect 11336 29291 11388 29300
rect 11336 29257 11345 29291
rect 11345 29257 11379 29291
rect 11379 29257 11388 29291
rect 11336 29248 11388 29257
rect 12532 29248 12584 29300
rect 13912 29248 13964 29300
rect 10876 29180 10928 29232
rect 6644 29112 6696 29164
rect 6736 29112 6788 29164
rect 10692 29155 10744 29164
rect 10692 29121 10701 29155
rect 10701 29121 10735 29155
rect 10735 29121 10744 29155
rect 10692 29112 10744 29121
rect 10784 29155 10836 29164
rect 10784 29121 10794 29155
rect 10794 29121 10828 29155
rect 10828 29121 10836 29155
rect 10784 29112 10836 29121
rect 11244 29112 11296 29164
rect 11428 29112 11480 29164
rect 12256 29155 12308 29164
rect 12256 29121 12266 29155
rect 12266 29121 12300 29155
rect 12300 29121 12308 29155
rect 12256 29112 12308 29121
rect 12900 29044 12952 29096
rect 13084 29112 13136 29164
rect 13176 29112 13228 29164
rect 15200 29248 15252 29300
rect 14924 29223 14976 29232
rect 14924 29189 14933 29223
rect 14933 29189 14967 29223
rect 14967 29189 14976 29223
rect 14924 29180 14976 29189
rect 15292 29223 15344 29232
rect 15292 29189 15301 29223
rect 15301 29189 15335 29223
rect 15335 29189 15344 29223
rect 15292 29180 15344 29189
rect 16304 29248 16356 29300
rect 18512 29248 18564 29300
rect 22836 29248 22888 29300
rect 24860 29291 24912 29300
rect 24860 29257 24869 29291
rect 24869 29257 24903 29291
rect 24903 29257 24912 29291
rect 24860 29248 24912 29257
rect 30012 29248 30064 29300
rect 15016 29155 15068 29164
rect 15016 29121 15061 29155
rect 15061 29121 15068 29155
rect 15016 29112 15068 29121
rect 15200 29155 15252 29164
rect 15200 29121 15209 29155
rect 15209 29121 15243 29155
rect 15243 29121 15252 29155
rect 15200 29112 15252 29121
rect 15384 29112 15436 29164
rect 18236 29180 18288 29232
rect 22100 29223 22152 29232
rect 22100 29189 22123 29223
rect 22123 29189 22152 29223
rect 22100 29180 22152 29189
rect 15660 29044 15712 29096
rect 18788 29112 18840 29164
rect 6644 28976 6696 29028
rect 6000 28908 6052 28960
rect 9496 28976 9548 29028
rect 7932 28908 7984 28960
rect 11060 28908 11112 28960
rect 13268 28908 13320 28960
rect 14464 28908 14516 28960
rect 16672 29087 16724 29096
rect 16672 29053 16681 29087
rect 16681 29053 16715 29087
rect 16715 29053 16724 29087
rect 16672 29044 16724 29053
rect 17684 29044 17736 29096
rect 18972 29155 19024 29164
rect 18972 29121 18981 29155
rect 18981 29121 19015 29155
rect 19015 29121 19024 29155
rect 18972 29112 19024 29121
rect 19248 29112 19300 29164
rect 21364 29112 21416 29164
rect 23756 29155 23808 29164
rect 23756 29121 23790 29155
rect 23790 29121 23808 29155
rect 23756 29112 23808 29121
rect 25044 29180 25096 29232
rect 26792 29180 26844 29232
rect 27712 29180 27764 29232
rect 30472 29180 30524 29232
rect 30104 29112 30156 29164
rect 32220 29291 32272 29300
rect 32220 29257 32229 29291
rect 32229 29257 32263 29291
rect 32263 29257 32272 29291
rect 32220 29248 32272 29257
rect 33140 29248 33192 29300
rect 33600 29248 33652 29300
rect 35624 29248 35676 29300
rect 37096 29248 37148 29300
rect 34152 29180 34204 29232
rect 32680 29112 32732 29164
rect 33232 29155 33284 29164
rect 33232 29121 33241 29155
rect 33241 29121 33275 29155
rect 33275 29121 33284 29155
rect 33232 29112 33284 29121
rect 33324 29112 33376 29164
rect 33508 29112 33560 29164
rect 34796 29112 34848 29164
rect 37464 29180 37516 29232
rect 18512 28951 18564 28960
rect 18512 28917 18521 28951
rect 18521 28917 18555 28951
rect 18555 28917 18564 28951
rect 18512 28908 18564 28917
rect 21548 29044 21600 29096
rect 24768 29044 24820 29096
rect 19432 28976 19484 29028
rect 20260 28908 20312 28960
rect 26148 28976 26200 29028
rect 28448 29044 28500 29096
rect 34060 29044 34112 29096
rect 39028 29112 39080 29164
rect 39212 29248 39264 29300
rect 39396 29248 39448 29300
rect 39856 29291 39908 29300
rect 39856 29257 39865 29291
rect 39865 29257 39899 29291
rect 39899 29257 39908 29291
rect 39856 29248 39908 29257
rect 40132 29248 40184 29300
rect 40224 29248 40276 29300
rect 40776 29291 40828 29300
rect 40776 29257 40778 29291
rect 40778 29257 40812 29291
rect 40812 29257 40828 29291
rect 40776 29248 40828 29257
rect 37280 29087 37332 29096
rect 37280 29053 37289 29087
rect 37289 29053 37323 29087
rect 37323 29053 37332 29087
rect 37280 29044 37332 29053
rect 32312 28976 32364 29028
rect 38752 29044 38804 29096
rect 39948 29180 40000 29232
rect 39488 29155 39540 29164
rect 39488 29121 39497 29155
rect 39497 29121 39531 29155
rect 39531 29121 39540 29155
rect 39488 29112 39540 29121
rect 40408 29112 40460 29164
rect 40868 29155 40920 29164
rect 40868 29121 40877 29155
rect 40877 29121 40911 29155
rect 40911 29121 40920 29155
rect 40868 29112 40920 29121
rect 39948 29044 40000 29096
rect 41788 29248 41840 29300
rect 42984 29248 43036 29300
rect 43260 29248 43312 29300
rect 43352 29248 43404 29300
rect 43812 29248 43864 29300
rect 43904 29248 43956 29300
rect 41512 29180 41564 29232
rect 41328 29112 41380 29164
rect 42708 29180 42760 29232
rect 40040 28976 40092 29028
rect 21272 28908 21324 28960
rect 28632 28908 28684 28960
rect 33140 28951 33192 28960
rect 33140 28917 33149 28951
rect 33149 28917 33183 28951
rect 33183 28917 33192 28951
rect 33140 28908 33192 28917
rect 41236 29087 41288 29096
rect 41236 29053 41245 29087
rect 41245 29053 41279 29087
rect 41279 29053 41288 29087
rect 41236 29044 41288 29053
rect 41972 29112 42024 29164
rect 42156 29112 42208 29164
rect 42248 29155 42300 29164
rect 42248 29121 42257 29155
rect 42257 29121 42291 29155
rect 42291 29121 42300 29155
rect 42248 29112 42300 29121
rect 42892 29112 42944 29164
rect 40868 28976 40920 29028
rect 41236 28908 41288 28960
rect 42616 29019 42668 29028
rect 42616 28985 42625 29019
rect 42625 28985 42659 29019
rect 42659 28985 42668 29019
rect 42616 28976 42668 28985
rect 43168 29112 43220 29164
rect 43444 29044 43496 29096
rect 43720 29155 43772 29164
rect 43720 29121 43729 29155
rect 43729 29121 43763 29155
rect 43763 29121 43772 29155
rect 43720 29112 43772 29121
rect 43812 29087 43864 29096
rect 43812 29053 43821 29087
rect 43821 29053 43855 29087
rect 43855 29053 43864 29087
rect 43812 29044 43864 29053
rect 43904 29087 43956 29096
rect 43904 29053 43913 29087
rect 43913 29053 43947 29087
rect 43947 29053 43956 29087
rect 43904 29044 43956 29053
rect 44088 29044 44140 29096
rect 43904 28908 43956 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6736 28704 6788 28756
rect 7932 28704 7984 28756
rect 5264 28611 5316 28620
rect 5264 28577 5273 28611
rect 5273 28577 5307 28611
rect 5307 28577 5316 28611
rect 5264 28568 5316 28577
rect 6000 28568 6052 28620
rect 8300 28636 8352 28688
rect 5816 28432 5868 28484
rect 6000 28432 6052 28484
rect 5448 28364 5500 28416
rect 5632 28407 5684 28416
rect 5632 28373 5641 28407
rect 5641 28373 5675 28407
rect 5675 28373 5684 28407
rect 5632 28364 5684 28373
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 6828 28500 6880 28552
rect 6368 28407 6420 28416
rect 6368 28373 6377 28407
rect 6377 28373 6411 28407
rect 6411 28373 6420 28407
rect 9128 28747 9180 28756
rect 9128 28713 9137 28747
rect 9137 28713 9171 28747
rect 9171 28713 9180 28747
rect 9128 28704 9180 28713
rect 10692 28704 10744 28756
rect 11244 28747 11296 28756
rect 11244 28713 11253 28747
rect 11253 28713 11287 28747
rect 11287 28713 11296 28747
rect 11244 28704 11296 28713
rect 12900 28747 12952 28756
rect 12900 28713 12909 28747
rect 12909 28713 12943 28747
rect 12943 28713 12952 28747
rect 12900 28704 12952 28713
rect 13544 28704 13596 28756
rect 15200 28704 15252 28756
rect 12716 28636 12768 28688
rect 13268 28636 13320 28688
rect 13820 28636 13872 28688
rect 8668 28568 8720 28620
rect 9220 28568 9272 28620
rect 9496 28568 9548 28620
rect 11060 28568 11112 28620
rect 7932 28543 7984 28552
rect 7932 28509 7941 28543
rect 7941 28509 7975 28543
rect 7975 28509 7984 28543
rect 7932 28500 7984 28509
rect 8484 28500 8536 28552
rect 10600 28500 10652 28552
rect 13452 28611 13504 28620
rect 13452 28577 13461 28611
rect 13461 28577 13495 28611
rect 13495 28577 13504 28611
rect 13452 28568 13504 28577
rect 16028 28568 16080 28620
rect 16396 28568 16448 28620
rect 13084 28543 13136 28552
rect 13084 28509 13093 28543
rect 13093 28509 13127 28543
rect 13127 28509 13136 28543
rect 13084 28500 13136 28509
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 13176 28500 13228 28509
rect 8576 28432 8628 28484
rect 8668 28475 8720 28484
rect 8668 28441 8677 28475
rect 8677 28441 8711 28475
rect 8711 28441 8720 28475
rect 8668 28432 8720 28441
rect 8944 28475 8996 28484
rect 8944 28441 8953 28475
rect 8953 28441 8987 28475
rect 8987 28441 8996 28475
rect 8944 28432 8996 28441
rect 13544 28475 13596 28484
rect 13544 28441 13553 28475
rect 13553 28441 13587 28475
rect 13587 28441 13596 28475
rect 13544 28432 13596 28441
rect 14464 28500 14516 28552
rect 15936 28500 15988 28552
rect 17132 28500 17184 28552
rect 18512 28704 18564 28756
rect 18972 28704 19024 28756
rect 21364 28747 21416 28756
rect 21364 28713 21373 28747
rect 21373 28713 21407 28747
rect 21407 28713 21416 28747
rect 21364 28704 21416 28713
rect 21456 28704 21508 28756
rect 22928 28704 22980 28756
rect 26424 28704 26476 28756
rect 26608 28704 26660 28756
rect 34796 28704 34848 28756
rect 17684 28543 17736 28552
rect 17684 28509 17693 28543
rect 17693 28509 17727 28543
rect 17727 28509 17736 28543
rect 17684 28500 17736 28509
rect 18788 28500 18840 28552
rect 19064 28568 19116 28620
rect 24216 28679 24268 28688
rect 24216 28645 24225 28679
rect 24225 28645 24259 28679
rect 24259 28645 24268 28679
rect 24216 28636 24268 28645
rect 33416 28636 33468 28688
rect 33876 28636 33928 28688
rect 35624 28636 35676 28688
rect 39120 28636 39172 28688
rect 21272 28611 21324 28620
rect 21272 28577 21281 28611
rect 21281 28577 21315 28611
rect 21315 28577 21324 28611
rect 21272 28568 21324 28577
rect 22008 28611 22060 28620
rect 22008 28577 22017 28611
rect 22017 28577 22051 28611
rect 22051 28577 22060 28611
rect 22008 28568 22060 28577
rect 23296 28568 23348 28620
rect 23480 28568 23532 28620
rect 27528 28568 27580 28620
rect 33048 28568 33100 28620
rect 34520 28568 34572 28620
rect 36084 28568 36136 28620
rect 38752 28611 38804 28620
rect 38752 28577 38761 28611
rect 38761 28577 38795 28611
rect 38795 28577 38804 28611
rect 38752 28568 38804 28577
rect 40408 28636 40460 28688
rect 19156 28500 19208 28552
rect 21732 28543 21784 28552
rect 21732 28509 21741 28543
rect 21741 28509 21775 28543
rect 21775 28509 21784 28543
rect 21732 28500 21784 28509
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 23940 28500 23992 28552
rect 24400 28500 24452 28552
rect 24860 28500 24912 28552
rect 28632 28500 28684 28552
rect 32680 28543 32732 28552
rect 32680 28509 32689 28543
rect 32689 28509 32723 28543
rect 32723 28509 32732 28543
rect 32680 28500 32732 28509
rect 33140 28500 33192 28552
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 19432 28432 19484 28484
rect 6368 28364 6420 28373
rect 8300 28407 8352 28416
rect 8300 28373 8309 28407
rect 8309 28373 8343 28407
rect 8343 28373 8352 28407
rect 8300 28364 8352 28373
rect 9036 28364 9088 28416
rect 9680 28364 9732 28416
rect 13820 28364 13872 28416
rect 14372 28364 14424 28416
rect 14832 28364 14884 28416
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 19248 28364 19300 28416
rect 25412 28432 25464 28484
rect 23020 28364 23072 28416
rect 31852 28432 31904 28484
rect 32680 28364 32732 28416
rect 33876 28475 33928 28484
rect 33876 28441 33911 28475
rect 33911 28441 33928 28475
rect 34152 28543 34204 28552
rect 34152 28509 34161 28543
rect 34161 28509 34195 28543
rect 34195 28509 34204 28543
rect 34152 28500 34204 28509
rect 34336 28543 34388 28552
rect 34336 28509 34345 28543
rect 34345 28509 34379 28543
rect 34379 28509 34388 28543
rect 34336 28500 34388 28509
rect 33876 28432 33928 28441
rect 34612 28432 34664 28484
rect 35900 28500 35952 28552
rect 38936 28543 38988 28552
rect 38936 28509 38945 28543
rect 38945 28509 38979 28543
rect 38979 28509 38988 28543
rect 38936 28500 38988 28509
rect 39396 28543 39448 28552
rect 39396 28509 39405 28543
rect 39405 28509 39439 28543
rect 39439 28509 39448 28543
rect 39396 28500 39448 28509
rect 35992 28364 36044 28416
rect 39764 28568 39816 28620
rect 42800 28704 42852 28756
rect 44088 28636 44140 28688
rect 42248 28568 42300 28620
rect 43444 28568 43496 28620
rect 40040 28543 40092 28552
rect 40040 28509 40049 28543
rect 40049 28509 40083 28543
rect 40083 28509 40092 28543
rect 40040 28500 40092 28509
rect 40316 28500 40368 28552
rect 40592 28500 40644 28552
rect 40868 28543 40920 28552
rect 40868 28509 40877 28543
rect 40877 28509 40911 28543
rect 40911 28509 40920 28543
rect 40868 28500 40920 28509
rect 41696 28500 41748 28552
rect 43536 28500 43588 28552
rect 43996 28500 44048 28552
rect 39948 28432 40000 28484
rect 43260 28432 43312 28484
rect 42892 28364 42944 28416
rect 43812 28364 43864 28416
rect 44180 28364 44232 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5264 28160 5316 28212
rect 4804 28092 4856 28144
rect 6184 28160 6236 28212
rect 6552 28160 6604 28212
rect 5632 28135 5684 28144
rect 5632 28101 5641 28135
rect 5641 28101 5675 28135
rect 5675 28101 5684 28135
rect 5632 28092 5684 28101
rect 940 28024 992 28076
rect 5540 28067 5592 28076
rect 5540 28033 5549 28067
rect 5549 28033 5583 28067
rect 5583 28033 5592 28067
rect 5540 28024 5592 28033
rect 5724 28024 5776 28076
rect 4804 27956 4856 28008
rect 6368 28067 6420 28076
rect 6368 28033 6377 28067
rect 6377 28033 6411 28067
rect 6411 28033 6420 28067
rect 6368 28024 6420 28033
rect 7840 28160 7892 28212
rect 9036 28160 9088 28212
rect 9404 28160 9456 28212
rect 7104 28092 7156 28144
rect 9220 28092 9272 28144
rect 6828 28024 6880 28076
rect 8116 28024 8168 28076
rect 9036 27956 9088 28008
rect 12440 28092 12492 28144
rect 9956 28024 10008 28076
rect 12716 28092 12768 28144
rect 1768 27820 1820 27872
rect 6920 27820 6972 27872
rect 8392 27820 8444 27872
rect 11060 27999 11112 28008
rect 11060 27965 11069 27999
rect 11069 27965 11103 27999
rect 11103 27965 11112 27999
rect 11060 27956 11112 27965
rect 11336 27999 11388 28008
rect 11336 27965 11345 27999
rect 11345 27965 11379 27999
rect 11379 27965 11388 27999
rect 11336 27956 11388 27965
rect 13452 28092 13504 28144
rect 13544 28092 13596 28144
rect 14280 28092 14332 28144
rect 13636 28067 13688 28076
rect 13636 28033 13645 28067
rect 13645 28033 13679 28067
rect 13679 28033 13688 28067
rect 13636 28024 13688 28033
rect 17592 28160 17644 28212
rect 21732 28160 21784 28212
rect 23756 28160 23808 28212
rect 24216 28160 24268 28212
rect 25412 28203 25464 28212
rect 25412 28169 25421 28203
rect 25421 28169 25455 28203
rect 25455 28169 25464 28203
rect 25412 28160 25464 28169
rect 14832 28135 14884 28144
rect 14832 28101 14849 28135
rect 14849 28101 14884 28135
rect 14832 28092 14884 28101
rect 16028 28092 16080 28144
rect 12532 27888 12584 27940
rect 14372 27999 14424 28008
rect 14372 27965 14381 27999
rect 14381 27965 14415 27999
rect 14415 27965 14424 27999
rect 14372 27956 14424 27965
rect 14464 27956 14516 28008
rect 15016 27956 15068 28008
rect 15752 28024 15804 28076
rect 19248 28092 19300 28144
rect 19156 28024 19208 28076
rect 20260 28067 20312 28076
rect 20260 28033 20294 28067
rect 20294 28033 20312 28067
rect 20260 28024 20312 28033
rect 21548 28024 21600 28076
rect 27436 28160 27488 28212
rect 38936 28203 38988 28212
rect 38936 28169 38945 28203
rect 38945 28169 38979 28203
rect 38979 28169 38988 28203
rect 38936 28160 38988 28169
rect 39764 28203 39816 28212
rect 39764 28169 39773 28203
rect 39773 28169 39807 28203
rect 39807 28169 39816 28203
rect 39764 28160 39816 28169
rect 42892 28160 42944 28212
rect 42984 28160 43036 28212
rect 43352 28160 43404 28212
rect 44088 28160 44140 28212
rect 44180 28160 44232 28212
rect 15384 27956 15436 28008
rect 17132 27956 17184 28008
rect 19064 27956 19116 28008
rect 12808 27863 12860 27872
rect 12808 27829 12817 27863
rect 12817 27829 12851 27863
rect 12851 27829 12860 27863
rect 12808 27820 12860 27829
rect 13636 27820 13688 27872
rect 23480 27956 23532 28008
rect 24676 27999 24728 28008
rect 24676 27965 24685 27999
rect 24685 27965 24719 27999
rect 24719 27965 24728 27999
rect 24676 27956 24728 27965
rect 24860 27999 24912 28008
rect 24860 27965 24869 27999
rect 24869 27965 24903 27999
rect 24903 27965 24912 27999
rect 24860 27956 24912 27965
rect 26424 28024 26476 28076
rect 34704 28024 34756 28076
rect 35256 28067 35308 28076
rect 35256 28033 35265 28067
rect 35265 28033 35299 28067
rect 35299 28033 35308 28067
rect 35256 28024 35308 28033
rect 35440 28024 35492 28076
rect 38844 28067 38896 28076
rect 38844 28033 38853 28067
rect 38853 28033 38887 28067
rect 38887 28033 38896 28067
rect 38844 28024 38896 28033
rect 39304 28024 39356 28076
rect 39488 28067 39540 28076
rect 39488 28033 39497 28067
rect 39497 28033 39531 28067
rect 39531 28033 39540 28067
rect 39488 28024 39540 28033
rect 40316 28024 40368 28076
rect 41328 28024 41380 28076
rect 42984 28067 43036 28076
rect 42984 28033 42993 28067
rect 42993 28033 43027 28067
rect 43027 28033 43036 28067
rect 42984 28024 43036 28033
rect 36728 27999 36780 28008
rect 14096 27820 14148 27872
rect 14280 27820 14332 27872
rect 14924 27820 14976 27872
rect 34796 27863 34848 27872
rect 34796 27829 34805 27863
rect 34805 27829 34839 27863
rect 34839 27829 34848 27863
rect 34796 27820 34848 27829
rect 36728 27965 36737 27999
rect 36737 27965 36771 27999
rect 36771 27965 36780 27999
rect 36728 27956 36780 27965
rect 43260 27956 43312 28008
rect 43904 28067 43956 28076
rect 43904 28033 43913 28067
rect 43913 28033 43947 28067
rect 43947 28033 43956 28067
rect 43904 28024 43956 28033
rect 43168 27888 43220 27940
rect 43444 27888 43496 27940
rect 35900 27820 35952 27872
rect 36084 27820 36136 27872
rect 36176 27863 36228 27872
rect 36176 27829 36185 27863
rect 36185 27829 36219 27863
rect 36219 27829 36228 27863
rect 36176 27820 36228 27829
rect 42984 27820 43036 27872
rect 44180 27820 44232 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4804 27659 4856 27668
rect 4804 27625 4813 27659
rect 4813 27625 4847 27659
rect 4847 27625 4856 27659
rect 4804 27616 4856 27625
rect 5448 27659 5500 27668
rect 5448 27625 5457 27659
rect 5457 27625 5491 27659
rect 5491 27625 5500 27659
rect 5448 27616 5500 27625
rect 5632 27616 5684 27668
rect 5632 27387 5684 27396
rect 5632 27353 5641 27387
rect 5641 27353 5675 27387
rect 5675 27353 5684 27387
rect 5632 27344 5684 27353
rect 6552 27616 6604 27668
rect 8300 27616 8352 27668
rect 8852 27616 8904 27668
rect 9128 27616 9180 27668
rect 11060 27616 11112 27668
rect 12808 27616 12860 27668
rect 13452 27616 13504 27668
rect 14280 27616 14332 27668
rect 16028 27659 16080 27668
rect 16028 27625 16037 27659
rect 16037 27625 16071 27659
rect 16071 27625 16080 27659
rect 16028 27616 16080 27625
rect 21548 27616 21600 27668
rect 11336 27480 11388 27532
rect 13728 27480 13780 27532
rect 16672 27480 16724 27532
rect 7012 27455 7064 27464
rect 7012 27421 7021 27455
rect 7021 27421 7055 27455
rect 7055 27421 7064 27455
rect 7012 27412 7064 27421
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 9220 27412 9272 27421
rect 9404 27455 9456 27464
rect 9404 27421 9413 27455
rect 9413 27421 9447 27455
rect 9447 27421 9456 27455
rect 9404 27412 9456 27421
rect 9680 27412 9732 27464
rect 13636 27344 13688 27396
rect 14556 27387 14608 27396
rect 14556 27353 14565 27387
rect 14565 27353 14599 27387
rect 14599 27353 14608 27387
rect 14556 27344 14608 27353
rect 8208 27276 8260 27328
rect 8392 27276 8444 27328
rect 18144 27344 18196 27396
rect 16304 27276 16356 27328
rect 20812 27412 20864 27464
rect 27712 27616 27764 27668
rect 31852 27616 31904 27668
rect 34520 27616 34572 27668
rect 36728 27659 36780 27668
rect 36728 27625 36737 27659
rect 36737 27625 36771 27659
rect 36771 27625 36780 27659
rect 36728 27616 36780 27625
rect 36820 27616 36872 27668
rect 39488 27616 39540 27668
rect 43076 27616 43128 27668
rect 43444 27616 43496 27668
rect 23112 27548 23164 27600
rect 34796 27548 34848 27600
rect 39304 27591 39356 27600
rect 39304 27557 39313 27591
rect 39313 27557 39347 27591
rect 39347 27557 39356 27591
rect 39304 27548 39356 27557
rect 39764 27548 39816 27600
rect 24676 27480 24728 27532
rect 26976 27480 27028 27532
rect 34612 27480 34664 27532
rect 42800 27480 42852 27532
rect 22192 27412 22244 27464
rect 22652 27412 22704 27464
rect 24584 27412 24636 27464
rect 25504 27412 25556 27464
rect 26424 27455 26476 27464
rect 26424 27421 26433 27455
rect 26433 27421 26467 27455
rect 26467 27421 26476 27455
rect 26424 27412 26476 27421
rect 34336 27455 34388 27464
rect 34336 27421 34345 27455
rect 34345 27421 34379 27455
rect 34379 27421 34388 27455
rect 34336 27412 34388 27421
rect 19340 27276 19392 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 25044 27276 25096 27328
rect 27712 27344 27764 27396
rect 35256 27455 35308 27464
rect 35256 27421 35265 27455
rect 35265 27421 35299 27455
rect 35299 27421 35308 27455
rect 35256 27412 35308 27421
rect 35440 27412 35492 27464
rect 35900 27412 35952 27464
rect 36084 27412 36136 27464
rect 36912 27412 36964 27464
rect 38844 27344 38896 27396
rect 40316 27455 40368 27464
rect 40316 27421 40325 27455
rect 40325 27421 40359 27455
rect 40359 27421 40368 27455
rect 40316 27412 40368 27421
rect 39764 27344 39816 27396
rect 28448 27319 28500 27328
rect 28448 27285 28457 27319
rect 28457 27285 28491 27319
rect 28491 27285 28500 27319
rect 28448 27276 28500 27285
rect 30656 27276 30708 27328
rect 34704 27276 34756 27328
rect 36360 27276 36412 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8484 27072 8536 27124
rect 8576 27072 8628 27124
rect 9036 27072 9088 27124
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 13728 27072 13780 27124
rect 14556 27072 14608 27124
rect 22192 27072 22244 27124
rect 23112 27072 23164 27124
rect 6920 27004 6972 27056
rect 7104 27004 7156 27056
rect 5540 26936 5592 26988
rect 8208 26936 8260 26988
rect 8116 26843 8168 26852
rect 8116 26809 8125 26843
rect 8125 26809 8159 26843
rect 8159 26809 8168 26843
rect 8116 26800 8168 26809
rect 8852 26979 8904 26988
rect 8852 26945 8861 26979
rect 8861 26945 8895 26979
rect 8895 26945 8904 26979
rect 8852 26936 8904 26945
rect 14740 27047 14792 27056
rect 14740 27013 14749 27047
rect 14749 27013 14783 27047
rect 14783 27013 14792 27047
rect 14740 27004 14792 27013
rect 9220 26936 9272 26988
rect 14096 26936 14148 26988
rect 14924 26936 14976 26988
rect 20628 27004 20680 27056
rect 9404 26868 9456 26920
rect 12072 26911 12124 26920
rect 12072 26877 12081 26911
rect 12081 26877 12115 26911
rect 12115 26877 12124 26911
rect 12072 26868 12124 26877
rect 20628 26868 20680 26920
rect 22468 27004 22520 27056
rect 20812 26936 20864 26988
rect 22652 26936 22704 26988
rect 22836 26911 22888 26920
rect 22836 26877 22845 26911
rect 22845 26877 22879 26911
rect 22879 26877 22888 26911
rect 22836 26868 22888 26877
rect 24400 27072 24452 27124
rect 25780 27115 25832 27124
rect 25780 27081 25789 27115
rect 25789 27081 25823 27115
rect 25823 27081 25832 27115
rect 25780 27072 25832 27081
rect 26424 27072 26476 27124
rect 28448 27072 28500 27124
rect 24768 27004 24820 27056
rect 29276 27072 29328 27124
rect 30104 27072 30156 27124
rect 34336 27072 34388 27124
rect 35256 27115 35308 27124
rect 35256 27081 35265 27115
rect 35265 27081 35299 27115
rect 35299 27081 35308 27115
rect 35256 27072 35308 27081
rect 36820 27072 36872 27124
rect 43168 27072 43220 27124
rect 23480 26868 23532 26920
rect 21364 26800 21416 26852
rect 24124 26800 24176 26852
rect 27436 26911 27488 26920
rect 27436 26877 27445 26911
rect 27445 26877 27479 26911
rect 27479 26877 27488 26911
rect 27436 26868 27488 26877
rect 27528 26911 27580 26920
rect 27528 26877 27537 26911
rect 27537 26877 27571 26911
rect 27571 26877 27580 26911
rect 27528 26868 27580 26877
rect 29000 26936 29052 26988
rect 30656 26936 30708 26988
rect 28816 26868 28868 26920
rect 29644 26911 29696 26920
rect 29644 26877 29653 26911
rect 29653 26877 29687 26911
rect 29687 26877 29696 26911
rect 29644 26868 29696 26877
rect 34428 26868 34480 26920
rect 34796 26936 34848 26988
rect 35624 27004 35676 27056
rect 36360 27004 36412 27056
rect 28632 26800 28684 26852
rect 35164 26800 35216 26852
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 17960 26775 18012 26784
rect 17960 26741 17969 26775
rect 17969 26741 18003 26775
rect 18003 26741 18012 26775
rect 17960 26732 18012 26741
rect 26148 26732 26200 26784
rect 35440 26868 35492 26920
rect 35808 26979 35860 26988
rect 35808 26945 35817 26979
rect 35817 26945 35851 26979
rect 35851 26945 35860 26979
rect 35808 26936 35860 26945
rect 35900 26979 35952 26988
rect 35900 26945 35909 26979
rect 35909 26945 35943 26979
rect 35943 26945 35952 26979
rect 35900 26936 35952 26945
rect 36176 26979 36228 26988
rect 36176 26945 36185 26979
rect 36185 26945 36219 26979
rect 36219 26945 36228 26979
rect 36176 26936 36228 26945
rect 42432 26979 42484 26988
rect 42432 26945 42441 26979
rect 42441 26945 42475 26979
rect 42475 26945 42484 26979
rect 42432 26936 42484 26945
rect 42708 26979 42760 26988
rect 42708 26945 42717 26979
rect 42717 26945 42751 26979
rect 42751 26945 42760 26979
rect 42708 26936 42760 26945
rect 42984 26936 43036 26988
rect 43996 26936 44048 26988
rect 43536 26911 43588 26920
rect 43536 26877 43545 26911
rect 43545 26877 43579 26911
rect 43579 26877 43588 26911
rect 43536 26868 43588 26877
rect 38108 26732 38160 26784
rect 42892 26732 42944 26784
rect 43076 26775 43128 26784
rect 43076 26741 43085 26775
rect 43085 26741 43119 26775
rect 43119 26741 43128 26775
rect 43076 26732 43128 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 12072 26528 12124 26580
rect 13084 26528 13136 26580
rect 18052 26528 18104 26580
rect 18420 26528 18472 26580
rect 27436 26528 27488 26580
rect 28816 26571 28868 26580
rect 28816 26537 28825 26571
rect 28825 26537 28859 26571
rect 28859 26537 28868 26571
rect 28816 26528 28868 26537
rect 29000 26528 29052 26580
rect 30012 26571 30064 26580
rect 30012 26537 30021 26571
rect 30021 26537 30055 26571
rect 30055 26537 30064 26571
rect 30012 26528 30064 26537
rect 34704 26528 34756 26580
rect 35348 26528 35400 26580
rect 35808 26528 35860 26580
rect 23020 26460 23072 26512
rect 11244 26392 11296 26444
rect 12440 26392 12492 26444
rect 17132 26392 17184 26444
rect 20536 26435 20588 26444
rect 20536 26401 20545 26435
rect 20545 26401 20579 26435
rect 20579 26401 20588 26435
rect 20536 26392 20588 26401
rect 21364 26435 21416 26444
rect 21364 26401 21373 26435
rect 21373 26401 21407 26435
rect 21407 26401 21416 26435
rect 21364 26392 21416 26401
rect 21548 26435 21600 26444
rect 21548 26401 21557 26435
rect 21557 26401 21591 26435
rect 21591 26401 21600 26435
rect 21548 26392 21600 26401
rect 26976 26460 27028 26512
rect 28632 26392 28684 26444
rect 10876 26324 10928 26376
rect 11796 26256 11848 26308
rect 15292 26256 15344 26308
rect 16304 26324 16356 26376
rect 16672 26324 16724 26376
rect 18144 26324 18196 26376
rect 19248 26324 19300 26376
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 24124 26324 24176 26376
rect 29000 26367 29052 26376
rect 29000 26333 29009 26367
rect 29009 26333 29043 26367
rect 29043 26333 29052 26367
rect 29000 26324 29052 26333
rect 10232 26188 10284 26240
rect 17040 26299 17092 26308
rect 17040 26265 17049 26299
rect 17049 26265 17083 26299
rect 17083 26265 17092 26299
rect 17040 26256 17092 26265
rect 20260 26256 20312 26308
rect 21640 26256 21692 26308
rect 24676 26256 24728 26308
rect 19432 26188 19484 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 27712 26256 27764 26308
rect 26148 26231 26200 26240
rect 26148 26197 26157 26231
rect 26157 26197 26191 26231
rect 26191 26197 26200 26231
rect 26148 26188 26200 26197
rect 29276 26367 29328 26376
rect 29276 26333 29285 26367
rect 29285 26333 29319 26367
rect 29319 26333 29328 26367
rect 29276 26324 29328 26333
rect 29460 26392 29512 26444
rect 33416 26503 33468 26512
rect 33416 26469 33425 26503
rect 33425 26469 33459 26503
rect 33459 26469 33468 26503
rect 33416 26460 33468 26469
rect 32220 26392 32272 26444
rect 33140 26435 33192 26444
rect 33140 26401 33149 26435
rect 33149 26401 33183 26435
rect 33183 26401 33192 26435
rect 33140 26392 33192 26401
rect 33324 26324 33376 26376
rect 29552 26299 29604 26308
rect 29552 26265 29561 26299
rect 29561 26265 29595 26299
rect 29595 26265 29604 26299
rect 29552 26256 29604 26265
rect 30840 26299 30892 26308
rect 30840 26265 30849 26299
rect 30849 26265 30883 26299
rect 30883 26265 30892 26299
rect 30840 26256 30892 26265
rect 31852 26256 31904 26308
rect 34612 26324 34664 26376
rect 39396 26392 39448 26444
rect 40500 26392 40552 26444
rect 40960 26392 41012 26444
rect 42616 26528 42668 26580
rect 42984 26528 43036 26580
rect 43996 26528 44048 26580
rect 36912 26324 36964 26376
rect 37280 26324 37332 26376
rect 39948 26324 40000 26376
rect 35348 26299 35400 26308
rect 35348 26265 35357 26299
rect 35357 26265 35391 26299
rect 35391 26265 35400 26299
rect 35348 26256 35400 26265
rect 29460 26188 29512 26240
rect 32128 26188 32180 26240
rect 33600 26231 33652 26240
rect 33600 26197 33609 26231
rect 33609 26197 33643 26231
rect 33643 26197 33652 26231
rect 33600 26188 33652 26197
rect 33968 26231 34020 26240
rect 33968 26197 33977 26231
rect 33977 26197 34011 26231
rect 34011 26197 34020 26231
rect 33968 26188 34020 26197
rect 34152 26231 34204 26240
rect 34152 26197 34161 26231
rect 34161 26197 34195 26231
rect 34195 26197 34204 26231
rect 34152 26188 34204 26197
rect 34796 26188 34848 26240
rect 37740 26299 37792 26308
rect 37740 26265 37749 26299
rect 37749 26265 37783 26299
rect 37783 26265 37792 26299
rect 37740 26256 37792 26265
rect 39488 26299 39540 26308
rect 39488 26265 39497 26299
rect 39497 26265 39531 26299
rect 39531 26265 39540 26299
rect 39488 26256 39540 26265
rect 39580 26256 39632 26308
rect 38752 26188 38804 26240
rect 40224 26367 40276 26376
rect 40224 26333 40233 26367
rect 40233 26333 40267 26367
rect 40267 26333 40276 26367
rect 40224 26324 40276 26333
rect 40868 26367 40920 26376
rect 40868 26333 40877 26367
rect 40877 26333 40911 26367
rect 40911 26333 40920 26367
rect 40868 26324 40920 26333
rect 41420 26367 41472 26376
rect 41420 26333 41429 26367
rect 41429 26333 41463 26367
rect 41463 26333 41472 26367
rect 41420 26324 41472 26333
rect 41512 26324 41564 26376
rect 42800 26392 42852 26444
rect 40592 26299 40644 26308
rect 40592 26265 40601 26299
rect 40601 26265 40635 26299
rect 40635 26265 40644 26299
rect 40592 26256 40644 26265
rect 41788 26299 41840 26308
rect 41144 26188 41196 26240
rect 41788 26265 41797 26299
rect 41797 26265 41831 26299
rect 41831 26265 41840 26299
rect 41788 26256 41840 26265
rect 42524 26256 42576 26308
rect 42892 26367 42944 26376
rect 42892 26333 42901 26367
rect 42901 26333 42935 26367
rect 42935 26333 42944 26367
rect 42892 26324 42944 26333
rect 43260 26299 43312 26308
rect 43260 26265 43269 26299
rect 43269 26265 43303 26299
rect 43303 26265 43312 26299
rect 43260 26256 43312 26265
rect 43720 26256 43772 26308
rect 42708 26188 42760 26240
rect 43352 26188 43404 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 7104 25984 7156 26036
rect 12440 25984 12492 26036
rect 9956 25916 10008 25968
rect 11612 25916 11664 25968
rect 17040 25984 17092 26036
rect 12992 25891 13044 25900
rect 12992 25857 13010 25891
rect 13010 25857 13044 25891
rect 12992 25848 13044 25857
rect 7748 25823 7800 25832
rect 7748 25789 7757 25823
rect 7757 25789 7791 25823
rect 7791 25789 7800 25823
rect 7748 25780 7800 25789
rect 9680 25823 9732 25832
rect 9680 25789 9689 25823
rect 9689 25789 9723 25823
rect 9723 25789 9732 25823
rect 9680 25780 9732 25789
rect 10876 25780 10928 25832
rect 13452 25848 13504 25900
rect 16764 25848 16816 25900
rect 18420 25984 18472 26036
rect 19340 25984 19392 26036
rect 19432 25984 19484 26036
rect 18696 25848 18748 25900
rect 16212 25780 16264 25832
rect 18604 25780 18656 25832
rect 19340 25848 19392 25900
rect 21364 25984 21416 26036
rect 21640 26027 21692 26036
rect 21640 25993 21649 26027
rect 21649 25993 21683 26027
rect 21683 25993 21692 26027
rect 21640 25984 21692 25993
rect 23020 25984 23072 26036
rect 24032 25984 24084 26036
rect 26148 25984 26200 26036
rect 29644 26027 29696 26036
rect 29644 25993 29653 26027
rect 29653 25993 29687 26027
rect 29687 25993 29696 26027
rect 29644 25984 29696 25993
rect 30840 25984 30892 26036
rect 27712 25916 27764 25968
rect 32128 25916 32180 25968
rect 33140 25984 33192 26036
rect 37740 25984 37792 26036
rect 39396 25984 39448 26036
rect 39580 25984 39632 26036
rect 39948 25984 40000 26036
rect 40224 26027 40276 26036
rect 40224 25993 40233 26027
rect 40233 25993 40267 26027
rect 40267 25993 40276 26027
rect 40224 25984 40276 25993
rect 41420 25984 41472 26036
rect 42432 26027 42484 26036
rect 42432 25993 42441 26027
rect 42441 25993 42475 26027
rect 42475 25993 42484 26027
rect 42432 25984 42484 25993
rect 23572 25891 23624 25900
rect 23572 25857 23581 25891
rect 23581 25857 23615 25891
rect 23615 25857 23624 25891
rect 23572 25848 23624 25857
rect 26608 25891 26660 25900
rect 26608 25857 26617 25891
rect 26617 25857 26651 25891
rect 26651 25857 26660 25891
rect 26608 25848 26660 25857
rect 29276 25848 29328 25900
rect 31576 25891 31628 25900
rect 31576 25857 31585 25891
rect 31585 25857 31619 25891
rect 31619 25857 31628 25891
rect 31576 25848 31628 25857
rect 32220 25891 32272 25900
rect 32220 25857 32229 25891
rect 32229 25857 32263 25891
rect 32263 25857 32272 25891
rect 32220 25848 32272 25857
rect 19432 25780 19484 25832
rect 22284 25823 22336 25832
rect 22284 25789 22293 25823
rect 22293 25789 22327 25823
rect 22327 25789 22336 25823
rect 22284 25780 22336 25789
rect 22468 25823 22520 25832
rect 22468 25789 22477 25823
rect 22477 25789 22511 25823
rect 22511 25789 22520 25823
rect 22468 25780 22520 25789
rect 22836 25823 22888 25832
rect 22836 25789 22845 25823
rect 22845 25789 22879 25823
rect 22879 25789 22888 25823
rect 22836 25780 22888 25789
rect 24768 25823 24820 25832
rect 24768 25789 24777 25823
rect 24777 25789 24811 25823
rect 24811 25789 24820 25823
rect 24768 25780 24820 25789
rect 26976 25823 27028 25832
rect 26976 25789 26985 25823
rect 26985 25789 27019 25823
rect 27019 25789 27028 25823
rect 26976 25780 27028 25789
rect 31484 25823 31536 25832
rect 31484 25789 31493 25823
rect 31493 25789 31527 25823
rect 31527 25789 31536 25823
rect 31484 25780 31536 25789
rect 32496 25848 32548 25900
rect 32680 25848 32732 25900
rect 33968 25891 34020 25900
rect 33968 25857 33977 25891
rect 33977 25857 34011 25891
rect 34011 25857 34020 25891
rect 33968 25848 34020 25857
rect 34152 25848 34204 25900
rect 39488 25848 39540 25900
rect 40868 25916 40920 25968
rect 41144 25959 41196 25968
rect 41144 25925 41153 25959
rect 41153 25925 41187 25959
rect 41187 25925 41196 25959
rect 41144 25916 41196 25925
rect 41512 25916 41564 25968
rect 33048 25780 33100 25832
rect 35348 25780 35400 25832
rect 38384 25823 38436 25832
rect 38384 25789 38393 25823
rect 38393 25789 38427 25823
rect 38427 25789 38436 25823
rect 38384 25780 38436 25789
rect 40500 25848 40552 25900
rect 40408 25780 40460 25832
rect 43168 25984 43220 26036
rect 43260 26027 43312 26036
rect 43260 25993 43269 26027
rect 43269 25993 43303 26027
rect 43303 25993 43312 26027
rect 43260 25984 43312 25993
rect 42064 25780 42116 25832
rect 42984 25891 43036 25900
rect 42984 25857 42993 25891
rect 42993 25857 43027 25891
rect 43027 25857 43036 25891
rect 42984 25848 43036 25857
rect 43076 25848 43128 25900
rect 44180 25848 44232 25900
rect 8208 25644 8260 25696
rect 9312 25644 9364 25696
rect 17960 25712 18012 25764
rect 29460 25712 29512 25764
rect 32128 25712 32180 25764
rect 42524 25712 42576 25764
rect 42892 25712 42944 25764
rect 43352 25780 43404 25832
rect 43168 25712 43220 25764
rect 43904 25712 43956 25764
rect 10324 25644 10376 25696
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 13360 25687 13412 25696
rect 13360 25653 13369 25687
rect 13369 25653 13403 25687
rect 13403 25653 13412 25687
rect 13360 25644 13412 25653
rect 15200 25644 15252 25696
rect 16120 25687 16172 25696
rect 16120 25653 16129 25687
rect 16129 25653 16163 25687
rect 16163 25653 16172 25687
rect 16120 25644 16172 25653
rect 19524 25644 19576 25696
rect 23756 25687 23808 25696
rect 23756 25653 23765 25687
rect 23765 25653 23799 25687
rect 23799 25653 23808 25687
rect 23756 25644 23808 25653
rect 29000 25644 29052 25696
rect 29552 25644 29604 25696
rect 29736 25644 29788 25696
rect 32404 25644 32456 25696
rect 38660 25687 38712 25696
rect 38660 25653 38669 25687
rect 38669 25653 38703 25687
rect 38703 25653 38712 25687
rect 38660 25644 38712 25653
rect 39028 25644 39080 25696
rect 42800 25644 42852 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7748 25440 7800 25492
rect 9680 25440 9732 25492
rect 11244 25440 11296 25492
rect 11796 25440 11848 25492
rect 12992 25440 13044 25492
rect 13360 25440 13412 25492
rect 15292 25440 15344 25492
rect 16120 25440 16172 25492
rect 16672 25440 16724 25492
rect 17040 25483 17092 25492
rect 17040 25449 17049 25483
rect 17049 25449 17083 25483
rect 17083 25449 17092 25483
rect 17040 25440 17092 25449
rect 18328 25440 18380 25492
rect 19524 25440 19576 25492
rect 20260 25440 20312 25492
rect 22836 25440 22888 25492
rect 26608 25440 26660 25492
rect 29552 25483 29604 25492
rect 29552 25449 29561 25483
rect 29561 25449 29595 25483
rect 29595 25449 29604 25483
rect 29552 25440 29604 25449
rect 31484 25440 31536 25492
rect 31576 25440 31628 25492
rect 31944 25440 31996 25492
rect 32680 25440 32732 25492
rect 33416 25440 33468 25492
rect 10232 25372 10284 25424
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 14924 25304 14976 25356
rect 17132 25304 17184 25356
rect 10876 25168 10928 25220
rect 11612 25168 11664 25220
rect 13636 25143 13688 25152
rect 13636 25109 13645 25143
rect 13645 25109 13679 25143
rect 13679 25109 13688 25143
rect 13636 25100 13688 25109
rect 15200 25236 15252 25288
rect 19432 25236 19484 25288
rect 23756 25304 23808 25356
rect 24124 25347 24176 25356
rect 24124 25313 24133 25347
rect 24133 25313 24167 25347
rect 24167 25313 24176 25347
rect 24124 25304 24176 25313
rect 24768 25304 24820 25356
rect 27528 25304 27580 25356
rect 29092 25347 29144 25356
rect 29092 25313 29101 25347
rect 29101 25313 29135 25347
rect 29135 25313 29144 25347
rect 29092 25304 29144 25313
rect 32128 25304 32180 25356
rect 33600 25372 33652 25424
rect 33416 25304 33468 25356
rect 14832 25168 14884 25220
rect 17592 25211 17644 25220
rect 17592 25177 17601 25211
rect 17601 25177 17635 25211
rect 17635 25177 17644 25211
rect 17592 25168 17644 25177
rect 18052 25168 18104 25220
rect 18144 25168 18196 25220
rect 24676 25168 24728 25220
rect 24952 25168 25004 25220
rect 22376 25143 22428 25152
rect 22376 25109 22385 25143
rect 22385 25109 22419 25143
rect 22419 25109 22428 25143
rect 31944 25279 31996 25288
rect 29828 25168 29880 25220
rect 31944 25245 31953 25279
rect 31953 25245 31987 25279
rect 31987 25245 31996 25279
rect 31944 25236 31996 25245
rect 22376 25100 22428 25109
rect 27160 25143 27212 25152
rect 27160 25109 27169 25143
rect 27169 25109 27203 25143
rect 27203 25109 27212 25143
rect 27160 25100 27212 25109
rect 29000 25100 29052 25152
rect 32220 25236 32272 25288
rect 33324 25279 33376 25288
rect 33324 25245 33333 25279
rect 33333 25245 33367 25279
rect 33367 25245 33376 25279
rect 33324 25236 33376 25245
rect 36268 25440 36320 25492
rect 38384 25440 38436 25492
rect 38660 25440 38712 25492
rect 37280 25304 37332 25356
rect 38476 25304 38528 25356
rect 34060 25279 34112 25288
rect 34060 25245 34069 25279
rect 34069 25245 34103 25279
rect 34103 25245 34112 25279
rect 34060 25236 34112 25245
rect 36912 25236 36964 25288
rect 43536 25440 43588 25492
rect 42064 25372 42116 25424
rect 42800 25236 42852 25288
rect 42892 25279 42944 25288
rect 42892 25245 42901 25279
rect 42901 25245 42935 25279
rect 42935 25245 42944 25279
rect 42892 25236 42944 25245
rect 31852 25100 31904 25152
rect 32404 25143 32456 25152
rect 32404 25109 32413 25143
rect 32413 25109 32447 25143
rect 32447 25109 32456 25143
rect 33876 25211 33928 25220
rect 33876 25177 33885 25211
rect 33885 25177 33919 25211
rect 33919 25177 33928 25211
rect 33876 25168 33928 25177
rect 33968 25211 34020 25220
rect 33968 25177 33977 25211
rect 33977 25177 34011 25211
rect 34011 25177 34020 25211
rect 33968 25168 34020 25177
rect 32404 25100 32456 25109
rect 33140 25100 33192 25152
rect 42984 25168 43036 25220
rect 43260 25168 43312 25220
rect 34796 25143 34848 25152
rect 34796 25109 34805 25143
rect 34805 25109 34839 25143
rect 34839 25109 34848 25143
rect 34796 25100 34848 25109
rect 34980 25100 35032 25152
rect 42340 25143 42392 25152
rect 42340 25109 42349 25143
rect 42349 25109 42383 25143
rect 42383 25109 42392 25143
rect 42340 25100 42392 25109
rect 42800 25100 42852 25152
rect 44364 25100 44416 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 10876 24939 10928 24948
rect 10876 24905 10885 24939
rect 10885 24905 10919 24939
rect 10919 24905 10928 24939
rect 10876 24896 10928 24905
rect 11612 24896 11664 24948
rect 13452 24896 13504 24948
rect 14832 24896 14884 24948
rect 16212 24939 16264 24948
rect 16212 24905 16221 24939
rect 16221 24905 16255 24939
rect 16255 24905 16264 24939
rect 16212 24896 16264 24905
rect 16764 24939 16816 24948
rect 16764 24905 16773 24939
rect 16773 24905 16807 24939
rect 16807 24905 16816 24939
rect 16764 24896 16816 24905
rect 17040 24896 17092 24948
rect 17592 24896 17644 24948
rect 18328 24939 18380 24948
rect 18328 24905 18337 24939
rect 18337 24905 18371 24939
rect 18371 24905 18380 24939
rect 18328 24896 18380 24905
rect 19340 24896 19392 24948
rect 20260 24939 20312 24948
rect 20260 24905 20269 24939
rect 20269 24905 20303 24939
rect 20303 24905 20312 24939
rect 20260 24896 20312 24905
rect 22376 24896 22428 24948
rect 23572 24896 23624 24948
rect 11520 24760 11572 24812
rect 11888 24760 11940 24812
rect 13728 24828 13780 24880
rect 24952 24896 25004 24948
rect 14924 24760 14976 24812
rect 15108 24803 15160 24812
rect 15108 24769 15142 24803
rect 15142 24769 15160 24803
rect 15108 24760 15160 24769
rect 15844 24760 15896 24812
rect 26976 24896 27028 24948
rect 29092 24896 29144 24948
rect 29276 24896 29328 24948
rect 29920 24896 29972 24948
rect 31944 24896 31996 24948
rect 13636 24692 13688 24744
rect 17224 24735 17276 24744
rect 17224 24701 17233 24735
rect 17233 24701 17267 24735
rect 17267 24701 17276 24735
rect 17224 24692 17276 24701
rect 22008 24760 22060 24812
rect 24676 24803 24728 24812
rect 24676 24769 24685 24803
rect 24685 24769 24719 24803
rect 24719 24769 24728 24803
rect 24676 24760 24728 24769
rect 28724 24803 28776 24812
rect 28724 24769 28733 24803
rect 28733 24769 28767 24803
rect 28767 24769 28776 24803
rect 28724 24760 28776 24769
rect 29276 24760 29328 24812
rect 29828 24803 29880 24812
rect 18420 24735 18472 24744
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 20352 24735 20404 24744
rect 20352 24701 20361 24735
rect 20361 24701 20395 24735
rect 20395 24701 20404 24735
rect 20352 24692 20404 24701
rect 20536 24735 20588 24744
rect 20536 24701 20545 24735
rect 20545 24701 20579 24735
rect 20579 24701 20588 24735
rect 20536 24692 20588 24701
rect 21916 24735 21968 24744
rect 21916 24701 21925 24735
rect 21925 24701 21959 24735
rect 21959 24701 21968 24735
rect 21916 24692 21968 24701
rect 24768 24692 24820 24744
rect 29828 24769 29837 24803
rect 29837 24769 29871 24803
rect 29871 24769 29880 24803
rect 29828 24760 29880 24769
rect 31852 24828 31904 24880
rect 32220 24828 32272 24880
rect 33324 24896 33376 24948
rect 33876 24896 33928 24948
rect 33968 24896 34020 24948
rect 39488 24896 39540 24948
rect 32128 24803 32180 24812
rect 24952 24556 25004 24608
rect 26976 24624 27028 24676
rect 26700 24599 26752 24608
rect 26700 24565 26709 24599
rect 26709 24565 26743 24599
rect 26743 24565 26752 24599
rect 29736 24735 29788 24744
rect 29736 24701 29745 24735
rect 29745 24701 29779 24735
rect 29779 24701 29788 24735
rect 29736 24692 29788 24701
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 34060 24828 34112 24880
rect 35440 24828 35492 24880
rect 42708 24828 42760 24880
rect 42800 24871 42852 24880
rect 42800 24837 42825 24871
rect 42825 24837 42852 24871
rect 42800 24828 42852 24837
rect 26700 24556 26752 24565
rect 29460 24556 29512 24608
rect 32680 24624 32732 24676
rect 33416 24803 33468 24812
rect 33416 24769 33425 24803
rect 33425 24769 33459 24803
rect 33459 24769 33468 24803
rect 33416 24760 33468 24769
rect 34980 24803 35032 24812
rect 34980 24769 34989 24803
rect 34989 24769 35023 24803
rect 35023 24769 35032 24803
rect 34980 24760 35032 24769
rect 33232 24735 33284 24744
rect 33232 24701 33241 24735
rect 33241 24701 33275 24735
rect 33275 24701 33284 24735
rect 33232 24692 33284 24701
rect 33600 24735 33652 24744
rect 33600 24701 33609 24735
rect 33609 24701 33643 24735
rect 33643 24701 33652 24735
rect 33600 24692 33652 24701
rect 38476 24692 38528 24744
rect 39120 24803 39172 24812
rect 39120 24769 39129 24803
rect 39129 24769 39163 24803
rect 39163 24769 39172 24803
rect 39120 24760 39172 24769
rect 40040 24760 40092 24812
rect 40684 24760 40736 24812
rect 40776 24803 40828 24812
rect 40776 24769 40785 24803
rect 40785 24769 40819 24803
rect 40819 24769 40828 24803
rect 40776 24760 40828 24769
rect 39396 24692 39448 24744
rect 41604 24692 41656 24744
rect 42340 24760 42392 24812
rect 43260 24896 43312 24948
rect 43076 24803 43128 24812
rect 43076 24769 43085 24803
rect 43085 24769 43119 24803
rect 43119 24769 43128 24803
rect 43076 24760 43128 24769
rect 37740 24556 37792 24608
rect 38752 24556 38804 24608
rect 43720 24624 43772 24676
rect 40132 24556 40184 24608
rect 41696 24599 41748 24608
rect 41696 24565 41705 24599
rect 41705 24565 41739 24599
rect 41739 24565 41748 24599
rect 41696 24556 41748 24565
rect 43168 24556 43220 24608
rect 44548 24599 44600 24608
rect 44548 24565 44557 24599
rect 44557 24565 44591 24599
rect 44591 24565 44600 24599
rect 44548 24556 44600 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8024 24352 8076 24404
rect 11060 24352 11112 24404
rect 15108 24352 15160 24404
rect 15844 24352 15896 24404
rect 16764 24352 16816 24404
rect 10968 24284 11020 24336
rect 14280 24284 14332 24336
rect 11244 24216 11296 24268
rect 12440 24216 12492 24268
rect 12808 24216 12860 24268
rect 18696 24352 18748 24404
rect 24676 24352 24728 24404
rect 29276 24395 29328 24404
rect 29276 24361 29285 24395
rect 29285 24361 29319 24395
rect 29319 24361 29328 24395
rect 29276 24352 29328 24361
rect 29736 24395 29788 24404
rect 29736 24361 29745 24395
rect 29745 24361 29779 24395
rect 29779 24361 29788 24395
rect 29736 24352 29788 24361
rect 32128 24352 32180 24404
rect 32680 24352 32732 24404
rect 37740 24352 37792 24404
rect 39120 24395 39172 24404
rect 39120 24361 39129 24395
rect 39129 24361 39163 24395
rect 39163 24361 39172 24395
rect 39120 24352 39172 24361
rect 41788 24352 41840 24404
rect 42708 24352 42760 24404
rect 44548 24352 44600 24404
rect 22376 24284 22428 24336
rect 27160 24284 27212 24336
rect 31944 24284 31996 24336
rect 32864 24284 32916 24336
rect 40776 24284 40828 24336
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 10968 24148 11020 24200
rect 11060 24148 11112 24200
rect 11796 24191 11848 24200
rect 11796 24157 11805 24191
rect 11805 24157 11839 24191
rect 11839 24157 11848 24191
rect 11796 24148 11848 24157
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 9220 24012 9272 24064
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10232 24055 10284 24064
rect 10232 24021 10241 24055
rect 10241 24021 10275 24055
rect 10275 24021 10284 24055
rect 10232 24012 10284 24021
rect 10600 24055 10652 24064
rect 10600 24021 10609 24055
rect 10609 24021 10643 24055
rect 10643 24021 10652 24055
rect 10600 24012 10652 24021
rect 12624 24080 12676 24132
rect 11888 24055 11940 24064
rect 11888 24021 11897 24055
rect 11897 24021 11931 24055
rect 11931 24021 11940 24055
rect 11888 24012 11940 24021
rect 12440 24055 12492 24064
rect 12440 24021 12449 24055
rect 12449 24021 12483 24055
rect 12483 24021 12492 24055
rect 12440 24012 12492 24021
rect 12532 24055 12584 24064
rect 12532 24021 12541 24055
rect 12541 24021 12575 24055
rect 12575 24021 12584 24055
rect 12532 24012 12584 24021
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 15200 24148 15252 24200
rect 17592 24080 17644 24132
rect 25320 24216 25372 24268
rect 18696 24148 18748 24200
rect 21916 24148 21968 24200
rect 23388 24148 23440 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 20260 24080 20312 24132
rect 26700 24080 26752 24132
rect 27804 24080 27856 24132
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29460 24080 29512 24132
rect 29920 24148 29972 24200
rect 32312 24148 32364 24200
rect 33508 24216 33560 24268
rect 38660 24216 38712 24268
rect 41420 24216 41472 24268
rect 42892 24216 42944 24268
rect 44364 24259 44416 24268
rect 44364 24225 44373 24259
rect 44373 24225 44407 24259
rect 44407 24225 44416 24259
rect 44364 24216 44416 24225
rect 33048 24191 33100 24200
rect 33048 24157 33057 24191
rect 33057 24157 33091 24191
rect 33091 24157 33100 24191
rect 33048 24148 33100 24157
rect 38752 24148 38804 24200
rect 39396 24191 39448 24200
rect 39396 24157 39405 24191
rect 39405 24157 39439 24191
rect 39439 24157 39448 24191
rect 39396 24148 39448 24157
rect 40132 24148 40184 24200
rect 40408 24191 40460 24200
rect 16672 24055 16724 24064
rect 16672 24021 16681 24055
rect 16681 24021 16715 24055
rect 16715 24021 16724 24055
rect 16672 24012 16724 24021
rect 18144 24012 18196 24064
rect 27712 24055 27764 24064
rect 27712 24021 27721 24055
rect 27721 24021 27755 24055
rect 27755 24021 27764 24055
rect 27712 24012 27764 24021
rect 28264 24055 28316 24064
rect 28264 24021 28273 24055
rect 28273 24021 28307 24055
rect 28307 24021 28316 24055
rect 28264 24012 28316 24021
rect 32680 24012 32732 24064
rect 32772 24012 32824 24064
rect 35808 24123 35860 24132
rect 35808 24089 35817 24123
rect 35817 24089 35851 24123
rect 35851 24089 35860 24123
rect 35808 24080 35860 24089
rect 37924 24080 37976 24132
rect 40408 24157 40417 24191
rect 40417 24157 40451 24191
rect 40451 24157 40460 24191
rect 40408 24148 40460 24157
rect 33692 24012 33744 24064
rect 35348 24012 35400 24064
rect 36452 24012 36504 24064
rect 37280 24055 37332 24064
rect 37280 24021 37289 24055
rect 37289 24021 37323 24055
rect 37323 24021 37332 24055
rect 37280 24012 37332 24021
rect 39212 24012 39264 24064
rect 40040 24055 40092 24064
rect 40040 24021 40067 24055
rect 40067 24021 40092 24055
rect 40040 24012 40092 24021
rect 42616 24080 42668 24132
rect 43720 24080 43772 24132
rect 42064 24012 42116 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 10416 23808 10468 23860
rect 10692 23808 10744 23860
rect 11060 23808 11112 23860
rect 12072 23808 12124 23860
rect 12532 23808 12584 23860
rect 12624 23851 12676 23860
rect 12624 23817 12633 23851
rect 12633 23817 12667 23851
rect 12667 23817 12676 23851
rect 12624 23808 12676 23817
rect 16764 23808 16816 23860
rect 17224 23808 17276 23860
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 18144 23808 18196 23860
rect 19432 23808 19484 23860
rect 34796 23808 34848 23860
rect 16672 23672 16724 23724
rect 17776 23715 17828 23724
rect 17776 23681 17785 23715
rect 17785 23681 17819 23715
rect 17819 23681 17828 23715
rect 17776 23672 17828 23681
rect 19432 23672 19484 23724
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 11244 23647 11296 23656
rect 11244 23613 11253 23647
rect 11253 23613 11287 23647
rect 11287 23613 11296 23647
rect 11244 23604 11296 23613
rect 11520 23647 11572 23656
rect 11520 23613 11529 23647
rect 11529 23613 11563 23647
rect 11563 23613 11572 23647
rect 11520 23604 11572 23613
rect 12440 23604 12492 23656
rect 12808 23647 12860 23656
rect 12808 23613 12817 23647
rect 12817 23613 12851 23647
rect 12851 23613 12860 23647
rect 12808 23604 12860 23613
rect 13636 23647 13688 23656
rect 13636 23613 13645 23647
rect 13645 23613 13679 23647
rect 13679 23613 13688 23647
rect 13636 23604 13688 23613
rect 14648 23604 14700 23656
rect 20076 23715 20128 23724
rect 20076 23681 20110 23715
rect 20110 23681 20128 23715
rect 20076 23672 20128 23681
rect 22744 23715 22796 23724
rect 22744 23681 22778 23715
rect 22778 23681 22796 23715
rect 22744 23672 22796 23681
rect 21916 23604 21968 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 12072 23536 12124 23588
rect 8576 23468 8628 23520
rect 26516 23783 26568 23792
rect 26516 23749 26525 23783
rect 26525 23749 26559 23783
rect 26559 23749 26568 23783
rect 26516 23740 26568 23749
rect 27344 23740 27396 23792
rect 28540 23740 28592 23792
rect 32680 23740 32732 23792
rect 32772 23740 32824 23792
rect 33232 23740 33284 23792
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27252 23647 27304 23656
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 27344 23604 27396 23656
rect 29368 23647 29420 23656
rect 29368 23613 29377 23647
rect 29377 23613 29411 23647
rect 29411 23613 29420 23647
rect 29368 23604 29420 23613
rect 23388 23468 23440 23520
rect 26240 23511 26292 23520
rect 26240 23477 26249 23511
rect 26249 23477 26283 23511
rect 26283 23477 26292 23511
rect 26240 23468 26292 23477
rect 31944 23536 31996 23588
rect 28816 23511 28868 23520
rect 28816 23477 28825 23511
rect 28825 23477 28859 23511
rect 28859 23477 28868 23511
rect 28816 23468 28868 23477
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32404 23715 32456 23724
rect 32404 23681 32413 23715
rect 32413 23681 32447 23715
rect 32447 23681 32456 23715
rect 32404 23672 32456 23681
rect 33048 23672 33100 23724
rect 35348 23808 35400 23860
rect 35808 23808 35860 23860
rect 37924 23808 37976 23860
rect 38568 23808 38620 23860
rect 39212 23808 39264 23860
rect 40408 23808 40460 23860
rect 40684 23808 40736 23860
rect 41604 23808 41656 23860
rect 41696 23808 41748 23860
rect 42064 23808 42116 23860
rect 42800 23851 42852 23860
rect 42800 23817 42809 23851
rect 42809 23817 42843 23851
rect 42843 23817 42852 23851
rect 42800 23808 42852 23817
rect 44548 23808 44600 23860
rect 45284 23808 45336 23860
rect 32772 23604 32824 23656
rect 33416 23647 33468 23656
rect 33416 23613 33425 23647
rect 33425 23613 33459 23647
rect 33459 23613 33468 23647
rect 33416 23604 33468 23613
rect 35440 23672 35492 23724
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 36544 23647 36596 23656
rect 36544 23613 36553 23647
rect 36553 23613 36587 23647
rect 36587 23613 36596 23647
rect 36544 23604 36596 23613
rect 37280 23604 37332 23656
rect 38660 23672 38712 23724
rect 41420 23672 41472 23724
rect 42616 23740 42668 23792
rect 41788 23604 41840 23656
rect 40040 23536 40092 23588
rect 36452 23511 36504 23520
rect 36452 23477 36461 23511
rect 36461 23477 36495 23511
rect 36495 23477 36504 23511
rect 36452 23468 36504 23477
rect 38568 23468 38620 23520
rect 41604 23468 41656 23520
rect 43260 23604 43312 23656
rect 44640 23511 44692 23520
rect 44640 23477 44649 23511
rect 44649 23477 44683 23511
rect 44683 23477 44692 23511
rect 44640 23468 44692 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 11520 23264 11572 23316
rect 17776 23264 17828 23316
rect 20076 23264 20128 23316
rect 22376 23307 22428 23316
rect 22376 23273 22385 23307
rect 22385 23273 22419 23307
rect 22419 23273 22428 23307
rect 22376 23264 22428 23273
rect 27252 23264 27304 23316
rect 29000 23264 29052 23316
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 19800 23196 19852 23248
rect 10232 23128 10284 23180
rect 8576 23060 8628 23112
rect 9220 23060 9272 23112
rect 10600 23060 10652 23112
rect 11612 23060 11664 23112
rect 12900 23060 12952 23112
rect 16028 23060 16080 23112
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 19984 23128 20036 23180
rect 16856 23060 16908 23112
rect 18144 23060 18196 23112
rect 8944 22967 8996 22976
rect 8944 22933 8953 22967
rect 8953 22933 8987 22967
rect 8987 22933 8996 22967
rect 8944 22924 8996 22933
rect 14096 22992 14148 23044
rect 14832 22992 14884 23044
rect 14924 23035 14976 23044
rect 14924 23001 14933 23035
rect 14933 23001 14967 23035
rect 14967 23001 14976 23035
rect 14924 22992 14976 23001
rect 17224 22992 17276 23044
rect 17868 22992 17920 23044
rect 16396 22967 16448 22976
rect 16396 22933 16405 22967
rect 16405 22933 16439 22967
rect 16439 22933 16448 22967
rect 16396 22924 16448 22933
rect 19248 22992 19300 23044
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 20260 23103 20312 23112
rect 20260 23069 20269 23103
rect 20269 23069 20303 23103
rect 20303 23069 20312 23103
rect 20260 23060 20312 23069
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 22468 23128 22520 23180
rect 23020 23171 23072 23180
rect 23020 23137 23029 23171
rect 23029 23137 23063 23171
rect 23063 23137 23072 23171
rect 23020 23128 23072 23137
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 25872 23128 25924 23180
rect 28816 23128 28868 23180
rect 22652 23060 22704 23112
rect 23388 23060 23440 23112
rect 24768 23060 24820 23112
rect 26240 23060 26292 23112
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 28264 23060 28316 23112
rect 29092 23103 29144 23112
rect 29092 23069 29101 23103
rect 29101 23069 29135 23103
rect 29135 23069 29144 23103
rect 29092 23060 29144 23069
rect 20812 22924 20864 22976
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 25504 22924 25556 22976
rect 27804 22924 27856 22976
rect 28816 22992 28868 23044
rect 29000 22992 29052 23044
rect 29368 23035 29420 23044
rect 29368 23001 29377 23035
rect 29377 23001 29411 23035
rect 29411 23001 29420 23035
rect 29368 22992 29420 23001
rect 28172 22924 28224 22976
rect 29092 22924 29144 22976
rect 32128 23264 32180 23316
rect 32404 23264 32456 23316
rect 33416 23264 33468 23316
rect 36544 23264 36596 23316
rect 38660 23264 38712 23316
rect 30932 23171 30984 23180
rect 30932 23137 30941 23171
rect 30941 23137 30975 23171
rect 30975 23137 30984 23171
rect 30932 23128 30984 23137
rect 30288 23103 30340 23112
rect 30288 23069 30297 23103
rect 30297 23069 30331 23103
rect 30331 23069 30340 23103
rect 30288 23060 30340 23069
rect 30380 22992 30432 23044
rect 30840 22992 30892 23044
rect 33692 23128 33744 23180
rect 41788 23264 41840 23316
rect 43260 23307 43312 23316
rect 43260 23273 43269 23307
rect 43269 23273 43303 23307
rect 43303 23273 43312 23307
rect 43260 23264 43312 23273
rect 32588 23103 32640 23112
rect 32588 23069 32597 23103
rect 32597 23069 32631 23103
rect 32631 23069 32640 23103
rect 32588 23060 32640 23069
rect 33048 23060 33100 23112
rect 34520 23060 34572 23112
rect 36360 23103 36412 23112
rect 36360 23069 36369 23103
rect 36369 23069 36403 23103
rect 36403 23069 36412 23103
rect 36360 23060 36412 23069
rect 35992 22992 36044 23044
rect 41604 23060 41656 23112
rect 43536 23060 43588 23112
rect 36636 22992 36688 23044
rect 34612 22924 34664 22976
rect 35624 22924 35676 22976
rect 36544 22924 36596 22976
rect 40500 23035 40552 23044
rect 40500 23001 40509 23035
rect 40509 23001 40543 23035
rect 40543 23001 40552 23035
rect 40500 22992 40552 23001
rect 43076 22924 43128 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9772 22763 9824 22772
rect 9772 22729 9781 22763
rect 9781 22729 9815 22763
rect 9815 22729 9824 22763
rect 9772 22720 9824 22729
rect 13636 22720 13688 22772
rect 14924 22720 14976 22772
rect 15660 22763 15712 22772
rect 15660 22729 15669 22763
rect 15669 22729 15703 22763
rect 15703 22729 15712 22763
rect 15660 22720 15712 22729
rect 16396 22720 16448 22772
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 18420 22720 18472 22772
rect 18880 22720 18932 22772
rect 20720 22720 20772 22772
rect 22376 22720 22428 22772
rect 22468 22720 22520 22772
rect 22744 22720 22796 22772
rect 24768 22720 24820 22772
rect 25504 22763 25556 22772
rect 25504 22729 25513 22763
rect 25513 22729 25547 22763
rect 25547 22729 25556 22763
rect 25504 22720 25556 22729
rect 26516 22720 26568 22772
rect 28172 22720 28224 22772
rect 29368 22720 29420 22772
rect 29736 22720 29788 22772
rect 30288 22720 30340 22772
rect 30380 22720 30432 22772
rect 30932 22720 30984 22772
rect 32588 22720 32640 22772
rect 8576 22652 8628 22704
rect 10968 22652 11020 22704
rect 11888 22652 11940 22704
rect 13544 22652 13596 22704
rect 16580 22652 16632 22704
rect 11612 22584 11664 22636
rect 14464 22627 14516 22636
rect 14464 22593 14473 22627
rect 14473 22593 14507 22627
rect 14507 22593 14516 22627
rect 14464 22584 14516 22593
rect 8944 22516 8996 22568
rect 18052 22627 18104 22636
rect 18052 22593 18061 22627
rect 18061 22593 18095 22627
rect 18095 22593 18104 22627
rect 18052 22584 18104 22593
rect 15384 22516 15436 22568
rect 17224 22559 17276 22568
rect 17224 22525 17233 22559
rect 17233 22525 17267 22559
rect 17267 22525 17276 22559
rect 17224 22516 17276 22525
rect 17868 22516 17920 22568
rect 20628 22652 20680 22704
rect 11796 22380 11848 22432
rect 12164 22380 12216 22432
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 18144 22423 18196 22432
rect 18144 22389 18153 22423
rect 18153 22389 18187 22423
rect 18187 22389 18196 22423
rect 18144 22380 18196 22389
rect 18420 22448 18472 22500
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 22468 22559 22520 22568
rect 22468 22525 22477 22559
rect 22477 22525 22511 22559
rect 22511 22525 22520 22559
rect 22468 22516 22520 22525
rect 23020 22516 23072 22568
rect 23112 22559 23164 22568
rect 23112 22525 23121 22559
rect 23121 22525 23155 22559
rect 23155 22525 23164 22559
rect 23112 22516 23164 22525
rect 19984 22380 20036 22432
rect 22376 22448 22428 22500
rect 24124 22584 24176 22636
rect 25320 22584 25372 22636
rect 27804 22584 27856 22636
rect 28172 22584 28224 22636
rect 28908 22584 28960 22636
rect 29184 22584 29236 22636
rect 29276 22584 29328 22636
rect 27528 22516 27580 22568
rect 33048 22652 33100 22704
rect 28540 22448 28592 22500
rect 30840 22448 30892 22500
rect 24308 22423 24360 22432
rect 24308 22389 24317 22423
rect 24317 22389 24351 22423
rect 24351 22389 24360 22423
rect 24308 22380 24360 22389
rect 29644 22380 29696 22432
rect 32128 22559 32180 22568
rect 32128 22525 32137 22559
rect 32137 22525 32171 22559
rect 32171 22525 32180 22559
rect 32128 22516 32180 22525
rect 32772 22516 32824 22568
rect 34612 22652 34664 22704
rect 35348 22695 35400 22704
rect 35348 22661 35357 22695
rect 35357 22661 35391 22695
rect 35391 22661 35400 22695
rect 35348 22652 35400 22661
rect 35624 22652 35676 22704
rect 36360 22720 36412 22772
rect 40500 22720 40552 22772
rect 35440 22516 35492 22568
rect 35624 22559 35676 22568
rect 35624 22525 35633 22559
rect 35633 22525 35667 22559
rect 35667 22525 35676 22559
rect 35624 22516 35676 22525
rect 36084 22627 36136 22636
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 34060 22423 34112 22432
rect 34060 22389 34069 22423
rect 34069 22389 34103 22423
rect 34103 22389 34112 22423
rect 34060 22380 34112 22389
rect 35624 22380 35676 22432
rect 36176 22448 36228 22500
rect 37740 22516 37792 22568
rect 40040 22559 40092 22568
rect 40040 22525 40049 22559
rect 40049 22525 40083 22559
rect 40083 22525 40092 22559
rect 40040 22516 40092 22525
rect 41788 22584 41840 22636
rect 36268 22423 36320 22432
rect 36268 22389 36277 22423
rect 36277 22389 36311 22423
rect 36311 22389 36320 22423
rect 36268 22380 36320 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14832 22176 14884 22228
rect 16580 22176 16632 22228
rect 18052 22176 18104 22228
rect 20536 22176 20588 22228
rect 16856 22040 16908 22092
rect 17408 22040 17460 22092
rect 23112 22040 23164 22092
rect 14648 21972 14700 22024
rect 24768 22108 24820 22160
rect 25320 22176 25372 22228
rect 29092 22219 29144 22228
rect 29092 22185 29101 22219
rect 29101 22185 29135 22219
rect 29135 22185 29144 22219
rect 29092 22176 29144 22185
rect 31944 22176 31996 22228
rect 34152 22176 34204 22228
rect 28172 22108 28224 22160
rect 25872 22083 25924 22092
rect 25872 22049 25881 22083
rect 25881 22049 25915 22083
rect 25915 22049 25924 22083
rect 25872 22040 25924 22049
rect 15752 21904 15804 21956
rect 13084 21836 13136 21888
rect 18144 21972 18196 22024
rect 22376 21972 22428 22024
rect 23204 21972 23256 22024
rect 29368 22108 29420 22160
rect 29644 22083 29696 22092
rect 29644 22049 29653 22083
rect 29653 22049 29687 22083
rect 29687 22049 29696 22083
rect 29644 22040 29696 22049
rect 19064 21904 19116 21956
rect 19248 21836 19300 21888
rect 23664 21836 23716 21888
rect 29276 21972 29328 22024
rect 35992 22176 36044 22228
rect 36268 22219 36320 22228
rect 36268 22185 36298 22219
rect 36298 22185 36320 22219
rect 36268 22176 36320 22185
rect 37740 22219 37792 22228
rect 37740 22185 37749 22219
rect 37749 22185 37783 22219
rect 37783 22185 37792 22219
rect 37740 22176 37792 22185
rect 38200 22040 38252 22092
rect 38752 22040 38804 22092
rect 39764 22040 39816 22092
rect 26148 21947 26200 21956
rect 26148 21913 26157 21947
rect 26157 21913 26191 21947
rect 26191 21913 26200 21947
rect 26148 21904 26200 21913
rect 27712 21904 27764 21956
rect 28540 21904 28592 21956
rect 25136 21836 25188 21888
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 28908 21904 28960 21956
rect 34060 21947 34112 21956
rect 34060 21913 34069 21947
rect 34069 21913 34103 21947
rect 34103 21913 34112 21947
rect 35348 22015 35400 22024
rect 35348 21981 35357 22015
rect 35357 21981 35391 22015
rect 35391 21981 35400 22015
rect 35348 21972 35400 21981
rect 35440 22015 35492 22024
rect 35440 21981 35449 22015
rect 35449 21981 35483 22015
rect 35483 21981 35492 22015
rect 35440 21972 35492 21981
rect 35532 22015 35584 22024
rect 35532 21981 35541 22015
rect 35541 21981 35575 22015
rect 35575 21981 35584 22015
rect 35532 21972 35584 21981
rect 34060 21904 34112 21913
rect 29736 21836 29788 21888
rect 35808 21879 35860 21888
rect 35808 21845 35817 21879
rect 35817 21845 35851 21879
rect 35851 21845 35860 21879
rect 35808 21836 35860 21845
rect 38108 21947 38160 21956
rect 38108 21913 38117 21947
rect 38117 21913 38151 21947
rect 38151 21913 38160 21947
rect 38108 21904 38160 21913
rect 38568 21904 38620 21956
rect 39856 21879 39908 21888
rect 39856 21845 39865 21879
rect 39865 21845 39899 21879
rect 39899 21845 39908 21879
rect 39856 21836 39908 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 14464 21632 14516 21684
rect 13084 21607 13136 21616
rect 13084 21573 13093 21607
rect 13093 21573 13127 21607
rect 13127 21573 13136 21607
rect 13084 21564 13136 21573
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 15752 21675 15804 21684
rect 15752 21641 15761 21675
rect 15761 21641 15795 21675
rect 15795 21641 15804 21675
rect 15752 21632 15804 21641
rect 16580 21632 16632 21684
rect 19064 21675 19116 21684
rect 19064 21641 19073 21675
rect 19073 21641 19107 21675
rect 19107 21641 19116 21675
rect 19064 21632 19116 21641
rect 19248 21632 19300 21684
rect 23204 21675 23256 21684
rect 23204 21641 23213 21675
rect 23213 21641 23247 21675
rect 23247 21641 23256 21675
rect 23204 21632 23256 21641
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 26148 21675 26200 21684
rect 26148 21641 26157 21675
rect 26157 21641 26191 21675
rect 26191 21641 26200 21675
rect 26148 21632 26200 21641
rect 14188 21496 14240 21548
rect 16028 21564 16080 21616
rect 16672 21496 16724 21548
rect 16764 21496 16816 21548
rect 11980 21428 12032 21480
rect 15108 21471 15160 21480
rect 15108 21437 15117 21471
rect 15117 21437 15151 21471
rect 15151 21437 15160 21471
rect 15108 21428 15160 21437
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 17868 21428 17920 21480
rect 18328 21428 18380 21480
rect 21456 21496 21508 21548
rect 19248 21428 19300 21480
rect 19984 21428 20036 21480
rect 13544 21292 13596 21344
rect 17224 21292 17276 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 23388 21471 23440 21480
rect 23388 21437 23397 21471
rect 23397 21437 23431 21471
rect 23431 21437 23440 21471
rect 23388 21428 23440 21437
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 24308 21428 24360 21480
rect 25136 21428 25188 21480
rect 28080 21632 28132 21684
rect 29736 21675 29788 21684
rect 29736 21641 29745 21675
rect 29745 21641 29779 21675
rect 29779 21641 29788 21675
rect 29736 21632 29788 21641
rect 35348 21675 35400 21684
rect 35348 21641 35357 21675
rect 35357 21641 35391 21675
rect 35391 21641 35400 21675
rect 35348 21632 35400 21641
rect 36084 21675 36136 21684
rect 36084 21641 36093 21675
rect 36093 21641 36127 21675
rect 36127 21641 36136 21675
rect 36084 21632 36136 21641
rect 36452 21632 36504 21684
rect 38108 21632 38160 21684
rect 39856 21632 39908 21684
rect 27620 21564 27672 21616
rect 29276 21564 29328 21616
rect 27528 21471 27580 21480
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 29644 21496 29696 21548
rect 35532 21564 35584 21616
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 23296 21292 23348 21344
rect 28908 21360 28960 21412
rect 35716 21539 35768 21548
rect 35716 21505 35725 21539
rect 35725 21505 35759 21539
rect 35759 21505 35768 21539
rect 35716 21496 35768 21505
rect 36084 21496 36136 21548
rect 35532 21471 35584 21480
rect 35532 21437 35541 21471
rect 35541 21437 35575 21471
rect 35575 21437 35584 21471
rect 35532 21428 35584 21437
rect 28080 21335 28132 21344
rect 28080 21301 28089 21335
rect 28089 21301 28123 21335
rect 28123 21301 28132 21335
rect 28080 21292 28132 21301
rect 29000 21292 29052 21344
rect 35440 21360 35492 21412
rect 36452 21539 36504 21548
rect 36452 21505 36461 21539
rect 36461 21505 36495 21539
rect 36495 21505 36504 21539
rect 36452 21496 36504 21505
rect 39396 21471 39448 21480
rect 39396 21437 39405 21471
rect 39405 21437 39439 21471
rect 39439 21437 39448 21471
rect 39396 21428 39448 21437
rect 35716 21292 35768 21344
rect 38844 21292 38896 21344
rect 39488 21292 39540 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 11428 21088 11480 21140
rect 13820 21088 13872 21140
rect 18696 21131 18748 21140
rect 18696 21097 18705 21131
rect 18705 21097 18739 21131
rect 18739 21097 18748 21131
rect 18696 21088 18748 21097
rect 23296 21088 23348 21140
rect 23204 20952 23256 21004
rect 24768 21088 24820 21140
rect 32312 21131 32364 21140
rect 32312 21097 32321 21131
rect 32321 21097 32355 21131
rect 32355 21097 32364 21131
rect 32312 21088 32364 21097
rect 23664 20952 23716 21004
rect 25136 20952 25188 21004
rect 10784 20884 10836 20936
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 14188 20884 14240 20936
rect 17408 20884 17460 20936
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 23388 20884 23440 20936
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 9772 20859 9824 20868
rect 9772 20825 9781 20859
rect 9781 20825 9815 20859
rect 9815 20825 9824 20859
rect 9772 20816 9824 20825
rect 12256 20859 12308 20868
rect 12256 20825 12265 20859
rect 12265 20825 12299 20859
rect 12299 20825 12308 20859
rect 12256 20816 12308 20825
rect 17776 20816 17828 20868
rect 14464 20748 14516 20800
rect 22744 20791 22796 20800
rect 22744 20757 22753 20791
rect 22753 20757 22787 20791
rect 22787 20757 22796 20791
rect 22744 20748 22796 20757
rect 23756 20791 23808 20800
rect 23756 20757 23765 20791
rect 23765 20757 23799 20791
rect 23799 20757 23808 20791
rect 23756 20748 23808 20757
rect 24216 20791 24268 20800
rect 24216 20757 24225 20791
rect 24225 20757 24259 20791
rect 24259 20757 24268 20791
rect 24216 20748 24268 20757
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 32036 20995 32088 21004
rect 32036 20961 32045 20995
rect 32045 20961 32079 20995
rect 32079 20961 32088 20995
rect 32036 20952 32088 20961
rect 39396 21088 39448 21140
rect 39488 20952 39540 21004
rect 32404 20884 32456 20936
rect 35532 20927 35584 20936
rect 35532 20893 35541 20927
rect 35541 20893 35575 20927
rect 35575 20893 35584 20927
rect 35532 20884 35584 20893
rect 35716 20927 35768 20936
rect 35716 20893 35725 20927
rect 35725 20893 35759 20927
rect 35759 20893 35768 20927
rect 35716 20884 35768 20893
rect 36452 20884 36504 20936
rect 38936 20927 38988 20936
rect 38936 20893 38945 20927
rect 38945 20893 38979 20927
rect 38979 20893 38988 20927
rect 38936 20884 38988 20893
rect 25964 20816 26016 20868
rect 27712 20816 27764 20868
rect 35440 20816 35492 20868
rect 28080 20748 28132 20800
rect 38752 20791 38804 20800
rect 38752 20757 38761 20791
rect 38761 20757 38795 20791
rect 38795 20757 38804 20791
rect 38752 20748 38804 20757
rect 39304 20748 39356 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 9772 20544 9824 20596
rect 11428 20544 11480 20596
rect 13820 20544 13872 20596
rect 12072 20476 12124 20528
rect 11244 20340 11296 20392
rect 12256 20340 12308 20392
rect 11888 20272 11940 20324
rect 15936 20544 15988 20596
rect 17776 20587 17828 20596
rect 17776 20553 17785 20587
rect 17785 20553 17819 20587
rect 17819 20553 17828 20587
rect 17776 20544 17828 20553
rect 18052 20544 18104 20596
rect 18696 20544 18748 20596
rect 20720 20544 20772 20596
rect 21272 20544 21324 20596
rect 21456 20544 21508 20596
rect 22744 20544 22796 20596
rect 23756 20544 23808 20596
rect 24216 20544 24268 20596
rect 24676 20544 24728 20596
rect 32036 20544 32088 20596
rect 32496 20544 32548 20596
rect 38752 20544 38804 20596
rect 38844 20544 38896 20596
rect 39488 20544 39540 20596
rect 13084 20340 13136 20392
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 15200 20340 15252 20392
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 19616 20408 19668 20460
rect 20076 20476 20128 20528
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 31300 20408 31352 20460
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 31944 20408 31996 20460
rect 32220 20408 32272 20460
rect 32404 20451 32456 20460
rect 32404 20417 32413 20451
rect 32413 20417 32447 20451
rect 32447 20417 32456 20451
rect 32404 20408 32456 20417
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 35808 20408 35860 20460
rect 36452 20408 36504 20460
rect 38200 20451 38252 20460
rect 38200 20417 38209 20451
rect 38209 20417 38243 20451
rect 38243 20417 38252 20451
rect 38200 20408 38252 20417
rect 17868 20340 17920 20392
rect 18420 20340 18472 20392
rect 19984 20340 20036 20392
rect 21732 20340 21784 20392
rect 17960 20272 18012 20324
rect 18328 20272 18380 20324
rect 22376 20340 22428 20392
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 31760 20272 31812 20324
rect 32772 20340 32824 20392
rect 13544 20204 13596 20256
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15384 20204 15436 20213
rect 32588 20204 32640 20256
rect 36820 20204 36872 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 12072 20000 12124 20052
rect 13452 20000 13504 20052
rect 19432 20000 19484 20052
rect 14096 19932 14148 19984
rect 15108 19975 15160 19984
rect 15108 19941 15117 19975
rect 15117 19941 15151 19975
rect 15151 19941 15160 19975
rect 15108 19932 15160 19941
rect 15476 19864 15528 19916
rect 15936 19864 15988 19916
rect 11980 19796 12032 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 16764 19796 16816 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 19616 19932 19668 19984
rect 19984 19864 20036 19916
rect 21272 19864 21324 19916
rect 22008 19864 22060 19916
rect 21916 19796 21968 19848
rect 29184 20000 29236 20052
rect 29460 20000 29512 20052
rect 25504 19864 25556 19916
rect 29000 19907 29052 19916
rect 29000 19873 29009 19907
rect 29009 19873 29043 19907
rect 29043 19873 29052 19907
rect 29000 19864 29052 19873
rect 29644 19907 29696 19916
rect 29644 19873 29653 19907
rect 29653 19873 29687 19907
rect 29687 19873 29696 19907
rect 29644 19864 29696 19873
rect 26792 19796 26844 19848
rect 28724 19796 28776 19848
rect 31024 19839 31076 19848
rect 31024 19805 31033 19839
rect 31033 19805 31067 19839
rect 31067 19805 31076 19839
rect 31024 19796 31076 19805
rect 31944 20000 31996 20052
rect 32220 20043 32272 20052
rect 32220 20009 32229 20043
rect 32229 20009 32263 20043
rect 32263 20009 32272 20043
rect 32220 20000 32272 20009
rect 32404 20000 32456 20052
rect 31392 19932 31444 19984
rect 31668 19907 31720 19916
rect 31668 19873 31677 19907
rect 31677 19873 31711 19907
rect 31711 19873 31720 19907
rect 31668 19864 31720 19873
rect 32496 19932 32548 19984
rect 35624 20000 35676 20052
rect 38936 20000 38988 20052
rect 35808 19932 35860 19984
rect 34704 19864 34756 19916
rect 35900 19864 35952 19916
rect 31392 19839 31444 19848
rect 31392 19805 31401 19839
rect 31401 19805 31435 19839
rect 31435 19805 31444 19839
rect 31392 19796 31444 19805
rect 10692 19728 10744 19780
rect 11060 19728 11112 19780
rect 12440 19771 12492 19780
rect 12440 19737 12452 19771
rect 12452 19737 12492 19771
rect 12440 19728 12492 19737
rect 15384 19728 15436 19780
rect 16028 19728 16080 19780
rect 11520 19703 11572 19712
rect 11520 19669 11529 19703
rect 11529 19669 11563 19703
rect 11563 19669 11572 19703
rect 11520 19660 11572 19669
rect 12072 19660 12124 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 19984 19660 20036 19712
rect 21548 19703 21600 19712
rect 21548 19669 21557 19703
rect 21557 19669 21591 19703
rect 21591 19669 21600 19703
rect 21548 19660 21600 19669
rect 23940 19728 23992 19780
rect 24400 19728 24452 19780
rect 26976 19728 27028 19780
rect 28908 19728 28960 19780
rect 22468 19660 22520 19712
rect 27160 19660 27212 19712
rect 29000 19660 29052 19712
rect 29736 19660 29788 19712
rect 31300 19728 31352 19780
rect 31944 19796 31996 19848
rect 32312 19839 32364 19848
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32312 19796 32364 19805
rect 32588 19796 32640 19848
rect 35440 19839 35492 19848
rect 35440 19805 35449 19839
rect 35449 19805 35483 19839
rect 35483 19805 35492 19839
rect 35440 19796 35492 19805
rect 35532 19839 35584 19848
rect 35532 19805 35541 19839
rect 35541 19805 35575 19839
rect 35575 19805 35584 19839
rect 35532 19796 35584 19805
rect 34888 19728 34940 19780
rect 36176 19839 36228 19848
rect 36176 19805 36185 19839
rect 36185 19805 36219 19839
rect 36219 19805 36228 19839
rect 36176 19796 36228 19805
rect 37280 19839 37332 19848
rect 37280 19805 37289 19839
rect 37289 19805 37323 19839
rect 37323 19805 37332 19839
rect 37280 19796 37332 19805
rect 39488 19796 39540 19848
rect 39304 19728 39356 19780
rect 31760 19660 31812 19712
rect 33048 19660 33100 19712
rect 34428 19660 34480 19712
rect 35716 19660 35768 19712
rect 35808 19660 35860 19712
rect 36636 19660 36688 19712
rect 36728 19660 36780 19712
rect 36912 19703 36964 19712
rect 36912 19669 36921 19703
rect 36921 19669 36955 19703
rect 36955 19669 36964 19703
rect 36912 19660 36964 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 11888 19499 11940 19508
rect 11888 19465 11897 19499
rect 11897 19465 11931 19499
rect 11931 19465 11940 19499
rect 11888 19456 11940 19465
rect 12440 19456 12492 19508
rect 12440 19320 12492 19372
rect 14464 19456 14516 19508
rect 14556 19456 14608 19508
rect 15200 19456 15252 19508
rect 16028 19456 16080 19508
rect 16120 19456 16172 19508
rect 13084 19431 13136 19440
rect 13084 19397 13093 19431
rect 13093 19397 13127 19431
rect 13127 19397 13136 19431
rect 13084 19388 13136 19397
rect 13544 19388 13596 19440
rect 15476 19388 15528 19440
rect 14096 19320 14148 19372
rect 15108 19320 15160 19372
rect 16764 19388 16816 19440
rect 17684 19456 17736 19508
rect 18696 19456 18748 19508
rect 20076 19456 20128 19508
rect 21180 19388 21232 19440
rect 23940 19456 23992 19508
rect 28724 19499 28776 19508
rect 12072 19252 12124 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 21824 19363 21876 19372
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 16028 19184 16080 19236
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 22376 19388 22428 19440
rect 23204 19388 23256 19440
rect 23388 19320 23440 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 25964 19388 26016 19440
rect 28724 19465 28733 19499
rect 28733 19465 28767 19499
rect 28767 19465 28776 19499
rect 28724 19456 28776 19465
rect 29644 19456 29696 19508
rect 29736 19456 29788 19508
rect 27160 19388 27212 19440
rect 27712 19388 27764 19440
rect 29276 19388 29328 19440
rect 31024 19456 31076 19508
rect 31392 19499 31444 19508
rect 31392 19465 31401 19499
rect 31401 19465 31435 19499
rect 31435 19465 31444 19499
rect 31392 19456 31444 19465
rect 31944 19499 31996 19508
rect 31944 19465 31953 19499
rect 31953 19465 31987 19499
rect 31987 19465 31996 19499
rect 31944 19456 31996 19465
rect 34704 19456 34756 19508
rect 34888 19499 34940 19508
rect 34888 19465 34897 19499
rect 34897 19465 34931 19499
rect 34931 19465 34940 19499
rect 34888 19456 34940 19465
rect 35532 19499 35584 19508
rect 35532 19465 35541 19499
rect 35541 19465 35575 19499
rect 35575 19465 35584 19499
rect 35532 19456 35584 19465
rect 20812 19252 20864 19304
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 15936 19116 15988 19168
rect 21456 19184 21508 19236
rect 21640 19116 21692 19168
rect 22468 19116 22520 19168
rect 26792 19320 26844 19372
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 26240 19295 26292 19304
rect 26240 19261 26249 19295
rect 26249 19261 26283 19295
rect 26283 19261 26292 19295
rect 26240 19252 26292 19261
rect 28724 19252 28776 19304
rect 29000 19320 29052 19372
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 29276 19252 29328 19304
rect 31484 19363 31536 19372
rect 31484 19329 31493 19363
rect 31493 19329 31527 19363
rect 31527 19329 31536 19363
rect 31484 19320 31536 19329
rect 33416 19320 33468 19372
rect 33876 19363 33928 19372
rect 33876 19329 33885 19363
rect 33885 19329 33919 19363
rect 33919 19329 33928 19363
rect 33876 19320 33928 19329
rect 28908 19184 28960 19236
rect 32128 19295 32180 19304
rect 32128 19261 32137 19295
rect 32137 19261 32171 19295
rect 32171 19261 32180 19295
rect 32128 19252 32180 19261
rect 33048 19252 33100 19304
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 34428 19320 34480 19329
rect 35348 19320 35400 19372
rect 35624 19320 35676 19372
rect 35900 19363 35952 19372
rect 35900 19329 35909 19363
rect 35909 19329 35943 19363
rect 35943 19329 35952 19363
rect 35900 19320 35952 19329
rect 36452 19363 36504 19372
rect 36452 19329 36461 19363
rect 36461 19329 36495 19363
rect 36495 19329 36504 19363
rect 36452 19320 36504 19329
rect 36544 19363 36596 19372
rect 36544 19329 36579 19363
rect 36579 19329 36596 19363
rect 36544 19320 36596 19329
rect 36728 19363 36780 19372
rect 36728 19329 36737 19363
rect 36737 19329 36771 19363
rect 36771 19329 36780 19363
rect 36728 19320 36780 19329
rect 36820 19363 36872 19372
rect 36820 19329 36829 19363
rect 36829 19329 36863 19363
rect 36863 19329 36872 19363
rect 36820 19320 36872 19329
rect 36912 19320 36964 19372
rect 37372 19320 37424 19372
rect 25504 19116 25556 19168
rect 36268 19184 36320 19236
rect 30748 19159 30800 19168
rect 30748 19125 30757 19159
rect 30757 19125 30791 19159
rect 30791 19125 30800 19159
rect 30748 19116 30800 19125
rect 31760 19116 31812 19168
rect 35900 19116 35952 19168
rect 37280 19116 37332 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1676 18912 1728 18964
rect 1768 18844 1820 18896
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 12440 18912 12492 18921
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 18052 18912 18104 18964
rect 17960 18844 18012 18896
rect 19156 18912 19208 18964
rect 11520 18776 11572 18828
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 15476 18776 15528 18828
rect 20812 18912 20864 18964
rect 21456 18912 21508 18964
rect 21640 18844 21692 18896
rect 21916 18887 21968 18896
rect 21916 18853 21925 18887
rect 21925 18853 21959 18887
rect 21959 18853 21968 18887
rect 21916 18844 21968 18853
rect 940 18708 992 18760
rect 15936 18751 15988 18760
rect 15936 18717 15970 18751
rect 15970 18717 15988 18751
rect 15936 18708 15988 18717
rect 18328 18708 18380 18760
rect 6920 18572 6972 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 10232 18615 10284 18624
rect 10232 18581 10241 18615
rect 10241 18581 10275 18615
rect 10275 18581 10284 18615
rect 10232 18572 10284 18581
rect 18972 18640 19024 18692
rect 15108 18572 15160 18624
rect 21088 18708 21140 18760
rect 20628 18640 20680 18692
rect 22744 18776 22796 18828
rect 22560 18640 22612 18692
rect 23020 18640 23072 18692
rect 23572 18912 23624 18964
rect 25596 18912 25648 18964
rect 23388 18776 23440 18828
rect 23664 18776 23716 18828
rect 24216 18776 24268 18828
rect 24492 18844 24544 18896
rect 26240 18844 26292 18896
rect 28816 18844 28868 18896
rect 33048 18912 33100 18964
rect 33416 18955 33468 18964
rect 33416 18921 33425 18955
rect 33425 18921 33459 18955
rect 33459 18921 33468 18955
rect 33416 18912 33468 18921
rect 25596 18708 25648 18760
rect 27712 18708 27764 18760
rect 28632 18819 28684 18828
rect 28632 18785 28641 18819
rect 28641 18785 28675 18819
rect 28675 18785 28684 18819
rect 28632 18776 28684 18785
rect 31760 18776 31812 18828
rect 30748 18708 30800 18760
rect 32220 18844 32272 18896
rect 32404 18844 32456 18896
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 31852 18640 31904 18692
rect 32036 18683 32088 18692
rect 32036 18649 32045 18683
rect 32045 18649 32079 18683
rect 32079 18649 32088 18683
rect 32036 18640 32088 18649
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 32496 18640 32548 18692
rect 34336 18751 34388 18760
rect 34336 18717 34345 18751
rect 34345 18717 34379 18751
rect 34379 18717 34388 18751
rect 34336 18708 34388 18717
rect 34612 18708 34664 18760
rect 34888 18751 34940 18760
rect 34888 18717 34897 18751
rect 34897 18717 34931 18751
rect 34931 18717 34940 18751
rect 34888 18708 34940 18717
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 22376 18572 22428 18581
rect 22468 18615 22520 18624
rect 22468 18581 22477 18615
rect 22477 18581 22511 18615
rect 22511 18581 22520 18615
rect 22468 18572 22520 18581
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 23756 18572 23808 18624
rect 25504 18572 25556 18624
rect 26148 18615 26200 18624
rect 26148 18581 26157 18615
rect 26157 18581 26191 18615
rect 26191 18581 26200 18615
rect 26148 18572 26200 18581
rect 32404 18572 32456 18624
rect 32588 18615 32640 18624
rect 32588 18581 32597 18615
rect 32597 18581 32631 18615
rect 32631 18581 32640 18615
rect 32588 18572 32640 18581
rect 33600 18572 33652 18624
rect 33692 18615 33744 18624
rect 33692 18581 33701 18615
rect 33701 18581 33735 18615
rect 33735 18581 33744 18615
rect 33692 18572 33744 18581
rect 34060 18683 34112 18692
rect 34060 18649 34069 18683
rect 34069 18649 34103 18683
rect 34103 18649 34112 18683
rect 34060 18640 34112 18649
rect 35532 18844 35584 18896
rect 35716 18955 35768 18964
rect 35716 18921 35725 18955
rect 35725 18921 35759 18955
rect 35759 18921 35768 18955
rect 35716 18912 35768 18921
rect 36176 18912 36228 18964
rect 36544 18912 36596 18964
rect 35256 18751 35308 18760
rect 35256 18717 35265 18751
rect 35265 18717 35299 18751
rect 35299 18717 35308 18751
rect 35256 18708 35308 18717
rect 37464 18776 37516 18828
rect 35624 18751 35676 18760
rect 35624 18717 35633 18751
rect 35633 18717 35667 18751
rect 35667 18717 35676 18751
rect 35624 18708 35676 18717
rect 35900 18708 35952 18760
rect 36268 18708 36320 18760
rect 37280 18640 37332 18692
rect 38568 18640 38620 18692
rect 38200 18615 38252 18624
rect 38200 18581 38209 18615
rect 38209 18581 38243 18615
rect 38243 18581 38252 18615
rect 38200 18572 38252 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9220 18368 9272 18420
rect 10232 18368 10284 18420
rect 16764 18368 16816 18420
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 18972 18368 19024 18420
rect 20628 18411 20680 18420
rect 20628 18377 20637 18411
rect 20637 18377 20671 18411
rect 20671 18377 20680 18411
rect 20628 18368 20680 18377
rect 15108 18343 15160 18352
rect 15108 18309 15117 18343
rect 15117 18309 15151 18343
rect 15151 18309 15160 18343
rect 15108 18300 15160 18309
rect 19156 18232 19208 18284
rect 11704 18207 11756 18216
rect 11704 18173 11713 18207
rect 11713 18173 11747 18207
rect 11747 18173 11756 18207
rect 11704 18164 11756 18173
rect 18328 18164 18380 18216
rect 14004 18096 14056 18148
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 11428 18028 11480 18080
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 18788 18207 18840 18216
rect 18788 18173 18797 18207
rect 18797 18173 18831 18207
rect 18831 18173 18840 18207
rect 18788 18164 18840 18173
rect 19064 18096 19116 18148
rect 21548 18368 21600 18420
rect 21732 18368 21784 18420
rect 22744 18368 22796 18420
rect 23020 18368 23072 18420
rect 23756 18411 23808 18420
rect 23756 18377 23765 18411
rect 23765 18377 23799 18411
rect 23799 18377 23808 18411
rect 23756 18368 23808 18377
rect 23940 18368 23992 18420
rect 25596 18411 25648 18420
rect 25596 18377 25605 18411
rect 25605 18377 25639 18411
rect 25639 18377 25648 18411
rect 25596 18368 25648 18377
rect 28632 18411 28684 18420
rect 28632 18377 28641 18411
rect 28641 18377 28675 18411
rect 28675 18377 28684 18411
rect 28632 18368 28684 18377
rect 32312 18368 32364 18420
rect 34336 18368 34388 18420
rect 35348 18368 35400 18420
rect 36176 18368 36228 18420
rect 38200 18368 38252 18420
rect 39304 18411 39356 18420
rect 39304 18377 39313 18411
rect 39313 18377 39347 18411
rect 39347 18377 39356 18411
rect 39304 18368 39356 18377
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 21824 18300 21876 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23388 18232 23440 18284
rect 26332 18300 26384 18352
rect 26700 18300 26752 18352
rect 26148 18275 26200 18284
rect 26148 18241 26157 18275
rect 26157 18241 26191 18275
rect 26191 18241 26200 18275
rect 26148 18232 26200 18241
rect 27712 18232 27764 18284
rect 28724 18232 28776 18284
rect 31852 18300 31904 18352
rect 32588 18300 32640 18352
rect 32036 18232 32088 18284
rect 21916 18096 21968 18148
rect 29000 18207 29052 18216
rect 29000 18173 29009 18207
rect 29009 18173 29043 18207
rect 29043 18173 29052 18207
rect 29000 18164 29052 18173
rect 30932 18164 30984 18216
rect 31484 18164 31536 18216
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 34060 18164 34112 18216
rect 36360 18164 36412 18216
rect 37464 18164 37516 18216
rect 37832 18207 37884 18216
rect 37832 18173 37841 18207
rect 37841 18173 37875 18207
rect 37875 18173 37884 18207
rect 37832 18164 37884 18173
rect 23480 18028 23532 18080
rect 26332 18071 26384 18080
rect 26332 18037 26341 18071
rect 26341 18037 26375 18071
rect 26375 18037 26384 18071
rect 26332 18028 26384 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 11704 17824 11756 17876
rect 22100 17824 22152 17876
rect 27712 17867 27764 17876
rect 27712 17833 27721 17867
rect 27721 17833 27755 17867
rect 27755 17833 27764 17867
rect 27712 17824 27764 17833
rect 30932 17867 30984 17876
rect 30932 17833 30941 17867
rect 30941 17833 30975 17867
rect 30975 17833 30984 17867
rect 30932 17824 30984 17833
rect 32220 17824 32272 17876
rect 6920 17799 6972 17808
rect 6920 17765 6929 17799
rect 6929 17765 6963 17799
rect 6963 17765 6972 17799
rect 6920 17756 6972 17765
rect 11060 17688 11112 17740
rect 11520 17688 11572 17740
rect 12348 17688 12400 17740
rect 21916 17688 21968 17740
rect 15568 17620 15620 17672
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 22744 17731 22796 17740
rect 22744 17697 22753 17731
rect 22753 17697 22787 17731
rect 22787 17697 22796 17731
rect 22744 17688 22796 17697
rect 23664 17688 23716 17740
rect 7196 17552 7248 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 10784 17552 10836 17604
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 12256 17484 12308 17536
rect 23756 17552 23808 17604
rect 15660 17484 15712 17536
rect 21824 17484 21876 17536
rect 22652 17527 22704 17536
rect 22652 17493 22661 17527
rect 22661 17493 22695 17527
rect 22695 17493 22704 17527
rect 22652 17484 22704 17493
rect 23940 17688 23992 17740
rect 26332 17688 26384 17740
rect 32404 17731 32456 17740
rect 32404 17697 32413 17731
rect 32413 17697 32447 17731
rect 32447 17697 32456 17731
rect 32404 17688 32456 17697
rect 33600 17824 33652 17876
rect 33692 17688 33744 17740
rect 34520 17731 34572 17740
rect 34520 17697 34529 17731
rect 34529 17697 34563 17731
rect 34563 17697 34572 17731
rect 34520 17688 34572 17697
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 26700 17552 26752 17604
rect 32128 17552 32180 17604
rect 32864 17552 32916 17604
rect 35808 17595 35860 17604
rect 35808 17561 35817 17595
rect 35817 17561 35851 17595
rect 35851 17561 35860 17595
rect 35808 17552 35860 17561
rect 27252 17484 27304 17536
rect 28080 17484 28132 17536
rect 37464 17484 37516 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7104 17280 7156 17332
rect 10784 17212 10836 17264
rect 11428 17212 11480 17264
rect 15660 17280 15712 17332
rect 12256 17212 12308 17264
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 15936 17212 15988 17264
rect 19248 17255 19300 17264
rect 19248 17221 19257 17255
rect 19257 17221 19291 17255
rect 19291 17221 19300 17255
rect 19248 17212 19300 17221
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 16488 17144 16540 17196
rect 19984 17323 20036 17332
rect 19984 17289 19993 17323
rect 19993 17289 20027 17323
rect 20027 17289 20036 17323
rect 19984 17280 20036 17289
rect 20352 17280 20404 17332
rect 23204 17212 23256 17264
rect 26700 17212 26752 17264
rect 27528 17212 27580 17264
rect 28908 17280 28960 17332
rect 37832 17280 37884 17332
rect 39120 17280 39172 17332
rect 40592 17280 40644 17332
rect 30932 17212 30984 17264
rect 32128 17212 32180 17264
rect 16856 17119 16908 17128
rect 16856 17085 16865 17119
rect 16865 17085 16899 17119
rect 16899 17085 16908 17119
rect 16856 17076 16908 17085
rect 17592 17076 17644 17128
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 17868 17119 17920 17128
rect 17868 17085 17902 17119
rect 17902 17085 17920 17119
rect 17868 17076 17920 17085
rect 16396 17008 16448 17060
rect 17500 17051 17552 17060
rect 17500 17017 17509 17051
rect 17509 17017 17543 17051
rect 17543 17017 17552 17051
rect 17500 17008 17552 17017
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 14280 16940 14332 16992
rect 16120 16940 16172 16992
rect 18696 17076 18748 17128
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 18972 17008 19024 17060
rect 22376 17144 22428 17196
rect 38016 17187 38068 17196
rect 38016 17153 38025 17187
rect 38025 17153 38059 17187
rect 38059 17153 38068 17187
rect 38016 17144 38068 17153
rect 21824 17119 21876 17128
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 22928 17008 22980 17060
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 20260 16983 20312 16992
rect 20260 16949 20269 16983
rect 20269 16949 20303 16983
rect 20303 16949 20312 16983
rect 20260 16940 20312 16949
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 28908 17076 28960 17128
rect 35440 17076 35492 17128
rect 44640 17008 44692 17060
rect 27620 16940 27672 16992
rect 31116 16983 31168 16992
rect 31116 16949 31125 16983
rect 31125 16949 31159 16983
rect 31159 16949 31168 16983
rect 31116 16940 31168 16949
rect 35900 16940 35952 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 14464 16600 14516 16652
rect 16856 16736 16908 16788
rect 17592 16736 17644 16788
rect 18788 16779 18840 16788
rect 18788 16745 18797 16779
rect 18797 16745 18831 16779
rect 18831 16745 18840 16779
rect 18788 16736 18840 16745
rect 20260 16736 20312 16788
rect 27528 16736 27580 16788
rect 28080 16736 28132 16788
rect 35992 16736 36044 16788
rect 37280 16736 37332 16788
rect 14832 16600 14884 16652
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 15108 16575 15160 16584
rect 15108 16541 15142 16575
rect 15142 16541 15160 16575
rect 15936 16600 15988 16652
rect 16120 16600 16172 16652
rect 16396 16600 16448 16652
rect 15108 16532 15160 16541
rect 9680 16464 9732 16516
rect 10784 16464 10836 16516
rect 15844 16464 15896 16516
rect 17500 16643 17552 16652
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 18420 16600 18472 16652
rect 23388 16600 23440 16652
rect 9496 16396 9548 16448
rect 15568 16396 15620 16448
rect 17132 16396 17184 16448
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 18972 16532 19024 16584
rect 23112 16532 23164 16584
rect 23480 16532 23532 16584
rect 23572 16532 23624 16584
rect 24492 16532 24544 16584
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 24952 16532 25004 16541
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 25412 16600 25464 16652
rect 25320 16532 25372 16584
rect 31944 16668 31996 16720
rect 27620 16643 27672 16652
rect 27620 16609 27629 16643
rect 27629 16609 27663 16643
rect 27663 16609 27672 16643
rect 27620 16600 27672 16609
rect 28908 16532 28960 16584
rect 29184 16532 29236 16584
rect 33048 16532 33100 16584
rect 34520 16600 34572 16652
rect 37464 16600 37516 16652
rect 38200 16532 38252 16584
rect 44548 16575 44600 16584
rect 44548 16541 44557 16575
rect 44557 16541 44591 16575
rect 44591 16541 44600 16575
rect 44548 16532 44600 16541
rect 28172 16464 28224 16516
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 18696 16396 18748 16448
rect 23664 16396 23716 16448
rect 36820 16464 36872 16516
rect 29368 16439 29420 16448
rect 29368 16405 29377 16439
rect 29377 16405 29411 16439
rect 29411 16405 29420 16439
rect 29368 16396 29420 16405
rect 32956 16439 33008 16448
rect 32956 16405 32965 16439
rect 32965 16405 32999 16439
rect 32999 16405 33008 16439
rect 32956 16396 33008 16405
rect 35440 16396 35492 16448
rect 36728 16439 36780 16448
rect 36728 16405 36737 16439
rect 36737 16405 36771 16439
rect 36771 16405 36780 16439
rect 36728 16396 36780 16405
rect 38384 16396 38436 16448
rect 44732 16439 44784 16448
rect 44732 16405 44741 16439
rect 44741 16405 44775 16439
rect 44775 16405 44784 16439
rect 44732 16396 44784 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 9680 16192 9732 16244
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 14096 16192 14148 16244
rect 15292 16192 15344 16244
rect 9496 16167 9548 16176
rect 9496 16133 9505 16167
rect 9505 16133 9539 16167
rect 9539 16133 9548 16167
rect 9496 16124 9548 16133
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 14924 16124 14976 16176
rect 17040 16192 17092 16244
rect 19432 16192 19484 16244
rect 7104 15988 7156 16040
rect 13912 16056 13964 16108
rect 14832 16056 14884 16108
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 8944 15988 8996 16040
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 1584 15920 1636 15972
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 13544 15852 13596 15904
rect 15568 16056 15620 16108
rect 15752 15852 15804 15904
rect 16120 15988 16172 16040
rect 16856 15988 16908 16040
rect 16028 15920 16080 15972
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 22284 16192 22336 16244
rect 22376 16192 22428 16244
rect 22928 16235 22980 16244
rect 22928 16201 22937 16235
rect 22937 16201 22971 16235
rect 22971 16201 22980 16235
rect 22928 16192 22980 16201
rect 23204 16192 23256 16244
rect 25136 16235 25188 16244
rect 25136 16201 25145 16235
rect 25145 16201 25179 16235
rect 25179 16201 25188 16235
rect 25136 16192 25188 16201
rect 28172 16192 28224 16244
rect 17408 16056 17460 16108
rect 18696 16056 18748 16108
rect 21088 16056 21140 16108
rect 23020 16124 23072 16176
rect 23572 16124 23624 16176
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 17868 15988 17920 16040
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 23388 16099 23440 16108
rect 23388 16065 23397 16099
rect 23397 16065 23431 16099
rect 23431 16065 23440 16099
rect 23388 16056 23440 16065
rect 23572 15988 23624 16040
rect 21824 15920 21876 15972
rect 22928 15920 22980 15972
rect 23020 15920 23072 15972
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 24492 15988 24544 16040
rect 23756 15920 23808 15972
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 27896 16167 27948 16176
rect 27896 16133 27905 16167
rect 27905 16133 27939 16167
rect 27939 16133 27948 16167
rect 27896 16124 27948 16133
rect 29184 16124 29236 16176
rect 30932 16124 30984 16176
rect 32956 16192 33008 16244
rect 35900 16192 35952 16244
rect 35992 16235 36044 16244
rect 35992 16201 36001 16235
rect 36001 16201 36035 16235
rect 36035 16201 36044 16235
rect 35992 16192 36044 16201
rect 36728 16192 36780 16244
rect 38016 16235 38068 16244
rect 38016 16201 38025 16235
rect 38025 16201 38059 16235
rect 38059 16201 38068 16235
rect 38016 16192 38068 16201
rect 32864 16124 32916 16176
rect 34152 16167 34204 16176
rect 34152 16133 34161 16167
rect 34161 16133 34195 16167
rect 34195 16133 34204 16167
rect 34152 16124 34204 16133
rect 25320 16099 25372 16108
rect 25320 16065 25329 16099
rect 25329 16065 25363 16099
rect 25363 16065 25372 16099
rect 25320 16056 25372 16065
rect 27620 16099 27672 16108
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 29368 16056 29420 16108
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 25412 16031 25464 16040
rect 25412 15997 25421 16031
rect 25421 15997 25455 16031
rect 25455 15997 25464 16031
rect 25412 15988 25464 15997
rect 25596 16031 25648 16040
rect 25596 15997 25605 16031
rect 25605 15997 25639 16031
rect 25639 15997 25648 16031
rect 25596 15988 25648 15997
rect 26056 15988 26108 16040
rect 31116 16056 31168 16108
rect 31208 16056 31260 16108
rect 31668 16099 31720 16108
rect 31668 16065 31670 16099
rect 31670 16065 31704 16099
rect 31704 16065 31720 16099
rect 31668 16056 31720 16065
rect 32220 16056 32272 16108
rect 37464 16124 37516 16176
rect 41880 16124 41932 16176
rect 37832 16056 37884 16108
rect 31484 16031 31536 16040
rect 31484 15997 31493 16031
rect 31493 15997 31527 16031
rect 31527 15997 31536 16031
rect 31484 15988 31536 15997
rect 33048 15988 33100 16040
rect 16764 15852 16816 15904
rect 17776 15852 17828 15904
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 20168 15852 20220 15904
rect 21732 15852 21784 15904
rect 23664 15852 23716 15904
rect 24492 15852 24544 15904
rect 29000 15852 29052 15904
rect 29368 15895 29420 15904
rect 29368 15861 29377 15895
rect 29377 15861 29411 15895
rect 29411 15861 29420 15895
rect 29368 15852 29420 15861
rect 30748 15895 30800 15904
rect 30748 15861 30757 15895
rect 30757 15861 30791 15895
rect 30791 15861 30800 15895
rect 30748 15852 30800 15861
rect 31760 15852 31812 15904
rect 31852 15895 31904 15904
rect 31852 15861 31861 15895
rect 31861 15861 31895 15895
rect 31895 15861 31904 15895
rect 31852 15852 31904 15861
rect 34060 15895 34112 15904
rect 34060 15861 34069 15895
rect 34069 15861 34103 15895
rect 34103 15861 34112 15895
rect 34060 15852 34112 15861
rect 41604 15988 41656 16040
rect 44364 15988 44416 16040
rect 43812 15963 43864 15972
rect 43812 15929 43821 15963
rect 43821 15929 43855 15963
rect 43855 15929 43864 15963
rect 43812 15920 43864 15929
rect 35808 15852 35860 15904
rect 37188 15852 37240 15904
rect 37924 15895 37976 15904
rect 37924 15861 37933 15895
rect 37933 15861 37967 15895
rect 37967 15861 37976 15895
rect 37924 15852 37976 15861
rect 38384 15895 38436 15904
rect 38384 15861 38393 15895
rect 38393 15861 38427 15895
rect 38427 15861 38436 15895
rect 38384 15852 38436 15861
rect 38568 15852 38620 15904
rect 39764 15852 39816 15904
rect 42248 15852 42300 15904
rect 43996 15895 44048 15904
rect 43996 15861 44005 15895
rect 44005 15861 44039 15895
rect 44039 15861 44048 15895
rect 43996 15852 44048 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8300 15648 8352 15700
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 14280 15648 14332 15700
rect 15108 15648 15160 15700
rect 13544 15580 13596 15632
rect 13176 15512 13228 15564
rect 17868 15648 17920 15700
rect 18052 15648 18104 15700
rect 20536 15691 20588 15700
rect 20536 15657 20545 15691
rect 20545 15657 20579 15691
rect 20579 15657 20588 15691
rect 20536 15648 20588 15657
rect 21088 15648 21140 15700
rect 21180 15648 21232 15700
rect 22468 15648 22520 15700
rect 14924 15512 14976 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 8392 15444 8444 15496
rect 8944 15487 8996 15496
rect 8944 15453 8953 15487
rect 8953 15453 8987 15487
rect 8987 15453 8996 15487
rect 8944 15444 8996 15453
rect 12164 15444 12216 15496
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 9680 15376 9732 15428
rect 11428 15419 11480 15428
rect 11428 15385 11437 15419
rect 11437 15385 11471 15419
rect 11471 15385 11480 15419
rect 11428 15376 11480 15385
rect 13636 15376 13688 15428
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 14004 15376 14056 15428
rect 15200 15487 15252 15496
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 15660 15580 15712 15632
rect 20628 15580 20680 15632
rect 15752 15512 15804 15564
rect 15292 15376 15344 15428
rect 15844 15444 15896 15496
rect 16028 15444 16080 15496
rect 16764 15444 16816 15496
rect 17408 15444 17460 15496
rect 17592 15512 17644 15564
rect 16672 15376 16724 15428
rect 14648 15308 14700 15360
rect 17408 15308 17460 15360
rect 18144 15376 18196 15428
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 21824 15580 21876 15632
rect 22744 15580 22796 15632
rect 21640 15555 21692 15564
rect 21640 15521 21649 15555
rect 21649 15521 21683 15555
rect 21683 15521 21692 15555
rect 21640 15512 21692 15521
rect 21732 15555 21784 15564
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 22376 15512 22428 15564
rect 23020 15648 23072 15700
rect 23112 15648 23164 15700
rect 24032 15648 24084 15700
rect 24308 15648 24360 15700
rect 24676 15648 24728 15700
rect 25044 15648 25096 15700
rect 26516 15648 26568 15700
rect 29000 15648 29052 15700
rect 30012 15648 30064 15700
rect 30564 15648 30616 15700
rect 34060 15648 34112 15700
rect 18328 15308 18380 15360
rect 19340 15308 19392 15360
rect 19708 15308 19760 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 20076 15308 20128 15360
rect 20812 15376 20864 15428
rect 21916 15487 21968 15496
rect 21916 15453 21925 15487
rect 21925 15453 21959 15487
rect 21959 15453 21968 15487
rect 21916 15444 21968 15453
rect 22100 15444 22152 15496
rect 21824 15376 21876 15428
rect 22468 15444 22520 15496
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 22652 15444 22704 15496
rect 23020 15444 23072 15496
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23388 15419 23440 15428
rect 23388 15385 23397 15419
rect 23397 15385 23431 15419
rect 23431 15385 23440 15419
rect 23388 15376 23440 15385
rect 24124 15512 24176 15564
rect 23756 15487 23808 15496
rect 23756 15453 23765 15487
rect 23765 15453 23799 15487
rect 23799 15453 23808 15487
rect 23756 15444 23808 15453
rect 25872 15512 25924 15564
rect 26792 15512 26844 15564
rect 29644 15512 29696 15564
rect 31668 15580 31720 15632
rect 24492 15376 24544 15428
rect 22744 15308 22796 15360
rect 22928 15308 22980 15360
rect 23848 15308 23900 15360
rect 24124 15308 24176 15360
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 29368 15444 29420 15496
rect 30288 15444 30340 15496
rect 30472 15444 30524 15496
rect 31208 15444 31260 15496
rect 31484 15487 31536 15496
rect 31484 15453 31493 15487
rect 31493 15453 31527 15487
rect 31527 15453 31536 15487
rect 31484 15444 31536 15453
rect 31760 15487 31812 15496
rect 31760 15453 31769 15487
rect 31769 15453 31803 15487
rect 31803 15453 31812 15487
rect 31760 15444 31812 15453
rect 37464 15648 37516 15700
rect 37924 15648 37976 15700
rect 41604 15691 41656 15700
rect 41604 15657 41613 15691
rect 41613 15657 41647 15691
rect 41647 15657 41656 15691
rect 41604 15648 41656 15657
rect 43812 15648 43864 15700
rect 39120 15555 39172 15564
rect 39120 15521 39129 15555
rect 39129 15521 39163 15555
rect 39163 15521 39172 15555
rect 39120 15512 39172 15521
rect 40684 15512 40736 15564
rect 42248 15512 42300 15564
rect 24676 15376 24728 15428
rect 24952 15376 25004 15428
rect 25136 15308 25188 15360
rect 26332 15351 26384 15360
rect 26332 15317 26341 15351
rect 26341 15317 26375 15351
rect 26375 15317 26384 15351
rect 26332 15308 26384 15317
rect 26884 15308 26936 15360
rect 31576 15376 31628 15428
rect 30564 15308 30616 15360
rect 32312 15376 32364 15428
rect 37740 15487 37792 15496
rect 37740 15453 37749 15487
rect 37749 15453 37783 15487
rect 37783 15453 37792 15487
rect 37740 15444 37792 15453
rect 35440 15419 35492 15428
rect 35440 15385 35449 15419
rect 35449 15385 35483 15419
rect 35483 15385 35492 15419
rect 35440 15376 35492 15385
rect 36820 15376 36872 15428
rect 35348 15351 35400 15360
rect 35348 15317 35357 15351
rect 35357 15317 35391 15351
rect 35391 15317 35400 15351
rect 35348 15308 35400 15317
rect 35900 15351 35952 15360
rect 35900 15317 35909 15351
rect 35909 15317 35943 15351
rect 35943 15317 35952 15351
rect 35900 15308 35952 15317
rect 38660 15419 38712 15428
rect 38660 15385 38678 15419
rect 38678 15385 38712 15419
rect 38660 15376 38712 15385
rect 38752 15351 38804 15360
rect 38752 15317 38761 15351
rect 38761 15317 38795 15351
rect 38795 15317 38804 15351
rect 38752 15308 38804 15317
rect 39028 15308 39080 15360
rect 39764 15308 39816 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 13084 15104 13136 15156
rect 13176 15104 13228 15156
rect 13452 15036 13504 15088
rect 13820 15036 13872 15088
rect 7012 14968 7064 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 8760 14900 8812 14952
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 12164 14968 12216 15020
rect 12256 14968 12308 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 13176 15011 13228 15020
rect 13176 14977 13179 15011
rect 13179 14977 13213 15011
rect 13213 14977 13228 15011
rect 13176 14968 13228 14977
rect 14464 15104 14516 15156
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 15200 15104 15252 15156
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 17040 15104 17092 15156
rect 17316 15104 17368 15156
rect 18512 15104 18564 15156
rect 18604 15104 18656 15156
rect 16304 15036 16356 15088
rect 17500 15036 17552 15088
rect 18052 15036 18104 15088
rect 20812 15104 20864 15156
rect 22560 15104 22612 15156
rect 22744 15104 22796 15156
rect 23664 15104 23716 15156
rect 15752 14968 15804 15020
rect 16672 14968 16724 15020
rect 18512 14968 18564 15020
rect 18604 14968 18656 15020
rect 16948 14900 17000 14952
rect 12900 14764 12952 14816
rect 13820 14832 13872 14884
rect 14280 14875 14332 14884
rect 14280 14841 14289 14875
rect 14289 14841 14323 14875
rect 14323 14841 14332 14875
rect 14280 14832 14332 14841
rect 14372 14764 14424 14816
rect 15568 14764 15620 14816
rect 16764 14764 16816 14816
rect 17040 14764 17092 14816
rect 17684 14943 17736 14952
rect 17684 14909 17693 14943
rect 17693 14909 17727 14943
rect 17727 14909 17736 14943
rect 17684 14900 17736 14909
rect 17776 14943 17828 14952
rect 17776 14909 17785 14943
rect 17785 14909 17819 14943
rect 17819 14909 17828 14943
rect 17776 14900 17828 14909
rect 19984 14968 20036 15020
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 20536 14968 20588 15020
rect 20628 14968 20680 15020
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21916 15036 21968 15088
rect 19156 14832 19208 14884
rect 17592 14764 17644 14816
rect 20076 14900 20128 14952
rect 22468 14968 22520 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23480 15036 23532 15088
rect 30748 15104 30800 15156
rect 34520 15104 34572 15156
rect 35900 15104 35952 15156
rect 37280 15147 37332 15156
rect 37280 15113 37289 15147
rect 37289 15113 37323 15147
rect 37323 15113 37332 15147
rect 37280 15104 37332 15113
rect 43996 15104 44048 15156
rect 44548 15104 44600 15156
rect 25596 14968 25648 15020
rect 25964 15011 26016 15020
rect 25964 14977 25973 15011
rect 25973 14977 26007 15011
rect 26007 14977 26016 15011
rect 25964 14968 26016 14977
rect 20720 14875 20772 14884
rect 20720 14841 20729 14875
rect 20729 14841 20763 14875
rect 20763 14841 20772 14875
rect 20720 14832 20772 14841
rect 26884 14968 26936 15020
rect 29000 14968 29052 15020
rect 25872 14900 25924 14952
rect 26332 14900 26384 14952
rect 27068 14900 27120 14952
rect 29644 15011 29696 15020
rect 29644 14977 29653 15011
rect 29653 14977 29687 15011
rect 29687 14977 29696 15011
rect 29644 14968 29696 14977
rect 30012 14968 30064 15020
rect 30288 14968 30340 15020
rect 30472 15011 30524 15020
rect 30472 14977 30481 15011
rect 30481 14977 30515 15011
rect 30515 14977 30524 15011
rect 30472 14968 30524 14977
rect 30564 14968 30616 15020
rect 34428 15036 34480 15088
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 31484 14968 31536 15020
rect 35348 15036 35400 15088
rect 31208 14900 31260 14952
rect 35716 14943 35768 14952
rect 35716 14909 35725 14943
rect 35725 14909 35759 14943
rect 35759 14909 35768 14943
rect 35716 14900 35768 14909
rect 37832 14943 37884 14952
rect 37832 14909 37841 14943
rect 37841 14909 37875 14943
rect 37875 14909 37884 14943
rect 37832 14900 37884 14909
rect 19616 14764 19668 14816
rect 20352 14764 20404 14816
rect 20444 14764 20496 14816
rect 20812 14764 20864 14816
rect 22560 14807 22612 14816
rect 22560 14773 22569 14807
rect 22569 14773 22603 14807
rect 22603 14773 22612 14807
rect 22560 14764 22612 14773
rect 23756 14764 23808 14816
rect 26148 14764 26200 14816
rect 29460 14764 29512 14816
rect 30288 14807 30340 14816
rect 30288 14773 30297 14807
rect 30297 14773 30331 14807
rect 30331 14773 30340 14807
rect 30288 14764 30340 14773
rect 31484 14764 31536 14816
rect 35348 14764 35400 14816
rect 36360 14764 36412 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7012 14560 7064 14612
rect 8760 14603 8812 14612
rect 8760 14569 8769 14603
rect 8769 14569 8803 14603
rect 8803 14569 8812 14603
rect 8760 14560 8812 14569
rect 10232 14560 10284 14612
rect 11980 14603 12032 14612
rect 11980 14569 11989 14603
rect 11989 14569 12023 14603
rect 12023 14569 12032 14603
rect 11980 14560 12032 14569
rect 12164 14603 12216 14612
rect 12164 14569 12173 14603
rect 12173 14569 12207 14603
rect 12207 14569 12216 14603
rect 12164 14560 12216 14569
rect 12532 14560 12584 14612
rect 13820 14560 13872 14612
rect 14096 14560 14148 14612
rect 15292 14560 15344 14612
rect 15844 14603 15896 14612
rect 15844 14569 15853 14603
rect 15853 14569 15887 14603
rect 15887 14569 15896 14603
rect 15844 14560 15896 14569
rect 8944 14467 8996 14476
rect 8944 14433 8953 14467
rect 8953 14433 8987 14467
rect 8987 14433 8996 14467
rect 8944 14424 8996 14433
rect 11796 14492 11848 14544
rect 13636 14492 13688 14544
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 16764 14492 16816 14544
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 18144 14560 18196 14612
rect 20444 14560 20496 14612
rect 20812 14560 20864 14612
rect 22560 14560 22612 14612
rect 23204 14560 23256 14612
rect 23388 14560 23440 14612
rect 25136 14603 25188 14612
rect 25136 14569 25145 14603
rect 25145 14569 25179 14603
rect 25179 14569 25188 14603
rect 25136 14560 25188 14569
rect 26148 14603 26200 14612
rect 26148 14569 26157 14603
rect 26157 14569 26191 14603
rect 26191 14569 26200 14603
rect 26148 14560 26200 14569
rect 26976 14560 27028 14612
rect 29368 14560 29420 14612
rect 30288 14560 30340 14612
rect 31576 14560 31628 14612
rect 35716 14560 35768 14612
rect 7288 14331 7340 14340
rect 7288 14297 7297 14331
rect 7297 14297 7331 14331
rect 7331 14297 7340 14331
rect 7288 14288 7340 14297
rect 9680 14288 9732 14340
rect 15108 14399 15160 14408
rect 15108 14365 15117 14399
rect 15117 14365 15151 14399
rect 15151 14365 15160 14399
rect 15108 14356 15160 14365
rect 15568 14424 15620 14476
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 16672 14467 16724 14476
rect 16672 14433 16681 14467
rect 16681 14433 16715 14467
rect 16715 14433 16724 14467
rect 16672 14424 16724 14433
rect 16948 14424 17000 14476
rect 17960 14467 18012 14476
rect 17960 14433 17969 14467
rect 17969 14433 18003 14467
rect 18003 14433 18012 14467
rect 17960 14424 18012 14433
rect 18144 14424 18196 14476
rect 19248 14492 19300 14544
rect 19616 14492 19668 14544
rect 10692 14263 10744 14272
rect 10692 14229 10701 14263
rect 10701 14229 10735 14263
rect 10735 14229 10744 14263
rect 10692 14220 10744 14229
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 11888 14220 11940 14272
rect 13176 14220 13228 14272
rect 13360 14220 13412 14272
rect 14556 14220 14608 14272
rect 15108 14220 15160 14272
rect 15752 14288 15804 14340
rect 16028 14356 16080 14408
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17500 14356 17552 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 15384 14220 15436 14272
rect 15936 14220 15988 14272
rect 16396 14220 16448 14272
rect 17960 14288 18012 14340
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 19156 14356 19208 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 20536 14288 20588 14340
rect 18972 14220 19024 14272
rect 19432 14220 19484 14272
rect 20260 14220 20312 14272
rect 21824 14424 21876 14476
rect 25872 14424 25924 14476
rect 26792 14424 26844 14476
rect 21732 14288 21784 14340
rect 25596 14263 25648 14272
rect 25596 14229 25605 14263
rect 25605 14229 25639 14263
rect 25639 14229 25648 14263
rect 25596 14220 25648 14229
rect 26516 14263 26568 14272
rect 26516 14229 26525 14263
rect 26525 14229 26559 14263
rect 26559 14229 26568 14263
rect 26516 14220 26568 14229
rect 30012 14424 30064 14476
rect 31760 14424 31812 14476
rect 30380 14356 30432 14408
rect 31852 14288 31904 14340
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32128 14356 32180 14365
rect 34520 14424 34572 14476
rect 35348 14424 35400 14476
rect 35992 14356 36044 14408
rect 36820 14356 36872 14408
rect 38660 14356 38712 14408
rect 33140 14288 33192 14340
rect 26700 14220 26752 14272
rect 27068 14220 27120 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 7288 14016 7340 14068
rect 11520 14016 11572 14068
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 11980 13880 12032 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 14096 14016 14148 14068
rect 14280 14016 14332 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 15292 14016 15344 14068
rect 13360 13948 13412 14000
rect 13820 13948 13872 14000
rect 17776 14016 17828 14068
rect 20444 14016 20496 14068
rect 24308 14059 24360 14068
rect 24308 14025 24317 14059
rect 24317 14025 24351 14059
rect 24351 14025 24360 14059
rect 24308 14016 24360 14025
rect 24860 14016 24912 14068
rect 25044 14059 25096 14068
rect 25044 14025 25053 14059
rect 25053 14025 25087 14059
rect 25087 14025 25096 14059
rect 25044 14016 25096 14025
rect 26148 14016 26200 14068
rect 26608 14016 26660 14068
rect 26700 14016 26752 14068
rect 27252 14016 27304 14068
rect 28908 14016 28960 14068
rect 13084 13880 13136 13932
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 13820 13812 13872 13864
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 14188 13812 14240 13864
rect 15200 13812 15252 13864
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 15752 13880 15804 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16396 13880 16448 13932
rect 18512 13948 18564 14000
rect 18788 13948 18840 14000
rect 20076 13948 20128 14000
rect 20720 13880 20772 13932
rect 16580 13812 16632 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 17500 13812 17552 13864
rect 19156 13812 19208 13864
rect 11244 13676 11296 13728
rect 11336 13676 11388 13728
rect 14004 13676 14056 13728
rect 14740 13676 14792 13728
rect 16304 13676 16356 13728
rect 17040 13676 17092 13728
rect 17224 13676 17276 13728
rect 17592 13676 17644 13728
rect 18972 13676 19024 13728
rect 24124 13744 24176 13796
rect 24676 13880 24728 13932
rect 25596 13880 25648 13932
rect 30840 13948 30892 14000
rect 31392 13948 31444 14000
rect 32128 14016 32180 14068
rect 37280 14016 37332 14068
rect 31024 13880 31076 13932
rect 24584 13812 24636 13864
rect 24952 13744 25004 13796
rect 26792 13744 26844 13796
rect 29092 13855 29144 13864
rect 29092 13821 29101 13855
rect 29101 13821 29135 13855
rect 29135 13821 29144 13855
rect 29092 13812 29144 13821
rect 31944 13880 31996 13932
rect 33140 13991 33192 14000
rect 33140 13957 33149 13991
rect 33149 13957 33183 13991
rect 33183 13957 33192 13991
rect 33140 13948 33192 13957
rect 35992 13948 36044 14000
rect 36360 13948 36412 14000
rect 36820 13948 36872 14000
rect 34428 13880 34480 13932
rect 37740 13880 37792 13932
rect 35992 13812 36044 13864
rect 30932 13676 30984 13728
rect 31116 13676 31168 13728
rect 34612 13719 34664 13728
rect 34612 13685 34621 13719
rect 34621 13685 34655 13719
rect 34655 13685 34664 13719
rect 34612 13676 34664 13685
rect 39580 13719 39632 13728
rect 39580 13685 39589 13719
rect 39589 13685 39623 13719
rect 39623 13685 39632 13719
rect 39580 13676 39632 13685
rect 40684 13744 40736 13796
rect 41236 13744 41288 13796
rect 43628 13744 43680 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7196 13472 7248 13524
rect 6920 13447 6972 13456
rect 6920 13413 6929 13447
rect 6929 13413 6963 13447
rect 6963 13413 6972 13447
rect 6920 13404 6972 13413
rect 7012 13336 7064 13388
rect 11336 13472 11388 13524
rect 12348 13472 12400 13524
rect 12532 13472 12584 13524
rect 14004 13472 14056 13524
rect 24952 13472 25004 13524
rect 26608 13515 26660 13524
rect 26608 13481 26617 13515
rect 26617 13481 26651 13515
rect 26651 13481 26660 13515
rect 26608 13472 26660 13481
rect 26792 13472 26844 13524
rect 34152 13472 34204 13524
rect 37832 13472 37884 13524
rect 16672 13404 16724 13456
rect 22284 13404 22336 13456
rect 24124 13447 24176 13456
rect 24124 13413 24133 13447
rect 24133 13413 24167 13447
rect 24167 13413 24176 13447
rect 24124 13404 24176 13413
rect 25596 13404 25648 13456
rect 26056 13447 26108 13456
rect 26056 13413 26065 13447
rect 26065 13413 26099 13447
rect 26099 13413 26108 13447
rect 26056 13404 26108 13413
rect 8944 13379 8996 13388
rect 8944 13345 8953 13379
rect 8953 13345 8987 13379
rect 8987 13345 8996 13379
rect 8944 13336 8996 13345
rect 11796 13336 11848 13388
rect 14740 13336 14792 13388
rect 15108 13336 15160 13388
rect 19340 13336 19392 13388
rect 21916 13379 21968 13388
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 23020 13336 23072 13388
rect 24860 13336 24912 13388
rect 9220 13243 9272 13252
rect 9220 13209 9229 13243
rect 9229 13209 9263 13243
rect 9263 13209 9272 13243
rect 9220 13200 9272 13209
rect 9956 13200 10008 13252
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12900 13200 12952 13252
rect 11336 13132 11388 13184
rect 11428 13132 11480 13184
rect 12624 13132 12676 13184
rect 13084 13268 13136 13320
rect 13636 13268 13688 13320
rect 15476 13268 15528 13320
rect 16580 13268 16632 13320
rect 13728 13200 13780 13252
rect 16672 13200 16724 13252
rect 17960 13268 18012 13320
rect 19156 13268 19208 13320
rect 20812 13268 20864 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 22376 13311 22428 13320
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 24400 13268 24452 13320
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 27252 13447 27304 13456
rect 27252 13413 27261 13447
rect 27261 13413 27295 13447
rect 27295 13413 27304 13447
rect 27252 13404 27304 13413
rect 31024 13404 31076 13456
rect 31208 13404 31260 13456
rect 31576 13447 31628 13456
rect 31576 13413 31585 13447
rect 31585 13413 31619 13447
rect 31619 13413 31628 13447
rect 31576 13404 31628 13413
rect 31852 13404 31904 13456
rect 27712 13379 27764 13388
rect 27712 13345 27721 13379
rect 27721 13345 27755 13379
rect 27755 13345 27764 13379
rect 27712 13336 27764 13345
rect 18236 13200 18288 13252
rect 20260 13200 20312 13252
rect 22192 13200 22244 13252
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 15936 13132 15988 13184
rect 16764 13132 16816 13184
rect 19340 13132 19392 13184
rect 20628 13132 20680 13184
rect 25780 13200 25832 13252
rect 26608 13268 26660 13320
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 26976 13268 27028 13320
rect 29276 13311 29328 13320
rect 29276 13277 29285 13311
rect 29285 13277 29319 13311
rect 29319 13277 29328 13311
rect 29276 13268 29328 13277
rect 30932 13268 30984 13320
rect 31668 13268 31720 13320
rect 31760 13311 31812 13320
rect 31760 13277 31769 13311
rect 31769 13277 31803 13311
rect 31803 13277 31812 13311
rect 31760 13268 31812 13277
rect 32128 13268 32180 13320
rect 38752 13336 38804 13388
rect 39580 13336 39632 13388
rect 32680 13268 32732 13320
rect 34152 13268 34204 13320
rect 34612 13268 34664 13320
rect 35624 13311 35676 13320
rect 35624 13277 35633 13311
rect 35633 13277 35667 13311
rect 35667 13277 35676 13311
rect 35624 13268 35676 13277
rect 36084 13268 36136 13320
rect 26240 13132 26292 13184
rect 26516 13132 26568 13184
rect 27620 13175 27672 13184
rect 27620 13141 27629 13175
rect 27629 13141 27663 13175
rect 27663 13141 27672 13175
rect 27620 13132 27672 13141
rect 28448 13175 28500 13184
rect 28448 13141 28457 13175
rect 28457 13141 28491 13175
rect 28491 13141 28500 13175
rect 28448 13132 28500 13141
rect 28908 13175 28960 13184
rect 28908 13141 28917 13175
rect 28917 13141 28951 13175
rect 28951 13141 28960 13175
rect 28908 13132 28960 13141
rect 29000 13132 29052 13184
rect 29920 13132 29972 13184
rect 31944 13243 31996 13252
rect 31944 13209 31953 13243
rect 31953 13209 31987 13243
rect 31987 13209 31996 13243
rect 31944 13200 31996 13209
rect 36728 13311 36780 13320
rect 36728 13277 36737 13311
rect 36737 13277 36771 13311
rect 36771 13277 36780 13311
rect 36728 13268 36780 13277
rect 37096 13268 37148 13320
rect 37464 13311 37516 13320
rect 37464 13277 37473 13311
rect 37473 13277 37507 13311
rect 37507 13277 37516 13311
rect 37464 13268 37516 13277
rect 37924 13268 37976 13320
rect 39028 13268 39080 13320
rect 41236 13336 41288 13388
rect 41328 13268 41380 13320
rect 34704 13132 34756 13184
rect 34888 13175 34940 13184
rect 34888 13141 34897 13175
rect 34897 13141 34931 13175
rect 34931 13141 34940 13175
rect 34888 13132 34940 13141
rect 35440 13132 35492 13184
rect 40500 13175 40552 13184
rect 40500 13141 40509 13175
rect 40509 13141 40543 13175
rect 40543 13141 40552 13175
rect 40500 13132 40552 13141
rect 43812 13243 43864 13252
rect 43812 13209 43821 13243
rect 43821 13209 43855 13243
rect 43855 13209 43864 13243
rect 43812 13200 43864 13209
rect 44364 13132 44416 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9220 12928 9272 12980
rect 11612 12928 11664 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 7012 12860 7064 12912
rect 12072 12860 12124 12912
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 11612 12792 11664 12844
rect 11980 12792 12032 12844
rect 13084 12928 13136 12980
rect 13360 12928 13412 12980
rect 14832 12928 14884 12980
rect 12348 12792 12400 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 1584 12656 1636 12708
rect 12992 12656 13044 12708
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 15844 12928 15896 12980
rect 16488 12928 16540 12980
rect 16672 12928 16724 12980
rect 14556 12724 14608 12776
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 15476 12724 15528 12776
rect 15660 12724 15712 12776
rect 16764 12860 16816 12912
rect 9956 12588 10008 12640
rect 11612 12588 11664 12640
rect 12440 12588 12492 12640
rect 12532 12588 12584 12640
rect 13728 12588 13780 12640
rect 14832 12588 14884 12640
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 18788 12928 18840 12980
rect 19432 12928 19484 12980
rect 20168 12928 20220 12980
rect 21916 12928 21968 12980
rect 22100 12928 22152 12980
rect 23204 12971 23256 12980
rect 23204 12937 23213 12971
rect 23213 12937 23247 12971
rect 23247 12937 23256 12971
rect 23204 12928 23256 12937
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 26240 12928 26292 12980
rect 27252 12928 27304 12980
rect 28908 12928 28960 12980
rect 29276 12928 29328 12980
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 19156 12860 19208 12912
rect 18236 12792 18288 12844
rect 18604 12792 18656 12844
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 18696 12724 18748 12776
rect 19156 12724 19208 12776
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 18328 12656 18380 12708
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 23756 12860 23808 12912
rect 20444 12656 20496 12708
rect 21364 12656 21416 12708
rect 23020 12792 23072 12844
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 24952 12860 25004 12912
rect 25228 12860 25280 12912
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 24308 12835 24360 12844
rect 23388 12767 23440 12776
rect 23388 12733 23397 12767
rect 23397 12733 23431 12767
rect 23431 12733 23440 12767
rect 23388 12724 23440 12733
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 27160 12792 27212 12844
rect 25044 12724 25096 12776
rect 25412 12724 25464 12776
rect 25872 12767 25924 12776
rect 25872 12733 25881 12767
rect 25881 12733 25915 12767
rect 25915 12733 25924 12767
rect 25872 12724 25924 12733
rect 29644 12835 29696 12844
rect 29644 12801 29653 12835
rect 29653 12801 29687 12835
rect 29687 12801 29696 12835
rect 29644 12792 29696 12801
rect 31852 12928 31904 12980
rect 34704 12928 34756 12980
rect 35348 12928 35400 12980
rect 35624 12928 35676 12980
rect 37096 12928 37148 12980
rect 37924 12928 37976 12980
rect 40500 12928 40552 12980
rect 43812 12928 43864 12980
rect 29828 12767 29880 12776
rect 29828 12733 29837 12767
rect 29837 12733 29871 12767
rect 29871 12733 29880 12767
rect 29828 12724 29880 12733
rect 30472 12724 30524 12776
rect 31760 12860 31812 12912
rect 31852 12792 31904 12844
rect 31760 12767 31812 12776
rect 31760 12733 31769 12767
rect 31769 12733 31803 12767
rect 31803 12733 31812 12767
rect 32496 12792 32548 12844
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 31760 12724 31812 12733
rect 24400 12656 24452 12708
rect 24492 12699 24544 12708
rect 24492 12665 24501 12699
rect 24501 12665 24535 12699
rect 24535 12665 24544 12699
rect 24492 12656 24544 12665
rect 16120 12588 16172 12640
rect 16672 12588 16724 12640
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 18788 12588 18840 12640
rect 19524 12588 19576 12640
rect 20536 12588 20588 12640
rect 22468 12631 22520 12640
rect 22468 12597 22477 12631
rect 22477 12597 22511 12631
rect 22511 12597 22520 12631
rect 22468 12588 22520 12597
rect 29000 12656 29052 12708
rect 31300 12656 31352 12708
rect 27620 12588 27672 12640
rect 30748 12588 30800 12640
rect 31576 12588 31628 12640
rect 31760 12588 31812 12640
rect 34704 12792 34756 12844
rect 34888 12792 34940 12844
rect 44364 12903 44416 12912
rect 44364 12869 44373 12903
rect 44373 12869 44407 12903
rect 44407 12869 44416 12903
rect 44364 12860 44416 12869
rect 40684 12767 40736 12776
rect 40684 12733 40693 12767
rect 40693 12733 40727 12767
rect 40727 12733 40736 12767
rect 40684 12724 40736 12733
rect 41328 12656 41380 12708
rect 44640 12656 44692 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12256 12384 12308 12436
rect 11980 12316 12032 12368
rect 13084 12384 13136 12436
rect 13176 12384 13228 12436
rect 14004 12384 14056 12436
rect 14096 12384 14148 12436
rect 14924 12384 14976 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15292 12384 15344 12436
rect 12440 12359 12492 12368
rect 12440 12325 12449 12359
rect 12449 12325 12483 12359
rect 12483 12325 12492 12359
rect 12440 12316 12492 12325
rect 13728 12316 13780 12368
rect 15200 12316 15252 12368
rect 15476 12384 15528 12436
rect 11612 12112 11664 12164
rect 11888 12112 11940 12164
rect 12532 12180 12584 12232
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 14004 12180 14056 12232
rect 14280 12180 14332 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 15108 12112 15160 12164
rect 15660 12316 15712 12368
rect 17040 12316 17092 12368
rect 16120 12248 16172 12300
rect 17316 12248 17368 12300
rect 20904 12384 20956 12436
rect 21180 12427 21232 12436
rect 21180 12393 21189 12427
rect 21189 12393 21223 12427
rect 21223 12393 21232 12427
rect 21180 12384 21232 12393
rect 22836 12384 22888 12436
rect 27712 12384 27764 12436
rect 29644 12384 29696 12436
rect 30748 12427 30800 12436
rect 30748 12393 30757 12427
rect 30757 12393 30791 12427
rect 30791 12393 30800 12427
rect 30748 12384 30800 12393
rect 19340 12316 19392 12368
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 16212 12180 16264 12232
rect 16488 12180 16540 12232
rect 16948 12180 17000 12232
rect 18604 12180 18656 12232
rect 19432 12248 19484 12300
rect 19524 12180 19576 12232
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 19984 12180 20036 12232
rect 20628 12316 20680 12368
rect 21364 12291 21416 12300
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 20260 12180 20312 12232
rect 20536 12223 20588 12232
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 20812 12180 20864 12232
rect 21732 12316 21784 12368
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 23756 12248 23808 12300
rect 22928 12180 22980 12232
rect 28356 12223 28408 12232
rect 28356 12189 28365 12223
rect 28365 12189 28399 12223
rect 28399 12189 28408 12223
rect 28356 12180 28408 12189
rect 29000 12180 29052 12232
rect 29092 12180 29144 12232
rect 29460 12180 29512 12232
rect 29920 12155 29972 12164
rect 29920 12121 29929 12155
rect 29929 12121 29963 12155
rect 29963 12121 29972 12155
rect 29920 12112 29972 12121
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 30656 12180 30708 12232
rect 32496 12384 32548 12436
rect 36084 12427 36136 12436
rect 36084 12393 36093 12427
rect 36093 12393 36127 12427
rect 36127 12393 36136 12427
rect 36084 12384 36136 12393
rect 31208 12180 31260 12232
rect 32404 12316 32456 12368
rect 34612 12316 34664 12368
rect 31392 12248 31444 12300
rect 31484 12180 31536 12232
rect 31668 12223 31720 12232
rect 31668 12189 31677 12223
rect 31677 12189 31711 12223
rect 31711 12189 31720 12223
rect 31668 12180 31720 12189
rect 31760 12180 31812 12232
rect 37464 12248 37516 12300
rect 37832 12291 37884 12300
rect 37832 12257 37841 12291
rect 37841 12257 37875 12291
rect 37875 12257 37884 12291
rect 37832 12248 37884 12257
rect 30748 12112 30800 12164
rect 31392 12112 31444 12164
rect 32128 12180 32180 12232
rect 32220 12223 32272 12232
rect 32220 12189 32229 12223
rect 32229 12189 32263 12223
rect 32263 12189 32272 12223
rect 32220 12180 32272 12189
rect 37004 12112 37056 12164
rect 39028 12112 39080 12164
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 12532 12044 12584 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 12900 12044 12952 12096
rect 13360 12044 13412 12096
rect 13452 12044 13504 12096
rect 14464 12044 14516 12096
rect 14924 12044 14976 12096
rect 15476 12044 15528 12096
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 18236 12044 18288 12096
rect 18512 12044 18564 12096
rect 18972 12044 19024 12096
rect 19340 12044 19392 12096
rect 20168 12044 20220 12096
rect 20628 12044 20680 12096
rect 22744 12044 22796 12096
rect 28816 12044 28868 12096
rect 30288 12044 30340 12096
rect 31208 12044 31260 12096
rect 34612 12044 34664 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 11704 11840 11756 11892
rect 12716 11840 12768 11892
rect 13912 11840 13964 11892
rect 14372 11840 14424 11892
rect 14740 11840 14792 11892
rect 15016 11840 15068 11892
rect 11428 11704 11480 11756
rect 11612 11636 11664 11688
rect 14556 11772 14608 11824
rect 15384 11840 15436 11892
rect 18420 11840 18472 11892
rect 18972 11840 19024 11892
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 12072 11636 12124 11688
rect 12808 11704 12860 11756
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 13820 11704 13872 11756
rect 14188 11704 14240 11756
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 14004 11636 14056 11688
rect 15292 11704 15344 11756
rect 16948 11704 17000 11756
rect 19156 11772 19208 11824
rect 19524 11840 19576 11892
rect 20076 11840 20128 11892
rect 20168 11840 20220 11892
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 23572 11840 23624 11892
rect 23940 11840 23992 11892
rect 25228 11883 25280 11892
rect 25228 11849 25237 11883
rect 25237 11849 25271 11883
rect 25271 11849 25280 11883
rect 25228 11840 25280 11849
rect 27068 11883 27120 11892
rect 27068 11849 27077 11883
rect 27077 11849 27111 11883
rect 27111 11849 27120 11883
rect 27068 11840 27120 11849
rect 29828 11840 29880 11892
rect 30564 11840 30616 11892
rect 13084 11568 13136 11620
rect 18604 11636 18656 11688
rect 19708 11747 19760 11756
rect 19708 11713 19717 11747
rect 19717 11713 19751 11747
rect 19751 11713 19760 11747
rect 19708 11704 19760 11713
rect 11704 11500 11756 11552
rect 13820 11500 13872 11552
rect 16120 11500 16172 11552
rect 17960 11500 18012 11552
rect 18328 11500 18380 11552
rect 18972 11568 19024 11620
rect 19340 11568 19392 11620
rect 20168 11704 20220 11756
rect 20628 11815 20680 11824
rect 20628 11781 20637 11815
rect 20637 11781 20671 11815
rect 20671 11781 20680 11815
rect 20628 11772 20680 11781
rect 27528 11815 27580 11824
rect 27528 11781 27537 11815
rect 27537 11781 27571 11815
rect 27571 11781 27580 11815
rect 27528 11772 27580 11781
rect 30380 11772 30432 11824
rect 20444 11704 20496 11756
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 25964 11747 26016 11756
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 27988 11704 28040 11756
rect 21180 11636 21232 11688
rect 24768 11636 24820 11688
rect 25412 11679 25464 11688
rect 25412 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25464 11679
rect 25412 11636 25464 11645
rect 26056 11679 26108 11688
rect 26056 11645 26065 11679
rect 26065 11645 26099 11679
rect 26099 11645 26108 11679
rect 26056 11636 26108 11645
rect 26148 11679 26200 11688
rect 26148 11645 26157 11679
rect 26157 11645 26191 11679
rect 26191 11645 26200 11679
rect 26148 11636 26200 11645
rect 27068 11636 27120 11688
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 30012 11636 30064 11688
rect 28816 11568 28868 11620
rect 30564 11747 30616 11756
rect 30564 11713 30573 11747
rect 30573 11713 30607 11747
rect 30607 11713 30616 11747
rect 30564 11704 30616 11713
rect 31024 11704 31076 11756
rect 31484 11747 31536 11756
rect 31484 11713 31493 11747
rect 31493 11713 31527 11747
rect 31527 11713 31536 11747
rect 31484 11704 31536 11713
rect 31852 11704 31904 11756
rect 32128 11704 32180 11756
rect 19984 11500 20036 11552
rect 26976 11500 27028 11552
rect 27252 11500 27304 11552
rect 28540 11543 28592 11552
rect 28540 11509 28549 11543
rect 28549 11509 28583 11543
rect 28583 11509 28592 11543
rect 28540 11500 28592 11509
rect 30104 11500 30156 11552
rect 31760 11636 31812 11688
rect 32220 11500 32272 11552
rect 35348 11772 35400 11824
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 37464 11704 37516 11756
rect 34428 11568 34480 11620
rect 37004 11568 37056 11620
rect 34704 11500 34756 11552
rect 35624 11500 35676 11552
rect 36452 11500 36504 11552
rect 36728 11500 36780 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12164 11296 12216 11348
rect 14648 11296 14700 11348
rect 16212 11296 16264 11348
rect 17960 11296 18012 11348
rect 19064 11296 19116 11348
rect 14464 11228 14516 11280
rect 15936 11228 15988 11280
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 23204 11296 23256 11348
rect 24860 11339 24912 11348
rect 24860 11305 24869 11339
rect 24869 11305 24903 11339
rect 24903 11305 24912 11339
rect 24860 11296 24912 11305
rect 25136 11296 25188 11348
rect 27528 11296 27580 11348
rect 28540 11296 28592 11348
rect 29000 11339 29052 11348
rect 29000 11305 29009 11339
rect 29009 11305 29043 11339
rect 29043 11305 29052 11339
rect 29000 11296 29052 11305
rect 30104 11296 30156 11348
rect 30564 11296 30616 11348
rect 31392 11296 31444 11348
rect 32220 11296 32272 11348
rect 17316 11160 17368 11212
rect 17500 11160 17552 11212
rect 13360 11092 13412 11144
rect 11428 11024 11480 11076
rect 14096 11024 14148 11076
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 15660 11092 15712 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 18236 11203 18288 11212
rect 18236 11169 18245 11203
rect 18245 11169 18279 11203
rect 18279 11169 18288 11203
rect 18236 11160 18288 11169
rect 23204 11160 23256 11212
rect 24676 11160 24728 11212
rect 17960 11092 18012 11144
rect 16120 11024 16172 11076
rect 12532 10956 12584 11008
rect 12992 10956 13044 11008
rect 16580 10956 16632 11008
rect 17224 10956 17276 11008
rect 17408 10956 17460 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 18144 11024 18196 11076
rect 18604 11024 18656 11076
rect 19340 11092 19392 11144
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 22652 11092 22704 11144
rect 24492 11092 24544 11144
rect 26148 11228 26200 11280
rect 27252 11160 27304 11212
rect 31300 11228 31352 11280
rect 31668 11228 31720 11280
rect 25320 11135 25372 11144
rect 25320 11101 25329 11135
rect 25329 11101 25363 11135
rect 25363 11101 25372 11135
rect 25320 11092 25372 11101
rect 19156 11024 19208 11076
rect 19064 10956 19116 11008
rect 23388 11024 23440 11076
rect 26056 11092 26108 11144
rect 28448 11160 28500 11212
rect 28908 11092 28960 11144
rect 29920 11092 29972 11144
rect 30748 11092 30800 11144
rect 31852 11203 31904 11212
rect 31852 11169 31861 11203
rect 31861 11169 31895 11203
rect 31895 11169 31904 11203
rect 31852 11160 31904 11169
rect 37372 11296 37424 11348
rect 38568 11228 38620 11280
rect 31300 11135 31352 11144
rect 31300 11101 31309 11135
rect 31309 11101 31343 11135
rect 31343 11101 31352 11135
rect 31300 11092 31352 11101
rect 31392 11135 31444 11144
rect 31392 11101 31401 11135
rect 31401 11101 31435 11135
rect 31435 11101 31444 11135
rect 31392 11092 31444 11101
rect 28264 11067 28316 11076
rect 28264 11033 28273 11067
rect 28273 11033 28307 11067
rect 28307 11033 28316 11067
rect 28264 11024 28316 11033
rect 32128 11135 32180 11144
rect 32128 11101 32137 11135
rect 32137 11101 32171 11135
rect 32171 11101 32180 11135
rect 32128 11092 32180 11101
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 37188 11160 37240 11212
rect 32404 11092 32456 11144
rect 34704 11135 34756 11144
rect 34704 11101 34713 11135
rect 34713 11101 34747 11135
rect 34747 11101 34756 11135
rect 34704 11092 34756 11101
rect 36360 11135 36412 11144
rect 36360 11101 36369 11135
rect 36369 11101 36403 11135
rect 36403 11101 36412 11135
rect 36360 11092 36412 11101
rect 38936 11135 38988 11144
rect 38936 11101 38945 11135
rect 38945 11101 38979 11135
rect 38979 11101 38988 11135
rect 38936 11092 38988 11101
rect 30748 10999 30800 11008
rect 30748 10965 30757 10999
rect 30757 10965 30791 10999
rect 30791 10965 30800 10999
rect 30748 10956 30800 10965
rect 30840 10956 30892 11008
rect 32496 11024 32548 11076
rect 36636 11067 36688 11076
rect 36636 11033 36645 11067
rect 36645 11033 36679 11067
rect 36679 11033 36688 11067
rect 36636 11024 36688 11033
rect 32128 10956 32180 11008
rect 35440 10999 35492 11008
rect 35440 10965 35449 10999
rect 35449 10965 35483 10999
rect 35483 10965 35492 10999
rect 35440 10956 35492 10965
rect 37004 10956 37056 11008
rect 38844 11024 38896 11076
rect 39120 10999 39172 11008
rect 39120 10965 39129 10999
rect 39129 10965 39163 10999
rect 39163 10965 39172 10999
rect 39120 10956 39172 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 12532 10752 12584 10804
rect 12716 10752 12768 10804
rect 11612 10616 11664 10668
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 12348 10548 12400 10600
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 15936 10752 15988 10804
rect 17224 10752 17276 10804
rect 18696 10752 18748 10804
rect 19156 10752 19208 10804
rect 19340 10752 19392 10804
rect 20536 10752 20588 10804
rect 22560 10795 22612 10804
rect 22560 10761 22569 10795
rect 22569 10761 22603 10795
rect 22603 10761 22612 10795
rect 22560 10752 22612 10761
rect 22652 10795 22704 10804
rect 22652 10761 22661 10795
rect 22661 10761 22695 10795
rect 22695 10761 22704 10795
rect 22652 10752 22704 10761
rect 24032 10752 24084 10804
rect 25320 10752 25372 10804
rect 26056 10752 26108 10804
rect 13084 10548 13136 10600
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 13636 10684 13688 10736
rect 13912 10548 13964 10600
rect 14832 10684 14884 10736
rect 15476 10684 15528 10736
rect 15752 10684 15804 10736
rect 14924 10616 14976 10668
rect 16304 10616 16356 10668
rect 17040 10684 17092 10736
rect 23020 10684 23072 10736
rect 23296 10684 23348 10736
rect 23756 10684 23808 10736
rect 23940 10684 23992 10736
rect 15200 10548 15252 10600
rect 15844 10548 15896 10600
rect 13728 10480 13780 10532
rect 11244 10412 11296 10464
rect 11796 10412 11848 10464
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 13544 10412 13596 10464
rect 13820 10412 13872 10464
rect 14556 10412 14608 10464
rect 14648 10412 14700 10464
rect 15384 10412 15436 10464
rect 16120 10412 16172 10464
rect 16304 10412 16356 10464
rect 16580 10548 16632 10600
rect 17500 10616 17552 10668
rect 18880 10616 18932 10668
rect 18972 10616 19024 10668
rect 22468 10616 22520 10668
rect 23572 10616 23624 10668
rect 23664 10659 23716 10668
rect 23664 10625 23673 10659
rect 23673 10625 23707 10659
rect 23707 10625 23716 10659
rect 23664 10616 23716 10625
rect 17224 10523 17276 10532
rect 17224 10489 17233 10523
rect 17233 10489 17267 10523
rect 17267 10489 17276 10523
rect 17224 10480 17276 10489
rect 18512 10480 18564 10532
rect 18880 10480 18932 10532
rect 19340 10480 19392 10532
rect 17960 10412 18012 10464
rect 19064 10412 19116 10464
rect 23480 10548 23532 10600
rect 29644 10752 29696 10804
rect 29828 10752 29880 10804
rect 31024 10795 31076 10804
rect 31024 10761 31033 10795
rect 31033 10761 31067 10795
rect 31067 10761 31076 10795
rect 31024 10752 31076 10761
rect 34704 10752 34756 10804
rect 36636 10752 36688 10804
rect 39120 10752 39172 10804
rect 26792 10616 26844 10668
rect 27068 10616 27120 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 27528 10659 27580 10668
rect 27528 10625 27561 10659
rect 27561 10625 27580 10659
rect 25412 10480 25464 10532
rect 26240 10591 26292 10600
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 27528 10616 27580 10625
rect 28080 10548 28132 10600
rect 26516 10480 26568 10532
rect 28264 10616 28316 10668
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 29092 10616 29144 10668
rect 29644 10616 29696 10668
rect 29920 10616 29972 10668
rect 30012 10659 30064 10668
rect 30012 10625 30021 10659
rect 30021 10625 30055 10659
rect 30055 10625 30064 10659
rect 30012 10616 30064 10625
rect 30104 10616 30156 10668
rect 31576 10684 31628 10736
rect 31668 10684 31720 10736
rect 31852 10684 31904 10736
rect 29184 10591 29236 10600
rect 29184 10557 29193 10591
rect 29193 10557 29227 10591
rect 29227 10557 29236 10591
rect 29184 10548 29236 10557
rect 29000 10480 29052 10532
rect 22100 10412 22152 10464
rect 22836 10455 22888 10464
rect 22836 10421 22845 10455
rect 22845 10421 22879 10455
rect 22879 10421 22888 10455
rect 22836 10412 22888 10421
rect 27528 10412 27580 10464
rect 28172 10455 28224 10464
rect 28172 10421 28181 10455
rect 28181 10421 28215 10455
rect 28215 10421 28224 10455
rect 28172 10412 28224 10421
rect 29276 10412 29328 10464
rect 29828 10412 29880 10464
rect 30840 10412 30892 10464
rect 31392 10616 31444 10668
rect 32036 10616 32088 10668
rect 34428 10684 34480 10736
rect 36452 10684 36504 10736
rect 31484 10480 31536 10532
rect 37372 10616 37424 10668
rect 38844 10616 38896 10668
rect 40684 10616 40736 10668
rect 37832 10591 37884 10600
rect 37832 10557 37841 10591
rect 37841 10557 37875 10591
rect 37875 10557 37884 10591
rect 37832 10548 37884 10557
rect 40224 10548 40276 10600
rect 31668 10455 31720 10464
rect 31668 10421 31677 10455
rect 31677 10421 31711 10455
rect 31711 10421 31720 10455
rect 31668 10412 31720 10421
rect 32220 10455 32272 10464
rect 32220 10421 32229 10455
rect 32229 10421 32263 10455
rect 32263 10421 32272 10455
rect 32220 10412 32272 10421
rect 34704 10412 34756 10464
rect 35348 10412 35400 10464
rect 38384 10455 38436 10464
rect 38384 10421 38393 10455
rect 38393 10421 38427 10455
rect 38427 10421 38436 10455
rect 38384 10412 38436 10421
rect 41236 10412 41288 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12256 10208 12308 10260
rect 12348 10208 12400 10260
rect 12164 10140 12216 10192
rect 12624 10208 12676 10260
rect 11520 10072 11572 10124
rect 15568 10208 15620 10260
rect 16856 10208 16908 10260
rect 19064 10208 19116 10260
rect 13084 10072 13136 10124
rect 14188 10072 14240 10124
rect 19432 10140 19484 10192
rect 11888 10047 11940 10056
rect 11888 10013 11906 10047
rect 11906 10013 11940 10047
rect 11888 10004 11940 10013
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 14280 10004 14332 10056
rect 14648 10004 14700 10056
rect 16120 10072 16172 10124
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 16672 10072 16724 10124
rect 16856 10072 16908 10124
rect 17868 10072 17920 10124
rect 20076 10208 20128 10260
rect 19984 10140 20036 10192
rect 16948 10004 17000 10056
rect 18052 10004 18104 10056
rect 20352 10140 20404 10192
rect 22744 10208 22796 10260
rect 22836 10208 22888 10260
rect 26792 10208 26844 10260
rect 23848 10072 23900 10124
rect 25412 10140 25464 10192
rect 25136 10072 25188 10124
rect 25780 10072 25832 10124
rect 26148 10072 26200 10124
rect 26516 10115 26568 10124
rect 26516 10081 26534 10115
rect 26534 10081 26568 10115
rect 26516 10072 26568 10081
rect 27160 10140 27212 10192
rect 27988 10208 28040 10260
rect 29000 10251 29052 10260
rect 29000 10217 29009 10251
rect 29009 10217 29043 10251
rect 29043 10217 29052 10251
rect 29000 10208 29052 10217
rect 29184 10251 29236 10260
rect 29184 10217 29193 10251
rect 29193 10217 29227 10251
rect 29227 10217 29236 10251
rect 29184 10208 29236 10217
rect 29276 10208 29328 10260
rect 31300 10208 31352 10260
rect 31392 10208 31444 10260
rect 31576 10251 31628 10260
rect 31576 10217 31585 10251
rect 31585 10217 31619 10251
rect 31619 10217 31628 10251
rect 31576 10208 31628 10217
rect 35348 10208 35400 10260
rect 36360 10208 36412 10260
rect 27252 10072 27304 10124
rect 30748 10140 30800 10192
rect 31208 10140 31260 10192
rect 12256 9868 12308 9920
rect 12532 9868 12584 9920
rect 12716 9868 12768 9920
rect 12808 9868 12860 9920
rect 14556 9868 14608 9920
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 16672 9868 16724 9877
rect 18972 9868 19024 9920
rect 19156 9868 19208 9920
rect 19984 9868 20036 9920
rect 20352 10004 20404 10056
rect 20444 10049 20496 10058
rect 20444 10015 20453 10049
rect 20453 10015 20487 10049
rect 20487 10015 20496 10049
rect 20444 10006 20496 10015
rect 20720 10004 20772 10056
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 27436 10004 27488 10056
rect 22560 9979 22612 9988
rect 22560 9945 22569 9979
rect 22569 9945 22603 9979
rect 22603 9945 22612 9979
rect 22560 9936 22612 9945
rect 20536 9868 20588 9920
rect 20996 9868 21048 9920
rect 22192 9868 22244 9920
rect 25596 9868 25648 9920
rect 29184 9936 29236 9988
rect 29460 9936 29512 9988
rect 30012 10004 30064 10056
rect 31300 10004 31352 10056
rect 31760 10047 31812 10056
rect 31760 10013 31769 10047
rect 31769 10013 31803 10047
rect 31803 10013 31812 10047
rect 31760 10004 31812 10013
rect 32128 10004 32180 10056
rect 35440 10140 35492 10192
rect 34612 10072 34664 10124
rect 40224 10208 40276 10260
rect 39212 10115 39264 10124
rect 39212 10081 39221 10115
rect 39221 10081 39255 10115
rect 39255 10081 39264 10115
rect 39212 10072 39264 10081
rect 41236 10072 41288 10124
rect 43628 10072 43680 10124
rect 39304 10047 39356 10056
rect 39304 10013 39313 10047
rect 39313 10013 39347 10047
rect 39347 10013 39356 10047
rect 39304 10004 39356 10013
rect 37280 9936 37332 9988
rect 37556 9979 37608 9988
rect 37556 9945 37565 9979
rect 37565 9945 37599 9979
rect 37599 9945 37608 9979
rect 37556 9936 37608 9945
rect 38844 9936 38896 9988
rect 29644 9868 29696 9920
rect 31300 9868 31352 9920
rect 31668 9868 31720 9920
rect 33968 9911 34020 9920
rect 33968 9877 33977 9911
rect 33977 9877 34011 9911
rect 34011 9877 34020 9911
rect 33968 9868 34020 9877
rect 34244 9911 34296 9920
rect 34244 9877 34253 9911
rect 34253 9877 34287 9911
rect 34287 9877 34296 9911
rect 34244 9868 34296 9877
rect 39028 9911 39080 9920
rect 39028 9877 39037 9911
rect 39037 9877 39071 9911
rect 39071 9877 39080 9911
rect 39028 9868 39080 9877
rect 39856 9911 39908 9920
rect 39856 9877 39865 9911
rect 39865 9877 39899 9911
rect 39899 9877 39908 9911
rect 39856 9868 39908 9877
rect 40868 9936 40920 9988
rect 43168 9979 43220 9988
rect 43168 9945 43177 9979
rect 43177 9945 43211 9979
rect 43211 9945 43220 9979
rect 43168 9936 43220 9945
rect 41696 9911 41748 9920
rect 41696 9877 41705 9911
rect 41705 9877 41739 9911
rect 41739 9877 41748 9911
rect 41696 9868 41748 9877
rect 42156 9868 42208 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 11980 9664 12032 9716
rect 11244 9460 11296 9512
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 16028 9707 16080 9716
rect 16028 9673 16037 9707
rect 16037 9673 16071 9707
rect 16071 9673 16080 9707
rect 16028 9664 16080 9673
rect 16212 9664 16264 9716
rect 16304 9664 16356 9716
rect 12348 9528 12400 9580
rect 12808 9528 12860 9580
rect 12992 9528 13044 9580
rect 14648 9596 14700 9648
rect 11428 9392 11480 9444
rect 12900 9460 12952 9512
rect 11796 9392 11848 9444
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13544 9528 13596 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 15292 9596 15344 9648
rect 13820 9460 13872 9512
rect 13912 9460 13964 9512
rect 14372 9460 14424 9512
rect 16212 9528 16264 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 18972 9639 19024 9648
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 16580 9460 16632 9512
rect 16396 9392 16448 9444
rect 11980 9324 12032 9376
rect 14004 9324 14056 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 14832 9324 14884 9376
rect 16580 9324 16632 9376
rect 16856 9324 16908 9376
rect 17408 9392 17460 9444
rect 18972 9605 18981 9639
rect 18981 9605 19015 9639
rect 19015 9605 19024 9639
rect 18972 9596 19024 9605
rect 19616 9664 19668 9716
rect 19800 9664 19852 9716
rect 20536 9664 20588 9716
rect 23480 9664 23532 9716
rect 23664 9664 23716 9716
rect 26792 9664 26844 9716
rect 27068 9664 27120 9716
rect 27344 9664 27396 9716
rect 28908 9664 28960 9716
rect 22376 9596 22428 9648
rect 18052 9528 18104 9580
rect 18512 9528 18564 9580
rect 18236 9392 18288 9444
rect 18696 9392 18748 9444
rect 18880 9460 18932 9512
rect 19984 9528 20036 9580
rect 19340 9460 19392 9512
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 22192 9528 22244 9580
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 23388 9528 23440 9580
rect 23572 9596 23624 9648
rect 23756 9528 23808 9580
rect 23940 9528 23992 9580
rect 26240 9460 26292 9512
rect 27252 9460 27304 9512
rect 25964 9392 26016 9444
rect 17592 9324 17644 9376
rect 18144 9324 18196 9376
rect 19156 9324 19208 9376
rect 19340 9324 19392 9376
rect 20076 9324 20128 9376
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 22468 9367 22520 9376
rect 22468 9333 22477 9367
rect 22477 9333 22511 9367
rect 22511 9333 22520 9367
rect 22468 9324 22520 9333
rect 23020 9324 23072 9376
rect 25688 9367 25740 9376
rect 25688 9333 25697 9367
rect 25697 9333 25731 9367
rect 25731 9333 25740 9367
rect 25688 9324 25740 9333
rect 28356 9596 28408 9648
rect 30196 9596 30248 9648
rect 31024 9664 31076 9716
rect 31484 9664 31536 9716
rect 32128 9664 32180 9716
rect 34428 9664 34480 9716
rect 37372 9664 37424 9716
rect 30012 9528 30064 9580
rect 30288 9528 30340 9580
rect 29644 9503 29696 9512
rect 29644 9469 29653 9503
rect 29653 9469 29687 9503
rect 29687 9469 29696 9503
rect 29644 9460 29696 9469
rect 29552 9392 29604 9444
rect 30656 9528 30708 9580
rect 31300 9571 31352 9580
rect 30564 9460 30616 9512
rect 31300 9537 31309 9571
rect 31309 9537 31343 9571
rect 31343 9537 31352 9571
rect 31300 9528 31352 9537
rect 31852 9528 31904 9580
rect 34704 9596 34756 9648
rect 39304 9664 39356 9716
rect 36820 9571 36872 9580
rect 34244 9460 34296 9512
rect 36820 9537 36829 9571
rect 36829 9537 36863 9571
rect 36863 9537 36872 9571
rect 36820 9528 36872 9537
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 37188 9528 37240 9580
rect 37556 9460 37608 9512
rect 37832 9460 37884 9512
rect 27436 9324 27488 9376
rect 27528 9324 27580 9376
rect 29920 9324 29972 9376
rect 30564 9324 30616 9376
rect 38384 9460 38436 9512
rect 38844 9528 38896 9580
rect 39120 9639 39172 9648
rect 39120 9605 39129 9639
rect 39129 9605 39163 9639
rect 39163 9605 39172 9639
rect 39120 9596 39172 9605
rect 41880 9639 41932 9648
rect 41880 9605 41907 9639
rect 41907 9605 41932 9639
rect 41880 9596 41932 9605
rect 43168 9664 43220 9716
rect 38568 9503 38620 9512
rect 38568 9469 38577 9503
rect 38577 9469 38611 9503
rect 38611 9469 38620 9503
rect 38568 9460 38620 9469
rect 39856 9460 39908 9512
rect 39028 9392 39080 9444
rect 42156 9528 42208 9580
rect 42708 9528 42760 9580
rect 42064 9392 42116 9444
rect 31392 9367 31444 9376
rect 31392 9333 31401 9367
rect 31401 9333 31435 9367
rect 31435 9333 31444 9367
rect 31392 9324 31444 9333
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 33140 9367 33192 9376
rect 33140 9333 33149 9367
rect 33149 9333 33183 9367
rect 33183 9333 33192 9367
rect 33140 9324 33192 9333
rect 39120 9324 39172 9376
rect 39304 9367 39356 9376
rect 39304 9333 39313 9367
rect 39313 9333 39347 9367
rect 39347 9333 39356 9367
rect 39304 9324 39356 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6920 9120 6972 9172
rect 11980 9120 12032 9172
rect 12808 9120 12860 9172
rect 13360 9120 13412 9172
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 14832 9120 14884 9172
rect 17132 9120 17184 9172
rect 12992 9052 13044 9104
rect 11520 8984 11572 9036
rect 940 8916 992 8968
rect 11796 8916 11848 8968
rect 12256 8916 12308 8968
rect 11704 8891 11756 8900
rect 11704 8857 11713 8891
rect 11713 8857 11747 8891
rect 11747 8857 11756 8891
rect 11704 8848 11756 8857
rect 13820 8916 13872 8968
rect 14004 8984 14056 9036
rect 14648 8984 14700 9036
rect 15660 9052 15712 9104
rect 16396 8984 16448 9036
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 13084 8780 13136 8832
rect 13728 8780 13780 8832
rect 13820 8780 13872 8832
rect 15844 8916 15896 8968
rect 16212 8916 16264 8968
rect 16488 8916 16540 8968
rect 16764 9052 16816 9104
rect 17776 9120 17828 9172
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 20352 9120 20404 9172
rect 22468 9120 22520 9172
rect 17960 9052 18012 9104
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 16672 8891 16724 8900
rect 16672 8857 16681 8891
rect 16681 8857 16715 8891
rect 16715 8857 16724 8891
rect 16672 8848 16724 8857
rect 14648 8780 14700 8832
rect 15936 8780 15988 8832
rect 16764 8780 16816 8832
rect 17408 8959 17460 8968
rect 17408 8925 17418 8959
rect 17418 8925 17460 8959
rect 17408 8916 17460 8925
rect 19984 8984 20036 9036
rect 17132 8848 17184 8900
rect 19524 8916 19576 8968
rect 22560 9052 22612 9104
rect 20628 8916 20680 8968
rect 22284 8916 22336 8968
rect 23388 9120 23440 9172
rect 25688 9120 25740 9172
rect 25780 9120 25832 9172
rect 27344 9163 27396 9172
rect 27344 9129 27353 9163
rect 27353 9129 27387 9163
rect 27387 9129 27396 9163
rect 27344 9120 27396 9129
rect 27528 9120 27580 9172
rect 28080 9163 28132 9172
rect 28080 9129 28089 9163
rect 28089 9129 28123 9163
rect 28123 9129 28132 9163
rect 28080 9120 28132 9129
rect 28448 9120 28500 9172
rect 30288 9163 30340 9172
rect 30288 9129 30297 9163
rect 30297 9129 30331 9163
rect 30331 9129 30340 9163
rect 30288 9120 30340 9129
rect 31392 9120 31444 9172
rect 31760 9120 31812 9172
rect 32404 9120 32456 9172
rect 33140 9120 33192 9172
rect 37372 9163 37424 9172
rect 37372 9129 37381 9163
rect 37381 9129 37415 9163
rect 37415 9129 37424 9163
rect 37372 9120 37424 9129
rect 38568 9120 38620 9172
rect 38936 9120 38988 9172
rect 39304 9120 39356 9172
rect 41880 9163 41932 9172
rect 41880 9129 41889 9163
rect 41889 9129 41923 9163
rect 41923 9129 41932 9163
rect 41880 9120 41932 9129
rect 23020 8959 23072 8968
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 23204 8959 23256 8968
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 26148 8984 26200 9036
rect 24400 8916 24452 8968
rect 25044 8959 25096 8968
rect 25044 8925 25053 8959
rect 25053 8925 25087 8959
rect 25087 8925 25096 8959
rect 27344 8984 27396 9036
rect 25044 8916 25096 8925
rect 27528 8959 27580 8968
rect 27528 8925 27537 8959
rect 27537 8925 27571 8959
rect 27571 8925 27580 8959
rect 27528 8916 27580 8925
rect 17040 8780 17092 8832
rect 17224 8780 17276 8832
rect 17592 8780 17644 8832
rect 20076 8891 20128 8900
rect 20076 8857 20085 8891
rect 20085 8857 20119 8891
rect 20119 8857 20128 8891
rect 20076 8848 20128 8857
rect 20536 8848 20588 8900
rect 22192 8848 22244 8900
rect 23756 8891 23808 8900
rect 23756 8857 23765 8891
rect 23765 8857 23799 8891
rect 23799 8857 23808 8891
rect 23756 8848 23808 8857
rect 25780 8848 25832 8900
rect 28172 8848 28224 8900
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 28540 8916 28592 8968
rect 30104 9052 30156 9104
rect 30840 9095 30892 9104
rect 30840 9061 30849 9095
rect 30849 9061 30883 9095
rect 30883 9061 30892 9095
rect 30840 9052 30892 9061
rect 29644 8916 29696 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 29828 8959 29880 8968
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 29828 8916 29880 8925
rect 28908 8891 28960 8900
rect 28908 8857 28935 8891
rect 28935 8857 28960 8891
rect 28908 8848 28960 8857
rect 29184 8848 29236 8900
rect 29920 8894 29972 8946
rect 30472 8984 30524 9036
rect 30196 8848 30248 8900
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 23388 8823 23440 8832
rect 23388 8789 23397 8823
rect 23397 8789 23431 8823
rect 23431 8789 23440 8823
rect 23388 8780 23440 8789
rect 25228 8780 25280 8832
rect 29000 8780 29052 8832
rect 29644 8780 29696 8832
rect 30288 8780 30340 8832
rect 30840 8848 30892 8900
rect 31576 8984 31628 9036
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 41696 8984 41748 9036
rect 31484 8848 31536 8900
rect 38384 8916 38436 8968
rect 42708 8984 42760 9036
rect 41972 8959 42024 8968
rect 41972 8925 41981 8959
rect 41981 8925 42015 8959
rect 42015 8925 42024 8959
rect 41972 8916 42024 8925
rect 42248 8916 42300 8968
rect 42616 8959 42668 8968
rect 42616 8925 42625 8959
rect 42625 8925 42659 8959
rect 42659 8925 42668 8959
rect 42616 8916 42668 8925
rect 42892 8916 42944 8968
rect 36912 8848 36964 8900
rect 39028 8848 39080 8900
rect 39488 8848 39540 8900
rect 42064 8848 42116 8900
rect 43076 8848 43128 8900
rect 31116 8780 31168 8832
rect 31576 8823 31628 8832
rect 31576 8789 31585 8823
rect 31585 8789 31619 8823
rect 31619 8789 31628 8823
rect 31576 8780 31628 8789
rect 31668 8823 31720 8832
rect 31668 8789 31677 8823
rect 31677 8789 31711 8823
rect 31711 8789 31720 8823
rect 31668 8780 31720 8789
rect 34152 8823 34204 8832
rect 34152 8789 34161 8823
rect 34161 8789 34195 8823
rect 34195 8789 34204 8823
rect 34152 8780 34204 8789
rect 36820 8780 36872 8832
rect 37096 8780 37148 8832
rect 39212 8780 39264 8832
rect 43352 8780 43404 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 11704 8576 11756 8628
rect 13728 8508 13780 8560
rect 14832 8508 14884 8560
rect 15660 8576 15712 8628
rect 15936 8576 15988 8628
rect 12532 8440 12584 8492
rect 14372 8440 14424 8492
rect 15108 8440 15160 8492
rect 16488 8508 16540 8560
rect 20076 8576 20128 8628
rect 22008 8576 22060 8628
rect 23388 8576 23440 8628
rect 24400 8619 24452 8628
rect 24400 8585 24409 8619
rect 24409 8585 24443 8619
rect 24443 8585 24452 8619
rect 24400 8576 24452 8585
rect 25044 8576 25096 8628
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 25596 8576 25648 8628
rect 26332 8576 26384 8628
rect 28172 8576 28224 8628
rect 28356 8576 28408 8628
rect 28448 8576 28500 8628
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 12164 8372 12216 8424
rect 12256 8372 12308 8424
rect 14556 8372 14608 8424
rect 17132 8440 17184 8492
rect 19892 8508 19944 8560
rect 20628 8508 20680 8560
rect 17592 8440 17644 8492
rect 26700 8440 26752 8492
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 29092 8576 29144 8628
rect 29644 8576 29696 8628
rect 29828 8576 29880 8628
rect 30840 8576 30892 8628
rect 31116 8576 31168 8628
rect 32128 8576 32180 8628
rect 34152 8576 34204 8628
rect 42248 8619 42300 8628
rect 15844 8372 15896 8424
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 18972 8372 19024 8424
rect 19616 8372 19668 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 22192 8372 22244 8424
rect 25320 8372 25372 8424
rect 25780 8415 25832 8424
rect 25780 8381 25789 8415
rect 25789 8381 25823 8415
rect 25823 8381 25832 8415
rect 25780 8372 25832 8381
rect 27252 8372 27304 8424
rect 27896 8372 27948 8424
rect 29000 8440 29052 8492
rect 29184 8483 29236 8492
rect 29184 8449 29193 8483
rect 29193 8449 29227 8483
rect 29227 8449 29236 8483
rect 29184 8440 29236 8449
rect 30012 8483 30064 8492
rect 30012 8449 30020 8483
rect 30020 8449 30054 8483
rect 30054 8449 30064 8483
rect 30012 8440 30064 8449
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 30288 8440 30340 8492
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 31024 8440 31076 8492
rect 37004 8508 37056 8560
rect 42248 8585 42257 8619
rect 42257 8585 42291 8619
rect 42291 8585 42300 8619
rect 42248 8576 42300 8585
rect 42616 8576 42668 8628
rect 31576 8483 31628 8492
rect 11428 8304 11480 8356
rect 14924 8304 14976 8356
rect 16764 8304 16816 8356
rect 23388 8304 23440 8356
rect 26424 8304 26476 8356
rect 17408 8236 17460 8288
rect 22284 8236 22336 8288
rect 27436 8304 27488 8356
rect 31576 8449 31585 8483
rect 31585 8449 31619 8483
rect 31619 8449 31628 8483
rect 31576 8440 31628 8449
rect 31760 8483 31812 8492
rect 31760 8449 31773 8483
rect 31773 8449 31812 8483
rect 31760 8440 31812 8449
rect 40408 8440 40460 8492
rect 41696 8508 41748 8560
rect 41972 8508 42024 8560
rect 40592 8483 40644 8492
rect 40592 8449 40601 8483
rect 40601 8449 40635 8483
rect 40635 8449 40644 8483
rect 40592 8440 40644 8449
rect 41420 8372 41472 8424
rect 31668 8304 31720 8356
rect 34244 8304 34296 8356
rect 43720 8415 43772 8424
rect 43720 8381 43729 8415
rect 43729 8381 43763 8415
rect 43763 8381 43772 8415
rect 43720 8372 43772 8381
rect 30472 8279 30524 8288
rect 30472 8245 30481 8279
rect 30481 8245 30515 8279
rect 30515 8245 30524 8279
rect 30472 8236 30524 8245
rect 31484 8279 31536 8288
rect 31484 8245 31493 8279
rect 31493 8245 31527 8279
rect 31527 8245 31536 8279
rect 31484 8236 31536 8245
rect 33600 8279 33652 8288
rect 33600 8245 33609 8279
rect 33609 8245 33643 8279
rect 33643 8245 33652 8279
rect 33600 8236 33652 8245
rect 36360 8236 36412 8288
rect 40316 8279 40368 8288
rect 40316 8245 40325 8279
rect 40325 8245 40359 8279
rect 40359 8245 40368 8279
rect 40316 8236 40368 8245
rect 41236 8236 41288 8288
rect 42064 8279 42116 8288
rect 42064 8245 42073 8279
rect 42073 8245 42107 8279
rect 42107 8245 42116 8279
rect 42064 8236 42116 8245
rect 42432 8279 42484 8288
rect 42432 8245 42441 8279
rect 42441 8245 42475 8279
rect 42475 8245 42484 8279
rect 42432 8236 42484 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 12072 8032 12124 8084
rect 12624 8007 12676 8016
rect 12624 7973 12633 8007
rect 12633 7973 12667 8007
rect 12667 7973 12676 8007
rect 12624 7964 12676 7973
rect 11612 7896 11664 7948
rect 11796 7803 11848 7812
rect 11796 7769 11805 7803
rect 11805 7769 11839 7803
rect 11839 7769 11848 7803
rect 11796 7760 11848 7769
rect 11980 7760 12032 7812
rect 13268 8032 13320 8084
rect 13728 8032 13780 8084
rect 18788 8032 18840 8084
rect 19524 8032 19576 8084
rect 20076 8032 20128 8084
rect 19616 7964 19668 8016
rect 13268 7896 13320 7948
rect 15476 7896 15528 7948
rect 19432 7896 19484 7948
rect 19892 7896 19944 7948
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12716 7828 12768 7880
rect 16580 7828 16632 7880
rect 17684 7828 17736 7880
rect 13176 7760 13228 7812
rect 18144 7828 18196 7880
rect 11244 7692 11296 7744
rect 12256 7692 12308 7744
rect 14832 7692 14884 7744
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 18328 7692 18380 7744
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 23296 8075 23348 8084
rect 23296 8041 23305 8075
rect 23305 8041 23339 8075
rect 23339 8041 23348 8075
rect 23296 8032 23348 8041
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 25596 8032 25648 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 29736 8075 29788 8084
rect 29736 8041 29745 8075
rect 29745 8041 29779 8075
rect 29779 8041 29788 8075
rect 29736 8032 29788 8041
rect 30196 8032 30248 8084
rect 31024 8032 31076 8084
rect 19340 7760 19392 7812
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 20444 7828 20496 7880
rect 22100 7828 22152 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 27344 7964 27396 8016
rect 36636 7964 36688 8016
rect 27528 7896 27580 7948
rect 29092 7896 29144 7948
rect 21456 7803 21508 7812
rect 21456 7769 21465 7803
rect 21465 7769 21499 7803
rect 21499 7769 21508 7803
rect 21456 7760 21508 7769
rect 21548 7760 21600 7812
rect 27896 7871 27948 7880
rect 27896 7837 27905 7871
rect 27905 7837 27939 7871
rect 27939 7837 27948 7871
rect 27896 7828 27948 7837
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 27344 7760 27396 7812
rect 34704 7939 34756 7948
rect 34704 7905 34713 7939
rect 34713 7905 34747 7939
rect 34747 7905 34756 7939
rect 34704 7896 34756 7905
rect 20352 7692 20404 7744
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 24400 7692 24452 7744
rect 28080 7692 28132 7744
rect 30472 7760 30524 7812
rect 31484 7828 31536 7880
rect 31576 7828 31628 7880
rect 34980 7803 35032 7812
rect 34980 7769 34989 7803
rect 34989 7769 35023 7803
rect 35023 7769 35032 7803
rect 34980 7760 35032 7769
rect 36360 7760 36412 7812
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 36912 7828 36964 7880
rect 37740 7828 37792 7880
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 40316 8032 40368 8084
rect 42064 8032 42116 8084
rect 37096 7760 37148 7812
rect 38660 7760 38712 7812
rect 36544 7692 36596 7744
rect 36820 7735 36872 7744
rect 36820 7701 36829 7735
rect 36829 7701 36863 7735
rect 36863 7701 36872 7735
rect 36820 7692 36872 7701
rect 37464 7735 37516 7744
rect 37464 7701 37473 7735
rect 37473 7701 37507 7735
rect 37507 7701 37516 7735
rect 37464 7692 37516 7701
rect 37556 7735 37608 7744
rect 37556 7701 37565 7735
rect 37565 7701 37599 7735
rect 37599 7701 37608 7735
rect 37556 7692 37608 7701
rect 38752 7692 38804 7744
rect 41236 7828 41288 7880
rect 40224 7692 40276 7744
rect 41420 7692 41472 7744
rect 43628 7871 43680 7880
rect 43628 7837 43637 7871
rect 43637 7837 43671 7871
rect 43671 7837 43680 7871
rect 43628 7828 43680 7837
rect 43076 7760 43128 7812
rect 43444 7760 43496 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 12072 7488 12124 7540
rect 12532 7488 12584 7540
rect 13268 7531 13320 7540
rect 13268 7497 13298 7531
rect 13298 7497 13320 7531
rect 13268 7488 13320 7497
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 13084 7463 13136 7472
rect 13084 7429 13093 7463
rect 13093 7429 13127 7463
rect 13127 7429 13136 7463
rect 13084 7420 13136 7429
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 11704 7352 11756 7404
rect 12072 7352 12124 7404
rect 12256 7352 12308 7404
rect 14280 7420 14332 7472
rect 14832 7531 14884 7540
rect 14832 7497 14841 7531
rect 14841 7497 14875 7531
rect 14875 7497 14884 7531
rect 14832 7488 14884 7497
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 17684 7488 17736 7540
rect 15752 7420 15804 7472
rect 13360 7216 13412 7268
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14740 7352 14792 7404
rect 14924 7352 14976 7404
rect 17040 7327 17092 7336
rect 17040 7293 17049 7327
rect 17049 7293 17083 7327
rect 17083 7293 17092 7327
rect 17040 7284 17092 7293
rect 14832 7216 14884 7268
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 18328 7352 18380 7404
rect 18972 7420 19024 7472
rect 19340 7420 19392 7472
rect 19984 7488 20036 7540
rect 20536 7488 20588 7540
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 20352 7463 20404 7472
rect 20352 7429 20361 7463
rect 20361 7429 20395 7463
rect 20395 7429 20404 7463
rect 20352 7420 20404 7429
rect 20260 7352 20312 7404
rect 17960 7216 18012 7268
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 13176 7148 13228 7200
rect 15752 7148 15804 7200
rect 16304 7148 16356 7200
rect 19984 7284 20036 7336
rect 24584 7488 24636 7540
rect 25320 7488 25372 7540
rect 26884 7488 26936 7540
rect 27344 7531 27396 7540
rect 27344 7497 27353 7531
rect 27353 7497 27387 7531
rect 27387 7497 27396 7531
rect 27344 7488 27396 7497
rect 27896 7488 27948 7540
rect 34980 7488 35032 7540
rect 36636 7488 36688 7540
rect 36728 7488 36780 7540
rect 37280 7488 37332 7540
rect 23848 7420 23900 7472
rect 21088 7327 21140 7336
rect 21088 7293 21097 7327
rect 21097 7293 21131 7327
rect 21131 7293 21140 7327
rect 21088 7284 21140 7293
rect 21180 7216 21232 7268
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 24860 7395 24912 7404
rect 24860 7361 24869 7395
rect 24869 7361 24903 7395
rect 24903 7361 24912 7395
rect 24860 7352 24912 7361
rect 25964 7352 26016 7404
rect 23572 7284 23624 7336
rect 24400 7284 24452 7336
rect 25872 7284 25924 7336
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 38752 7420 38804 7472
rect 39212 7420 39264 7472
rect 20168 7148 20220 7200
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 36912 7395 36964 7404
rect 36912 7361 36921 7395
rect 36921 7361 36955 7395
rect 36955 7361 36964 7395
rect 36912 7352 36964 7361
rect 37004 7352 37056 7404
rect 37372 7352 37424 7404
rect 39120 7395 39172 7404
rect 39120 7361 39129 7395
rect 39129 7361 39163 7395
rect 39163 7361 39172 7395
rect 39120 7352 39172 7361
rect 39580 7352 39632 7404
rect 40224 7463 40276 7472
rect 40224 7429 40233 7463
rect 40233 7429 40267 7463
rect 40267 7429 40276 7463
rect 40224 7420 40276 7429
rect 41696 7488 41748 7540
rect 42248 7488 42300 7540
rect 43628 7488 43680 7540
rect 37556 7284 37608 7336
rect 38752 7327 38804 7336
rect 38752 7293 38761 7327
rect 38761 7293 38795 7327
rect 38795 7293 38804 7327
rect 38752 7284 38804 7293
rect 39028 7327 39080 7336
rect 39028 7293 39037 7327
rect 39037 7293 39071 7327
rect 39071 7293 39080 7327
rect 39028 7284 39080 7293
rect 40408 7395 40460 7404
rect 40408 7361 40417 7395
rect 40417 7361 40451 7395
rect 40451 7361 40460 7395
rect 40408 7352 40460 7361
rect 41328 7395 41380 7404
rect 41328 7361 41337 7395
rect 41337 7361 41371 7395
rect 41371 7361 41380 7395
rect 41328 7352 41380 7361
rect 41420 7284 41472 7336
rect 37648 7216 37700 7268
rect 39672 7216 39724 7268
rect 37740 7148 37792 7200
rect 39488 7148 39540 7200
rect 41788 7395 41840 7404
rect 41788 7361 41797 7395
rect 41797 7361 41831 7395
rect 41831 7361 41840 7395
rect 41788 7352 41840 7361
rect 42064 7352 42116 7404
rect 42248 7395 42300 7404
rect 42248 7361 42257 7395
rect 42257 7361 42291 7395
rect 42291 7361 42300 7395
rect 42248 7352 42300 7361
rect 42432 7395 42484 7404
rect 42432 7361 42441 7395
rect 42441 7361 42475 7395
rect 42475 7361 42484 7395
rect 42432 7352 42484 7361
rect 42708 7395 42760 7404
rect 42708 7361 42717 7395
rect 42717 7361 42751 7395
rect 42751 7361 42760 7395
rect 42708 7352 42760 7361
rect 43720 7216 43772 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6920 6944 6972 6996
rect 11612 6944 11664 6996
rect 11704 6944 11756 6996
rect 15936 6944 15988 6996
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9772 6740 9824 6792
rect 11336 6740 11388 6792
rect 12716 6876 12768 6928
rect 15016 6876 15068 6928
rect 13176 6808 13228 6860
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 15200 6808 15252 6860
rect 16028 6808 16080 6860
rect 7288 6672 7340 6724
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14372 6740 14424 6792
rect 14648 6783 14700 6792
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 15660 6783 15712 6792
rect 12348 6715 12400 6724
rect 12348 6681 12357 6715
rect 12357 6681 12391 6715
rect 12391 6681 12400 6715
rect 12348 6672 12400 6681
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 6368 6604 6420 6613
rect 9588 6604 9640 6656
rect 11796 6604 11848 6656
rect 12256 6604 12308 6656
rect 13544 6604 13596 6656
rect 13820 6672 13872 6724
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16212 6783 16264 6792
rect 16212 6749 16243 6783
rect 16243 6749 16264 6783
rect 16212 6740 16264 6749
rect 15292 6604 15344 6656
rect 15660 6604 15712 6656
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 17224 6944 17276 6996
rect 17776 6944 17828 6996
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 21088 6944 21140 6996
rect 21456 6944 21508 6996
rect 23572 6944 23624 6996
rect 23848 6944 23900 6996
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 17408 6740 17460 6792
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 17408 6604 17460 6656
rect 18604 6672 18656 6724
rect 20260 6783 20312 6792
rect 20260 6749 20294 6783
rect 20294 6749 20312 6783
rect 20260 6740 20312 6749
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 23572 6808 23624 6860
rect 25044 6944 25096 6996
rect 25320 6944 25372 6996
rect 27252 6944 27304 6996
rect 33600 6944 33652 6996
rect 36820 6944 36872 6996
rect 37372 6944 37424 6996
rect 39304 6944 39356 6996
rect 19156 6604 19208 6656
rect 24308 6740 24360 6792
rect 24400 6740 24452 6792
rect 42800 6919 42852 6928
rect 42800 6885 42809 6919
rect 42809 6885 42843 6919
rect 42843 6885 42852 6919
rect 42800 6876 42852 6885
rect 43536 6944 43588 6996
rect 25780 6808 25832 6860
rect 25872 6808 25924 6860
rect 24860 6672 24912 6724
rect 25964 6740 26016 6792
rect 31024 6808 31076 6860
rect 37464 6808 37516 6860
rect 37556 6851 37608 6860
rect 37556 6817 37565 6851
rect 37565 6817 37599 6851
rect 37599 6817 37608 6851
rect 37556 6808 37608 6817
rect 42708 6808 42760 6860
rect 42892 6851 42944 6860
rect 42892 6817 42901 6851
rect 42901 6817 42935 6851
rect 42935 6817 42944 6851
rect 42892 6808 42944 6817
rect 43076 6851 43128 6860
rect 43076 6817 43085 6851
rect 43085 6817 43119 6851
rect 43119 6817 43128 6851
rect 43076 6808 43128 6817
rect 43352 6851 43404 6860
rect 43352 6817 43361 6851
rect 43361 6817 43395 6851
rect 43395 6817 43404 6851
rect 43352 6808 43404 6817
rect 27068 6740 27120 6792
rect 23480 6604 23532 6656
rect 24768 6604 24820 6656
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 27528 6740 27580 6792
rect 34520 6740 34572 6792
rect 37924 6740 37976 6792
rect 39120 6740 39172 6792
rect 39672 6740 39724 6792
rect 31208 6715 31260 6724
rect 31208 6681 31217 6715
rect 31217 6681 31251 6715
rect 31251 6681 31260 6715
rect 31208 6672 31260 6681
rect 36360 6672 36412 6724
rect 36728 6672 36780 6724
rect 37004 6672 37056 6724
rect 39580 6715 39632 6724
rect 39580 6681 39589 6715
rect 39589 6681 39623 6715
rect 39623 6681 39632 6715
rect 39580 6672 39632 6681
rect 43444 6672 43496 6724
rect 25044 6604 25096 6613
rect 30196 6604 30248 6656
rect 31024 6647 31076 6656
rect 31024 6613 31033 6647
rect 31033 6613 31067 6647
rect 31067 6613 31076 6647
rect 31024 6604 31076 6613
rect 32220 6604 32272 6656
rect 33048 6604 33100 6656
rect 38200 6647 38252 6656
rect 38200 6613 38209 6647
rect 38209 6613 38243 6647
rect 38243 6613 38252 6647
rect 38200 6604 38252 6613
rect 38292 6647 38344 6656
rect 38292 6613 38301 6647
rect 38301 6613 38335 6647
rect 38335 6613 38344 6647
rect 38292 6604 38344 6613
rect 39212 6604 39264 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5724 6400 5776 6452
rect 6368 6400 6420 6452
rect 9496 6400 9548 6452
rect 13360 6400 13412 6452
rect 15292 6400 15344 6452
rect 5448 6332 5500 6384
rect 7288 6332 7340 6384
rect 13268 6332 13320 6384
rect 9588 6264 9640 6316
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 13820 6264 13872 6316
rect 15200 6375 15252 6384
rect 15200 6341 15209 6375
rect 15209 6341 15243 6375
rect 15243 6341 15252 6375
rect 15200 6332 15252 6341
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 3792 6060 3844 6112
rect 6920 6196 6972 6248
rect 8208 6196 8260 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 12164 6196 12216 6248
rect 10324 6060 10376 6112
rect 14096 6196 14148 6248
rect 14372 6196 14424 6248
rect 14740 6264 14792 6316
rect 14832 6264 14884 6316
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 15476 6264 15528 6316
rect 15936 6264 15988 6316
rect 16028 6264 16080 6316
rect 16488 6264 16540 6316
rect 13360 6171 13412 6180
rect 13360 6137 13369 6171
rect 13369 6137 13403 6171
rect 13403 6137 13412 6171
rect 13360 6128 13412 6137
rect 13452 6171 13504 6180
rect 13452 6137 13461 6171
rect 13461 6137 13495 6171
rect 13495 6137 13504 6171
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 17684 6400 17736 6452
rect 20260 6400 20312 6452
rect 17500 6375 17552 6384
rect 17500 6341 17509 6375
rect 17509 6341 17543 6375
rect 17543 6341 17552 6375
rect 17500 6332 17552 6341
rect 17132 6307 17184 6316
rect 17132 6273 17141 6307
rect 17141 6273 17175 6307
rect 17175 6273 17184 6307
rect 17132 6264 17184 6273
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 18512 6332 18564 6384
rect 19432 6332 19484 6384
rect 20444 6332 20496 6384
rect 18420 6196 18472 6248
rect 13452 6128 13504 6137
rect 14096 6060 14148 6112
rect 14740 6060 14792 6112
rect 15384 6060 15436 6112
rect 19156 6264 19208 6316
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 18880 6196 18932 6248
rect 19064 6128 19116 6180
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 23572 6307 23624 6316
rect 23572 6273 23581 6307
rect 23581 6273 23615 6307
rect 23615 6273 23624 6307
rect 23572 6264 23624 6273
rect 24308 6332 24360 6384
rect 33876 6400 33928 6452
rect 33968 6400 34020 6452
rect 36912 6400 36964 6452
rect 37924 6443 37976 6452
rect 24400 6307 24452 6316
rect 24400 6273 24409 6307
rect 24409 6273 24443 6307
rect 24443 6273 24452 6307
rect 24400 6264 24452 6273
rect 24768 6264 24820 6316
rect 30380 6264 30432 6316
rect 24860 6128 24912 6180
rect 15936 6060 15988 6112
rect 18604 6060 18656 6112
rect 19432 6060 19484 6112
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 23940 6060 23992 6112
rect 25044 6060 25096 6112
rect 25228 6103 25280 6112
rect 25228 6069 25237 6103
rect 25237 6069 25271 6103
rect 25271 6069 25280 6103
rect 25228 6060 25280 6069
rect 29460 6239 29512 6248
rect 29460 6205 29469 6239
rect 29469 6205 29503 6239
rect 29503 6205 29512 6239
rect 29460 6196 29512 6205
rect 30196 6239 30248 6248
rect 30196 6205 30205 6239
rect 30205 6205 30239 6239
rect 30239 6205 30248 6239
rect 30196 6196 30248 6205
rect 31668 6239 31720 6248
rect 31668 6205 31677 6239
rect 31677 6205 31711 6239
rect 31711 6205 31720 6239
rect 31668 6196 31720 6205
rect 26148 6060 26200 6112
rect 29552 6060 29604 6112
rect 29920 6060 29972 6112
rect 34520 6264 34572 6316
rect 37096 6375 37148 6384
rect 37096 6341 37105 6375
rect 37105 6341 37139 6375
rect 37139 6341 37148 6375
rect 37096 6332 37148 6341
rect 37648 6375 37700 6384
rect 37648 6341 37657 6375
rect 37657 6341 37691 6375
rect 37691 6341 37700 6375
rect 37648 6332 37700 6341
rect 37924 6409 37926 6443
rect 37926 6409 37960 6443
rect 37960 6409 37976 6443
rect 37924 6400 37976 6409
rect 38200 6400 38252 6452
rect 38292 6400 38344 6452
rect 41788 6400 41840 6452
rect 42708 6400 42760 6452
rect 42800 6400 42852 6452
rect 44640 6443 44692 6452
rect 44640 6409 44649 6443
rect 44649 6409 44683 6443
rect 44683 6409 44692 6443
rect 44640 6400 44692 6409
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 37464 6196 37516 6248
rect 37648 6196 37700 6248
rect 42248 6264 42300 6316
rect 38660 6196 38712 6248
rect 38752 6196 38804 6248
rect 42892 6264 42944 6316
rect 45284 6332 45336 6384
rect 32220 6060 32272 6112
rect 33140 6060 33192 6112
rect 36544 6060 36596 6112
rect 42984 6171 43036 6180
rect 42984 6137 42993 6171
rect 42993 6137 43027 6171
rect 43027 6137 43036 6171
rect 42984 6128 43036 6137
rect 37556 6060 37608 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5908 5856 5960 5908
rect 3240 5652 3292 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 5448 5584 5500 5636
rect 7288 5856 7340 5908
rect 8576 5856 8628 5908
rect 11980 5856 12032 5908
rect 14372 5856 14424 5908
rect 15384 5899 15436 5908
rect 15384 5865 15393 5899
rect 15393 5865 15427 5899
rect 15427 5865 15436 5899
rect 15384 5856 15436 5865
rect 6920 5720 6972 5772
rect 9588 5788 9640 5840
rect 12256 5788 12308 5840
rect 14004 5788 14056 5840
rect 14096 5788 14148 5840
rect 16948 5856 17000 5908
rect 18236 5856 18288 5908
rect 19248 5856 19300 5908
rect 20812 5856 20864 5908
rect 23756 5856 23808 5908
rect 23848 5856 23900 5908
rect 25228 5856 25280 5908
rect 26148 5856 26200 5908
rect 13360 5720 13412 5772
rect 14648 5720 14700 5772
rect 15292 5720 15344 5772
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 13636 5652 13688 5704
rect 7564 5584 7616 5636
rect 9680 5584 9732 5636
rect 10968 5584 11020 5636
rect 13084 5584 13136 5636
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 14004 5652 14056 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 15200 5652 15252 5704
rect 17592 5720 17644 5772
rect 16212 5695 16264 5704
rect 15568 5584 15620 5636
rect 9772 5516 9824 5568
rect 15108 5516 15160 5568
rect 15200 5516 15252 5568
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16488 5652 16540 5704
rect 16028 5584 16080 5636
rect 17408 5584 17460 5636
rect 17592 5627 17644 5636
rect 17592 5593 17601 5627
rect 17601 5593 17635 5627
rect 17635 5593 17644 5627
rect 17592 5584 17644 5593
rect 24308 5788 24360 5840
rect 21180 5652 21232 5704
rect 23940 5652 23992 5704
rect 24124 5652 24176 5704
rect 24400 5652 24452 5704
rect 25504 5695 25556 5704
rect 25504 5661 25513 5695
rect 25513 5661 25547 5695
rect 25547 5661 25556 5695
rect 25504 5652 25556 5661
rect 27068 5652 27120 5704
rect 29000 5652 29052 5704
rect 23572 5516 23624 5568
rect 24308 5516 24360 5568
rect 27344 5584 27396 5636
rect 25504 5516 25556 5568
rect 26148 5516 26200 5568
rect 27160 5516 27212 5568
rect 29460 5856 29512 5908
rect 31024 5856 31076 5908
rect 31208 5856 31260 5908
rect 31668 5856 31720 5908
rect 32312 5899 32364 5908
rect 32312 5865 32321 5899
rect 32321 5865 32355 5899
rect 32355 5865 32364 5899
rect 32312 5856 32364 5865
rect 33048 5856 33100 5908
rect 33140 5856 33192 5908
rect 29920 5720 29972 5772
rect 29552 5695 29604 5704
rect 29552 5661 29561 5695
rect 29561 5661 29595 5695
rect 29595 5661 29604 5695
rect 29552 5652 29604 5661
rect 31208 5652 31260 5704
rect 31576 5695 31628 5704
rect 31576 5661 31585 5695
rect 31585 5661 31619 5695
rect 31619 5661 31628 5695
rect 31576 5652 31628 5661
rect 31668 5652 31720 5704
rect 33876 5856 33928 5908
rect 39580 5856 39632 5908
rect 43076 5763 43128 5772
rect 43076 5729 43085 5763
rect 43085 5729 43119 5763
rect 43119 5729 43128 5763
rect 43076 5720 43128 5729
rect 37372 5652 37424 5704
rect 38016 5695 38068 5704
rect 38016 5661 38025 5695
rect 38025 5661 38059 5695
rect 38059 5661 38068 5695
rect 38016 5652 38068 5661
rect 30380 5584 30432 5636
rect 43352 5627 43404 5636
rect 43352 5593 43361 5627
rect 43361 5593 43395 5627
rect 43395 5593 43404 5627
rect 43352 5584 43404 5593
rect 43444 5584 43496 5636
rect 44824 5559 44876 5568
rect 44824 5525 44833 5559
rect 44833 5525 44867 5559
rect 44867 5525 44876 5559
rect 44824 5516 44876 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2688 5312 2740 5364
rect 4160 5312 4212 5364
rect 6920 5312 6972 5364
rect 10048 5312 10100 5364
rect 10416 5312 10468 5364
rect 13636 5312 13688 5364
rect 14832 5312 14884 5364
rect 9588 5244 9640 5296
rect 13912 5244 13964 5296
rect 15568 5244 15620 5296
rect 20076 5312 20128 5364
rect 19984 5244 20036 5296
rect 5448 5176 5500 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10600 5176 10652 5228
rect 10968 5108 11020 5160
rect 12624 5176 12676 5228
rect 17040 5176 17092 5228
rect 13176 5108 13228 5160
rect 19156 5108 19208 5160
rect 22192 5176 22244 5228
rect 20812 5108 20864 5160
rect 21272 5151 21324 5160
rect 21272 5117 21281 5151
rect 21281 5117 21315 5151
rect 21315 5117 21324 5151
rect 21272 5108 21324 5117
rect 22100 5108 22152 5160
rect 23296 5108 23348 5160
rect 18144 5040 18196 5092
rect 23112 5040 23164 5092
rect 23848 5108 23900 5160
rect 3240 4972 3292 5024
rect 8300 4972 8352 5024
rect 11980 5015 12032 5024
rect 11980 4981 11989 5015
rect 11989 4981 12023 5015
rect 12023 4981 12032 5015
rect 11980 4972 12032 4981
rect 14096 4972 14148 5024
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 20352 4972 20404 5024
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 24124 5040 24176 5092
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 24860 5176 24912 5228
rect 25228 5040 25280 5092
rect 23756 4972 23808 5024
rect 23848 5015 23900 5024
rect 23848 4981 23857 5015
rect 23857 4981 23891 5015
rect 23891 4981 23900 5015
rect 23848 4972 23900 4981
rect 24492 5015 24544 5024
rect 24492 4981 24501 5015
rect 24501 4981 24535 5015
rect 24535 4981 24544 5015
rect 24492 4972 24544 4981
rect 25412 5176 25464 5228
rect 26148 5176 26200 5228
rect 25504 5151 25556 5160
rect 25504 5117 25513 5151
rect 25513 5117 25547 5151
rect 25547 5117 25556 5151
rect 25504 5108 25556 5117
rect 25872 5040 25924 5092
rect 25964 5040 26016 5092
rect 26976 5312 27028 5364
rect 31576 5312 31628 5364
rect 35348 5312 35400 5364
rect 38752 5312 38804 5364
rect 41328 5312 41380 5364
rect 42156 5355 42208 5364
rect 42156 5321 42165 5355
rect 42165 5321 42199 5355
rect 42199 5321 42208 5355
rect 42156 5312 42208 5321
rect 29736 5244 29788 5296
rect 30288 5244 30340 5296
rect 37280 5287 37332 5296
rect 26976 5176 27028 5228
rect 37280 5253 37289 5287
rect 37289 5253 37323 5287
rect 37323 5253 37332 5287
rect 37280 5244 37332 5253
rect 34612 5176 34664 5228
rect 35440 5176 35492 5228
rect 29552 5151 29604 5160
rect 29552 5117 29561 5151
rect 29561 5117 29595 5151
rect 29595 5117 29604 5151
rect 29552 5108 29604 5117
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 31300 5108 31352 5160
rect 36544 5176 36596 5228
rect 36728 5176 36780 5228
rect 38752 5176 38804 5228
rect 39028 5176 39080 5228
rect 39212 5176 39264 5228
rect 27344 5083 27396 5092
rect 27344 5049 27353 5083
rect 27353 5049 27387 5083
rect 27387 5049 27396 5083
rect 27344 5040 27396 5049
rect 29000 5040 29052 5092
rect 36084 5151 36136 5160
rect 36084 5117 36093 5151
rect 36093 5117 36127 5151
rect 36127 5117 36136 5151
rect 36084 5108 36136 5117
rect 41512 5176 41564 5228
rect 42248 5219 42300 5228
rect 39580 5151 39632 5160
rect 39580 5117 39589 5151
rect 39589 5117 39623 5151
rect 39623 5117 39632 5151
rect 39580 5108 39632 5117
rect 41052 5151 41104 5160
rect 41052 5117 41061 5151
rect 41061 5117 41095 5151
rect 41095 5117 41104 5151
rect 41052 5108 41104 5117
rect 36452 5040 36504 5092
rect 41696 5040 41748 5092
rect 42248 5185 42257 5219
rect 42257 5185 42291 5219
rect 42291 5185 42300 5219
rect 42248 5176 42300 5185
rect 43352 5312 43404 5364
rect 42892 5108 42944 5160
rect 44824 5108 44876 5160
rect 34704 5015 34756 5024
rect 34704 4981 34713 5015
rect 34713 4981 34747 5015
rect 34747 4981 34756 5015
rect 34704 4972 34756 4981
rect 36176 5015 36228 5024
rect 36176 4981 36185 5015
rect 36185 4981 36219 5015
rect 36219 4981 36228 5015
rect 36176 4972 36228 4981
rect 42984 4972 43036 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1860 4768 1912 4820
rect 10048 4768 10100 4820
rect 13084 4700 13136 4752
rect 13176 4743 13228 4752
rect 13176 4709 13185 4743
rect 13185 4709 13219 4743
rect 13219 4709 13228 4743
rect 13176 4700 13228 4709
rect 3240 4632 3292 4684
rect 8484 4632 8536 4684
rect 10600 4632 10652 4684
rect 11980 4632 12032 4684
rect 13636 4632 13688 4684
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 8300 4564 8352 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9680 4564 9732 4616
rect 13544 4564 13596 4616
rect 2688 4496 2740 4548
rect 11980 4496 12032 4548
rect 7656 4428 7708 4480
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 13544 4428 13596 4437
rect 16120 4496 16172 4548
rect 16856 4539 16908 4548
rect 16856 4505 16865 4539
rect 16865 4505 16899 4539
rect 16899 4505 16908 4539
rect 16856 4496 16908 4505
rect 20352 4768 20404 4820
rect 21272 4768 21324 4820
rect 23204 4768 23256 4820
rect 23572 4811 23624 4820
rect 23572 4777 23581 4811
rect 23581 4777 23615 4811
rect 23615 4777 23624 4811
rect 23572 4768 23624 4777
rect 18696 4700 18748 4752
rect 17960 4564 18012 4616
rect 19156 4564 19208 4616
rect 20812 4632 20864 4684
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 22100 4632 22152 4684
rect 23848 4768 23900 4820
rect 34704 4768 34756 4820
rect 36176 4768 36228 4820
rect 37924 4768 37976 4820
rect 38016 4811 38068 4820
rect 38016 4777 38025 4811
rect 38025 4777 38059 4811
rect 38059 4777 38068 4811
rect 38016 4768 38068 4777
rect 23756 4632 23808 4684
rect 21548 4564 21600 4616
rect 23112 4564 23164 4616
rect 39580 4768 39632 4820
rect 40868 4768 40920 4820
rect 41052 4768 41104 4820
rect 42156 4768 42208 4820
rect 34520 4632 34572 4684
rect 35348 4632 35400 4684
rect 16580 4428 16632 4480
rect 18788 4428 18840 4480
rect 19984 4428 20036 4480
rect 24860 4564 24912 4616
rect 28540 4564 28592 4616
rect 29552 4607 29604 4616
rect 29552 4573 29561 4607
rect 29561 4573 29595 4607
rect 29595 4573 29604 4607
rect 29552 4564 29604 4573
rect 31300 4607 31352 4616
rect 31300 4573 31309 4607
rect 31309 4573 31343 4607
rect 31343 4573 31352 4607
rect 31300 4564 31352 4573
rect 32772 4607 32824 4616
rect 32772 4573 32781 4607
rect 32781 4573 32815 4607
rect 32815 4573 32824 4607
rect 32772 4564 32824 4573
rect 38752 4700 38804 4752
rect 38844 4632 38896 4684
rect 39580 4632 39632 4684
rect 33784 4496 33836 4548
rect 25412 4428 25464 4480
rect 33048 4428 33100 4480
rect 34612 4428 34664 4480
rect 36728 4496 36780 4548
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 40040 4607 40092 4616
rect 40040 4573 40049 4607
rect 40049 4573 40083 4607
rect 40083 4573 40092 4607
rect 40040 4564 40092 4573
rect 38016 4496 38068 4548
rect 36544 4428 36596 4480
rect 37188 4471 37240 4480
rect 37188 4437 37197 4471
rect 37197 4437 37231 4471
rect 37231 4437 37240 4471
rect 37188 4428 37240 4437
rect 38200 4428 38252 4480
rect 39304 4428 39356 4480
rect 41052 4564 41104 4616
rect 41328 4607 41380 4616
rect 41328 4573 41337 4607
rect 41337 4573 41371 4607
rect 41371 4573 41380 4607
rect 41328 4564 41380 4573
rect 41420 4607 41472 4616
rect 41420 4573 41429 4607
rect 41429 4573 41463 4607
rect 41463 4573 41472 4607
rect 41420 4564 41472 4573
rect 40776 4496 40828 4548
rect 40684 4428 40736 4480
rect 41512 4496 41564 4548
rect 42248 4564 42300 4616
rect 41696 4428 41748 4480
rect 41972 4496 42024 4548
rect 42892 4496 42944 4548
rect 43168 4496 43220 4548
rect 42800 4471 42852 4480
rect 42800 4437 42809 4471
rect 42809 4437 42843 4471
rect 42843 4437 42852 4471
rect 42800 4428 42852 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3056 4224 3108 4276
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 19156 4224 19208 4276
rect 20168 4224 20220 4276
rect 7288 4156 7340 4208
rect 3240 4088 3292 4140
rect 6184 4088 6236 4140
rect 7656 4088 7708 4140
rect 9680 4156 9732 4208
rect 10968 4156 11020 4208
rect 11980 4156 12032 4208
rect 4620 4020 4672 4072
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 14096 4088 14148 4140
rect 15568 4156 15620 4208
rect 18788 4156 18840 4208
rect 8024 4020 8076 4072
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 12532 4020 12584 4072
rect 13636 4020 13688 4072
rect 7748 3952 7800 4004
rect 8944 3952 8996 4004
rect 16304 4088 16356 4140
rect 16580 4088 16632 4140
rect 19616 4088 19668 4140
rect 19984 4088 20036 4140
rect 29000 4224 29052 4276
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 26056 4088 26108 4140
rect 27068 4088 27120 4140
rect 14280 4063 14332 4072
rect 14280 4029 14289 4063
rect 14289 4029 14323 4063
rect 14323 4029 14332 4063
rect 14280 4020 14332 4029
rect 6000 3884 6052 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 14832 3952 14884 4004
rect 15200 3995 15252 4004
rect 15200 3961 15209 3995
rect 15209 3961 15243 3995
rect 15243 3961 15252 3995
rect 15200 3952 15252 3961
rect 18052 4020 18104 4072
rect 20536 4020 20588 4072
rect 28540 4063 28592 4072
rect 28540 4029 28549 4063
rect 28549 4029 28583 4063
rect 28583 4029 28592 4063
rect 28540 4020 28592 4029
rect 28816 4063 28868 4072
rect 28816 4029 28825 4063
rect 28825 4029 28859 4063
rect 28859 4029 28868 4063
rect 28816 4020 28868 4029
rect 31392 4020 31444 4072
rect 19524 3952 19576 4004
rect 32220 4088 32272 4140
rect 33048 4088 33100 4140
rect 34244 4224 34296 4276
rect 34704 4224 34756 4276
rect 35440 4224 35492 4276
rect 34152 4131 34204 4140
rect 34152 4097 34161 4131
rect 34161 4097 34195 4131
rect 34195 4097 34204 4131
rect 34152 4088 34204 4097
rect 34244 4088 34296 4140
rect 34612 4131 34664 4140
rect 34612 4097 34621 4131
rect 34621 4097 34655 4131
rect 34655 4097 34664 4131
rect 34612 4088 34664 4097
rect 33968 4020 34020 4072
rect 34060 3952 34112 4004
rect 35900 4088 35952 4140
rect 36636 4224 36688 4276
rect 37832 4224 37884 4276
rect 38752 4224 38804 4276
rect 40040 4224 40092 4276
rect 41420 4224 41472 4276
rect 36176 4156 36228 4208
rect 37188 4156 37240 4208
rect 35716 4020 35768 4072
rect 36452 4020 36504 4072
rect 37096 4131 37148 4140
rect 37096 4097 37105 4131
rect 37105 4097 37139 4131
rect 37139 4097 37148 4131
rect 37096 4088 37148 4097
rect 38200 4131 38252 4140
rect 38200 4097 38209 4131
rect 38209 4097 38243 4131
rect 38243 4097 38252 4131
rect 38200 4088 38252 4097
rect 37280 4020 37332 4072
rect 38016 4063 38068 4072
rect 38016 4029 38025 4063
rect 38025 4029 38059 4063
rect 38059 4029 38068 4063
rect 38016 4020 38068 4029
rect 36084 3952 36136 4004
rect 17408 3884 17460 3936
rect 18696 3884 18748 3936
rect 25780 3927 25832 3936
rect 25780 3893 25789 3927
rect 25789 3893 25823 3927
rect 25823 3893 25832 3927
rect 25780 3884 25832 3893
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 27160 3884 27212 3893
rect 27344 3884 27396 3936
rect 31852 3884 31904 3936
rect 33232 3927 33284 3936
rect 33232 3893 33241 3927
rect 33241 3893 33275 3927
rect 33275 3893 33284 3927
rect 33232 3884 33284 3893
rect 33968 3927 34020 3936
rect 33968 3893 33977 3927
rect 33977 3893 34011 3927
rect 34011 3893 34020 3927
rect 33968 3884 34020 3893
rect 34152 3884 34204 3936
rect 34428 3927 34480 3936
rect 34428 3893 34437 3927
rect 34437 3893 34471 3927
rect 34471 3893 34480 3927
rect 34428 3884 34480 3893
rect 34520 3884 34572 3936
rect 35532 3884 35584 3936
rect 36728 3952 36780 4004
rect 36912 3995 36964 4004
rect 36912 3961 36921 3995
rect 36921 3961 36955 3995
rect 36955 3961 36964 3995
rect 36912 3952 36964 3961
rect 36544 3927 36596 3936
rect 36544 3893 36553 3927
rect 36553 3893 36587 3927
rect 36587 3893 36596 3927
rect 36544 3884 36596 3893
rect 43444 4224 43496 4276
rect 40500 4131 40552 4140
rect 40500 4097 40509 4131
rect 40509 4097 40543 4131
rect 40543 4097 40552 4131
rect 40500 4088 40552 4097
rect 40684 4131 40736 4140
rect 40684 4097 40693 4131
rect 40693 4097 40727 4131
rect 40727 4097 40736 4131
rect 40684 4088 40736 4097
rect 40868 4088 40920 4140
rect 40960 4131 41012 4140
rect 40960 4097 40969 4131
rect 40969 4097 41003 4131
rect 41003 4097 41012 4131
rect 40960 4088 41012 4097
rect 39120 4020 39172 4072
rect 41328 4088 41380 4140
rect 42340 4088 42392 4140
rect 42064 4020 42116 4072
rect 38384 3927 38436 3936
rect 38384 3893 38393 3927
rect 38393 3893 38427 3927
rect 38427 3893 38436 3927
rect 38384 3884 38436 3893
rect 41236 3927 41288 3936
rect 41236 3893 41245 3927
rect 41245 3893 41279 3927
rect 41279 3893 41288 3927
rect 41236 3884 41288 3893
rect 42800 4020 42852 4072
rect 43168 4020 43220 4072
rect 43076 3884 43128 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3240 3544 3292 3596
rect 7748 3680 7800 3732
rect 8208 3680 8260 3732
rect 9312 3680 9364 3732
rect 9588 3723 9640 3732
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 12992 3680 13044 3732
rect 16304 3680 16356 3732
rect 5540 3544 5592 3596
rect 5448 3476 5500 3528
rect 7288 3408 7340 3460
rect 7656 3408 7708 3460
rect 8024 3408 8076 3460
rect 9588 3544 9640 3596
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 11520 3544 11572 3596
rect 12900 3587 12952 3596
rect 12900 3553 12909 3587
rect 12909 3553 12943 3587
rect 12943 3553 12952 3587
rect 12900 3544 12952 3553
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 14280 3544 14332 3596
rect 19616 3680 19668 3732
rect 24492 3680 24544 3732
rect 25780 3680 25832 3732
rect 9772 3476 9824 3528
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 6920 3340 6972 3392
rect 11980 3408 12032 3460
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 16856 3544 16908 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 18696 3544 18748 3596
rect 25688 3544 25740 3596
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 28540 3680 28592 3732
rect 26516 3544 26568 3553
rect 28816 3680 28868 3732
rect 29828 3723 29880 3732
rect 29828 3689 29837 3723
rect 29837 3689 29871 3723
rect 29871 3689 29880 3723
rect 29828 3680 29880 3689
rect 32680 3723 32732 3732
rect 32680 3689 32710 3723
rect 32710 3689 32732 3723
rect 32680 3680 32732 3689
rect 34520 3723 34572 3732
rect 34520 3689 34529 3723
rect 34529 3689 34563 3723
rect 34563 3689 34572 3723
rect 34520 3680 34572 3689
rect 34612 3680 34664 3732
rect 35624 3680 35676 3732
rect 37096 3680 37148 3732
rect 38384 3680 38436 3732
rect 40500 3680 40552 3732
rect 33968 3612 34020 3664
rect 37372 3612 37424 3664
rect 30472 3587 30524 3596
rect 30472 3553 30481 3587
rect 30481 3553 30515 3587
rect 30515 3553 30524 3587
rect 30472 3544 30524 3553
rect 32772 3544 32824 3596
rect 33232 3544 33284 3596
rect 17592 3476 17644 3528
rect 18144 3476 18196 3528
rect 23756 3476 23808 3528
rect 25964 3476 26016 3528
rect 12716 3340 12768 3392
rect 16120 3340 16172 3392
rect 17960 3340 18012 3392
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 29000 3476 29052 3528
rect 30564 3476 30616 3528
rect 30840 3519 30892 3528
rect 30840 3485 30849 3519
rect 30849 3485 30883 3519
rect 30883 3485 30892 3519
rect 30840 3476 30892 3485
rect 34704 3544 34756 3596
rect 35440 3587 35492 3596
rect 35440 3553 35449 3587
rect 35449 3553 35483 3587
rect 35483 3553 35492 3587
rect 35440 3544 35492 3553
rect 35900 3587 35952 3596
rect 35900 3553 35909 3587
rect 35909 3553 35943 3587
rect 35943 3553 35952 3587
rect 35900 3544 35952 3553
rect 36912 3544 36964 3596
rect 37188 3587 37240 3596
rect 37188 3553 37197 3587
rect 37197 3553 37231 3587
rect 37231 3553 37240 3587
rect 37188 3544 37240 3553
rect 31852 3408 31904 3460
rect 34428 3408 34480 3460
rect 37556 3476 37608 3528
rect 38016 3476 38068 3528
rect 39580 3587 39632 3596
rect 39580 3553 39589 3587
rect 39589 3553 39623 3587
rect 39623 3553 39632 3587
rect 39580 3544 39632 3553
rect 39304 3519 39356 3528
rect 39304 3485 39313 3519
rect 39313 3485 39347 3519
rect 39347 3485 39356 3519
rect 39304 3476 39356 3485
rect 34152 3383 34204 3392
rect 34152 3349 34161 3383
rect 34161 3349 34195 3383
rect 34195 3349 34204 3383
rect 34152 3340 34204 3349
rect 34612 3340 34664 3392
rect 38568 3383 38620 3392
rect 38568 3349 38577 3383
rect 38577 3349 38611 3383
rect 38611 3349 38620 3383
rect 38568 3340 38620 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4528 3136 4580 3188
rect 5540 3136 5592 3188
rect 6000 3136 6052 3188
rect 6184 3136 6236 3188
rect 9496 3068 9548 3120
rect 12900 3136 12952 3188
rect 13728 3136 13780 3188
rect 14556 3136 14608 3188
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 9588 3000 9640 3052
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 12072 2932 12124 2984
rect 12716 3000 12768 3052
rect 13636 3000 13688 3052
rect 13544 2932 13596 2984
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 18144 3136 18196 3188
rect 17408 3111 17460 3120
rect 17408 3077 17417 3111
rect 17417 3077 17451 3111
rect 17451 3077 17460 3111
rect 17408 3068 17460 3077
rect 16120 2932 16172 2984
rect 17500 2932 17552 2984
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 25596 3136 25648 3188
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 27068 3136 27120 3188
rect 27344 3136 27396 3188
rect 29368 3136 29420 3188
rect 30472 3136 30524 3188
rect 30564 3136 30616 3188
rect 30840 3136 30892 3188
rect 29000 3068 29052 3120
rect 29736 3068 29788 3120
rect 34704 3179 34756 3188
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 35440 3136 35492 3188
rect 26516 3000 26568 3052
rect 10508 2907 10560 2916
rect 10508 2873 10517 2907
rect 10517 2873 10551 2907
rect 10551 2873 10560 2907
rect 10508 2864 10560 2873
rect 12808 2864 12860 2916
rect 18052 2864 18104 2916
rect 25872 2907 25924 2916
rect 25872 2873 25881 2907
rect 25881 2873 25915 2907
rect 25915 2873 25924 2907
rect 25872 2864 25924 2873
rect 26608 2907 26660 2916
rect 26608 2873 26617 2907
rect 26617 2873 26651 2907
rect 26651 2873 26660 2907
rect 26608 2864 26660 2873
rect 29000 2932 29052 2984
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 33784 3068 33836 3120
rect 34520 3068 34572 3120
rect 34612 3068 34664 3120
rect 30840 2907 30892 2916
rect 30840 2873 30849 2907
rect 30849 2873 30883 2907
rect 30883 2873 30892 2907
rect 30840 2864 30892 2873
rect 32220 2796 32272 2848
rect 32864 3000 32916 3052
rect 35532 3068 35584 3120
rect 37188 3136 37240 3188
rect 37556 3179 37608 3188
rect 37556 3145 37565 3179
rect 37565 3145 37599 3179
rect 37599 3145 37608 3179
rect 37556 3136 37608 3145
rect 39212 3136 39264 3188
rect 41236 3136 41288 3188
rect 42064 3179 42116 3188
rect 42064 3145 42073 3179
rect 42073 3145 42107 3179
rect 42107 3145 42116 3179
rect 42064 3136 42116 3145
rect 35348 3043 35400 3052
rect 35348 3009 35357 3043
rect 35357 3009 35391 3043
rect 35391 3009 35400 3043
rect 35348 3000 35400 3009
rect 36728 3000 36780 3052
rect 42340 3068 42392 3120
rect 34244 2864 34296 2916
rect 38568 2932 38620 2984
rect 34428 2796 34480 2848
rect 35716 2796 35768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 10508 2592 10560 2644
rect 12072 2592 12124 2644
rect 25872 2592 25924 2644
rect 26608 2592 26660 2644
rect 30288 2592 30340 2644
rect 32680 2635 32732 2644
rect 32680 2601 32689 2635
rect 32689 2601 32723 2635
rect 32723 2601 32732 2635
rect 32680 2592 32732 2601
rect 43904 2635 43956 2644
rect 43904 2601 43913 2635
rect 43913 2601 43947 2635
rect 43947 2601 43956 2635
rect 43904 2592 43956 2601
rect 18052 2524 18104 2576
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 8300 2456 8352 2508
rect 29184 2456 29236 2508
rect 32220 2499 32272 2508
rect 32220 2465 32229 2499
rect 32229 2465 32263 2499
rect 32263 2465 32272 2499
rect 32220 2456 32272 2465
rect 20 2388 72 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 26516 2431 26568 2440
rect 26516 2397 26525 2431
rect 26525 2397 26559 2431
rect 26559 2397 26568 2431
rect 26516 2388 26568 2397
rect 33232 2388 33284 2440
rect 43812 2388 43864 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 6458 47681 6514 48481
rect 14830 47681 14886 48481
rect 23846 47681 23902 48481
rect 32862 47818 32918 48481
rect 32862 47790 33088 47818
rect 32862 47681 32918 47790
rect 938 46336 994 46345
rect 938 46271 994 46280
rect 952 46034 980 46271
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 940 46028 992 46034
rect 940 45970 992 45976
rect 6472 45966 6500 47681
rect 14844 46170 14872 47681
rect 14832 46164 14884 46170
rect 14832 46106 14884 46112
rect 21824 46028 21876 46034
rect 21824 45970 21876 45976
rect 1676 45960 1728 45966
rect 1676 45902 1728 45908
rect 6460 45960 6512 45966
rect 6460 45902 6512 45908
rect 9864 45960 9916 45966
rect 9864 45902 9916 45908
rect 14832 45960 14884 45966
rect 14832 45902 14884 45908
rect 1688 45554 1716 45902
rect 7472 45824 7524 45830
rect 7472 45766 7524 45772
rect 8852 45824 8904 45830
rect 8852 45766 8904 45772
rect 1688 45526 1808 45554
rect 1780 41414 1808 45526
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 7484 43382 7512 45766
rect 8864 44878 8892 45766
rect 9036 45280 9088 45286
rect 9036 45222 9088 45228
rect 9048 45082 9076 45222
rect 9036 45076 9088 45082
rect 9036 45018 9088 45024
rect 8944 44940 8996 44946
rect 8944 44882 8996 44888
rect 8852 44872 8904 44878
rect 8852 44814 8904 44820
rect 8576 44736 8628 44742
rect 8576 44678 8628 44684
rect 8588 44402 8616 44678
rect 8956 44538 8984 44882
rect 9876 44538 9904 45902
rect 14004 45824 14056 45830
rect 14004 45766 14056 45772
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 13728 45552 13780 45558
rect 13728 45494 13780 45500
rect 9956 45416 10008 45422
rect 9956 45358 10008 45364
rect 9968 44538 9996 45358
rect 10060 44742 10088 45494
rect 10140 45484 10192 45490
rect 10140 45426 10192 45432
rect 11704 45484 11756 45490
rect 11704 45426 11756 45432
rect 13544 45484 13596 45490
rect 13544 45426 13596 45432
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 8944 44532 8996 44538
rect 8944 44474 8996 44480
rect 9864 44532 9916 44538
rect 9864 44474 9916 44480
rect 9956 44532 10008 44538
rect 9956 44474 10008 44480
rect 8576 44396 8628 44402
rect 8576 44338 8628 44344
rect 9312 44328 9364 44334
rect 9312 44270 9364 44276
rect 8208 44192 8260 44198
rect 8208 44134 8260 44140
rect 8220 43994 8248 44134
rect 8208 43988 8260 43994
rect 8208 43930 8260 43936
rect 8024 43648 8076 43654
rect 8024 43590 8076 43596
rect 8036 43450 8064 43590
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 8024 43444 8076 43450
rect 8024 43386 8076 43392
rect 7472 43376 7524 43382
rect 7472 43318 7524 43324
rect 6920 43240 6972 43246
rect 6920 43182 6972 43188
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 3884 42696 3936 42702
rect 3884 42638 3936 42644
rect 4896 42696 4948 42702
rect 4896 42638 4948 42644
rect 5356 42696 5408 42702
rect 5356 42638 5408 42644
rect 3896 42362 3924 42638
rect 4160 42560 4212 42566
rect 4160 42502 4212 42508
rect 4620 42560 4672 42566
rect 4620 42502 4672 42508
rect 3884 42356 3936 42362
rect 3884 42298 3936 42304
rect 3332 42152 3384 42158
rect 3332 42094 3384 42100
rect 3344 41682 3372 42094
rect 3896 41818 3924 42298
rect 4172 42106 4200 42502
rect 4080 42078 4200 42106
rect 3884 41812 3936 41818
rect 4080 41800 4108 42078
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4632 41818 4660 42502
rect 4712 42084 4764 42090
rect 4712 42026 4764 42032
rect 4620 41812 4672 41818
rect 4080 41772 4292 41800
rect 3884 41754 3936 41760
rect 2780 41676 2832 41682
rect 2780 41618 2832 41624
rect 3332 41676 3384 41682
rect 3332 41618 3384 41624
rect 1860 41608 1912 41614
rect 1860 41550 1912 41556
rect 1688 41386 1808 41414
rect 1492 38344 1544 38350
rect 1492 38286 1544 38292
rect 1504 37806 1532 38286
rect 1492 37800 1544 37806
rect 1492 37742 1544 37748
rect 940 37256 992 37262
rect 940 37198 992 37204
rect 952 36825 980 37198
rect 938 36816 994 36825
rect 1504 36786 1532 37742
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 938 36751 994 36760
rect 1492 36780 1544 36786
rect 1492 36722 1544 36728
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1504 31278 1532 32302
rect 1492 31272 1544 31278
rect 1492 31214 1544 31220
rect 1504 30802 1532 31214
rect 1492 30796 1544 30802
rect 1492 30738 1544 30744
rect 940 28076 992 28082
rect 940 28018 992 28024
rect 952 27985 980 28018
rect 938 27976 994 27985
rect 938 27911 994 27920
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1596 15978 1624 37062
rect 1688 18970 1716 41386
rect 1872 40594 1900 41550
rect 2792 41274 2820 41618
rect 2780 41268 2832 41274
rect 2780 41210 2832 41216
rect 1860 40588 1912 40594
rect 1860 40530 1912 40536
rect 3344 40458 3372 41618
rect 4264 41546 4292 41772
rect 4620 41754 4672 41760
rect 4344 41744 4396 41750
rect 4344 41686 4396 41692
rect 4252 41540 4304 41546
rect 4252 41482 4304 41488
rect 4160 41472 4212 41478
rect 4160 41414 4212 41420
rect 4172 41274 4200 41414
rect 4160 41268 4212 41274
rect 4160 41210 4212 41216
rect 4160 41132 4212 41138
rect 4160 41074 4212 41080
rect 3792 41064 3844 41070
rect 4172 41018 4200 41074
rect 3792 41006 3844 41012
rect 3516 40928 3568 40934
rect 3516 40870 3568 40876
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 3332 40452 3384 40458
rect 3332 40394 3384 40400
rect 1872 40186 1900 40394
rect 1860 40180 1912 40186
rect 1860 40122 1912 40128
rect 3528 39982 3556 40870
rect 3608 40588 3660 40594
rect 3608 40530 3660 40536
rect 3620 40050 3648 40530
rect 3608 40044 3660 40050
rect 3608 39986 3660 39992
rect 3516 39976 3568 39982
rect 3516 39918 3568 39924
rect 2596 39432 2648 39438
rect 2596 39374 2648 39380
rect 2504 39296 2556 39302
rect 2504 39238 2556 39244
rect 2136 38276 2188 38282
rect 2136 38218 2188 38224
rect 2148 38010 2176 38218
rect 2516 38010 2544 39238
rect 2608 39098 2636 39374
rect 3148 39296 3200 39302
rect 3148 39238 3200 39244
rect 2596 39092 2648 39098
rect 2596 39034 2648 39040
rect 2872 38956 2924 38962
rect 2872 38898 2924 38904
rect 2136 38004 2188 38010
rect 2136 37946 2188 37952
rect 2504 38004 2556 38010
rect 2504 37946 2556 37952
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2792 37466 2820 37810
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2884 37330 2912 38898
rect 3160 38894 3188 39238
rect 3148 38888 3200 38894
rect 3148 38830 3200 38836
rect 3620 37874 3648 39986
rect 3608 37868 3660 37874
rect 3608 37810 3660 37816
rect 2872 37324 2924 37330
rect 2872 37266 2924 37272
rect 1952 37120 2004 37126
rect 1952 37062 2004 37068
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 1964 36922 1992 37062
rect 2792 36922 2820 37062
rect 1952 36916 2004 36922
rect 1952 36858 2004 36864
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 3804 36802 3832 41006
rect 4080 40990 4200 41018
rect 4080 40610 4108 40990
rect 4264 40934 4292 41482
rect 4356 41414 4384 41686
rect 4356 41386 4660 41414
rect 4356 41138 4384 41386
rect 4528 41268 4580 41274
rect 4528 41210 4580 41216
rect 4540 41138 4568 41210
rect 4344 41132 4396 41138
rect 4344 41074 4396 41080
rect 4528 41132 4580 41138
rect 4528 41074 4580 41080
rect 4252 40928 4304 40934
rect 4252 40870 4304 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4632 40730 4660 41386
rect 4724 41138 4752 42026
rect 4908 41818 4936 42638
rect 5368 42294 5396 42638
rect 5448 42560 5500 42566
rect 5448 42502 5500 42508
rect 6460 42560 6512 42566
rect 6460 42502 6512 42508
rect 5460 42362 5488 42502
rect 6472 42362 6500 42502
rect 6932 42362 6960 43182
rect 7472 43104 7524 43110
rect 7472 43046 7524 43052
rect 7484 42906 7512 43046
rect 7760 42922 7788 43386
rect 7932 43376 7984 43382
rect 7932 43318 7984 43324
rect 7472 42900 7524 42906
rect 7472 42842 7524 42848
rect 7668 42894 7788 42922
rect 7472 42560 7524 42566
rect 7472 42502 7524 42508
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 6460 42356 6512 42362
rect 6460 42298 6512 42304
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 5356 42288 5408 42294
rect 5356 42230 5408 42236
rect 5368 42158 5396 42230
rect 6368 42220 6420 42226
rect 6368 42162 6420 42168
rect 5356 42152 5408 42158
rect 5356 42094 5408 42100
rect 6092 42152 6144 42158
rect 6092 42094 6144 42100
rect 5356 42016 5408 42022
rect 5356 41958 5408 41964
rect 5448 42016 5500 42022
rect 5448 41958 5500 41964
rect 5368 41818 5396 41958
rect 4896 41812 4948 41818
rect 4896 41754 4948 41760
rect 5356 41812 5408 41818
rect 5460 41800 5488 41958
rect 5460 41772 5580 41800
rect 5356 41754 5408 41760
rect 4804 41744 4856 41750
rect 4804 41686 4856 41692
rect 4816 41138 4844 41686
rect 5448 41676 5500 41682
rect 5448 41618 5500 41624
rect 4988 41608 5040 41614
rect 4988 41550 5040 41556
rect 5000 41274 5028 41550
rect 5264 41540 5316 41546
rect 5264 41482 5316 41488
rect 4988 41268 5040 41274
rect 4988 41210 5040 41216
rect 5000 41138 5028 41210
rect 5172 41200 5224 41206
rect 5172 41142 5224 41148
rect 4712 41132 4764 41138
rect 4712 41074 4764 41080
rect 4804 41132 4856 41138
rect 4804 41074 4856 41080
rect 4988 41132 5040 41138
rect 4988 41074 5040 41080
rect 4620 40724 4672 40730
rect 4620 40666 4672 40672
rect 4080 40594 4200 40610
rect 4816 40594 4844 41074
rect 4080 40588 4212 40594
rect 4080 40582 4160 40588
rect 4160 40530 4212 40536
rect 4804 40588 4856 40594
rect 4804 40530 4856 40536
rect 4620 40520 4672 40526
rect 4620 40462 4672 40468
rect 4344 40452 4396 40458
rect 4344 40394 4396 40400
rect 4068 40384 4120 40390
rect 4068 40326 4120 40332
rect 4080 40186 4108 40326
rect 4068 40180 4120 40186
rect 4068 40122 4120 40128
rect 4356 40118 4384 40394
rect 4344 40112 4396 40118
rect 4344 40054 4396 40060
rect 3976 39976 4028 39982
rect 3976 39918 4028 39924
rect 3988 39642 4016 39918
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 3976 39636 4028 39642
rect 3976 39578 4028 39584
rect 4528 39568 4580 39574
rect 4528 39510 4580 39516
rect 4540 38962 4568 39510
rect 4632 39098 4660 40462
rect 4816 39574 4844 40530
rect 4804 39568 4856 39574
rect 4804 39510 4856 39516
rect 4620 39092 4672 39098
rect 4620 39034 4672 39040
rect 4528 38956 4580 38962
rect 4528 38898 4580 38904
rect 5000 38894 5028 41074
rect 5080 40520 5132 40526
rect 5080 40462 5132 40468
rect 3976 38888 4028 38894
rect 3976 38830 4028 38836
rect 4988 38888 5040 38894
rect 4988 38830 5040 38836
rect 3988 38554 4016 38830
rect 4712 38820 4764 38826
rect 4712 38762 4764 38768
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 3976 38548 4028 38554
rect 3976 38490 4028 38496
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 38150
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 3712 36774 3832 36802
rect 3332 35692 3384 35698
rect 3332 35634 3384 35640
rect 2964 35488 3016 35494
rect 2964 35430 3016 35436
rect 2976 35086 3004 35430
rect 3344 35290 3372 35634
rect 3332 35284 3384 35290
rect 3332 35226 3384 35232
rect 2964 35080 3016 35086
rect 2964 35022 3016 35028
rect 2136 35012 2188 35018
rect 2136 34954 2188 34960
rect 2148 34746 2176 34954
rect 3056 34944 3108 34950
rect 3056 34886 3108 34892
rect 2136 34740 2188 34746
rect 2136 34682 2188 34688
rect 2872 34468 2924 34474
rect 2872 34410 2924 34416
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 2424 32910 2452 33798
rect 2504 33312 2556 33318
rect 2504 33254 2556 33260
rect 2596 33312 2648 33318
rect 2596 33254 2648 33260
rect 2516 32978 2544 33254
rect 2504 32972 2556 32978
rect 2504 32914 2556 32920
rect 2412 32904 2464 32910
rect 2412 32846 2464 32852
rect 1768 32768 1820 32774
rect 1768 32710 1820 32716
rect 1780 32502 1808 32710
rect 1768 32496 1820 32502
rect 1768 32438 1820 32444
rect 2424 31890 2452 32846
rect 2412 31884 2464 31890
rect 2412 31826 2464 31832
rect 2608 31754 2636 33254
rect 2884 32978 2912 34410
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 3068 32434 3096 34886
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3252 32570 3280 33934
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 3528 33114 3556 33458
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3712 32910 3740 36774
rect 3792 36712 3844 36718
rect 3792 36654 3844 36660
rect 3804 36378 3832 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3792 36372 3844 36378
rect 3792 36314 3844 36320
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 3792 34604 3844 34610
rect 3792 34546 3844 34552
rect 3700 32904 3752 32910
rect 3700 32846 3752 32852
rect 3804 32570 3832 34546
rect 3884 33924 3936 33930
rect 3884 33866 3936 33872
rect 3896 33658 3924 33866
rect 3884 33652 3936 33658
rect 3884 33594 3936 33600
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3792 32564 3844 32570
rect 3792 32506 3844 32512
rect 3056 32428 3108 32434
rect 3056 32370 3108 32376
rect 2516 31726 2636 31754
rect 2412 31680 2464 31686
rect 2412 31622 2464 31628
rect 2424 31482 2452 31622
rect 2412 31476 2464 31482
rect 2412 31418 2464 31424
rect 2516 31278 2544 31726
rect 3240 31680 3292 31686
rect 3240 31622 3292 31628
rect 2504 31272 2556 31278
rect 2504 31214 2556 31220
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 1860 31136 1912 31142
rect 1860 31078 1912 31084
rect 1872 30802 1900 31078
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 2516 30394 2544 31214
rect 2792 30938 2820 31214
rect 2780 30932 2832 30938
rect 2780 30874 2832 30880
rect 3252 30870 3280 31622
rect 3424 31272 3476 31278
rect 3424 31214 3476 31220
rect 3240 30864 3292 30870
rect 3240 30806 3292 30812
rect 3436 30734 3464 31214
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3804 30666 3832 32506
rect 4080 31482 4108 35974
rect 4724 35834 4752 38762
rect 5092 38554 5120 40462
rect 5080 38548 5132 38554
rect 5080 38490 5132 38496
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4908 37466 4936 37810
rect 4896 37460 4948 37466
rect 4896 37402 4948 37408
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 4712 35828 4764 35834
rect 4712 35770 4764 35776
rect 4620 35488 4672 35494
rect 4620 35430 4672 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 35430
rect 4816 35290 4844 37266
rect 4988 37120 5040 37126
rect 4988 37062 5040 37068
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 4804 35284 4856 35290
rect 4804 35226 4856 35232
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 4264 34746 4292 35022
rect 4252 34740 4304 34746
rect 4252 34682 4304 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4160 33924 4212 33930
rect 4160 33866 4212 33872
rect 4172 33522 4200 33866
rect 4160 33516 4212 33522
rect 4160 33458 4212 33464
rect 4632 33454 4660 35090
rect 4804 34400 4856 34406
rect 4804 34342 4856 34348
rect 4816 33658 4844 34342
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33390
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30682 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30938 4660 31962
rect 4896 31408 4948 31414
rect 4896 31350 4948 31356
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 3792 30660 3844 30666
rect 4080 30654 4200 30682
rect 3792 30602 3844 30608
rect 4172 30598 4200 30654
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4816 30394 4844 30534
rect 2504 30388 2556 30394
rect 2504 30330 2556 30336
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4908 30326 4936 31350
rect 4896 30320 4948 30326
rect 4896 30262 4948 30268
rect 4908 30054 4936 30262
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4804 28144 4856 28150
rect 4908 28132 4936 29990
rect 5000 29646 5028 37062
rect 5080 36032 5132 36038
rect 5080 35974 5132 35980
rect 5092 35018 5120 35974
rect 5080 35012 5132 35018
rect 5080 34954 5132 34960
rect 5184 34610 5212 41142
rect 5276 38758 5304 41482
rect 5460 40934 5488 41618
rect 5552 41614 5580 41772
rect 5540 41608 5592 41614
rect 5540 41550 5592 41556
rect 6104 41414 6132 42094
rect 6380 41818 6408 42162
rect 6368 41812 6420 41818
rect 6368 41754 6420 41760
rect 6472 41682 6500 42298
rect 7484 42226 7512 42502
rect 6736 42220 6788 42226
rect 6736 42162 6788 42168
rect 7472 42220 7524 42226
rect 7472 42162 7524 42168
rect 6460 41676 6512 41682
rect 6460 41618 6512 41624
rect 6104 41386 6224 41414
rect 6092 41064 6144 41070
rect 6092 41006 6144 41012
rect 5448 40928 5500 40934
rect 5448 40870 5500 40876
rect 6104 39846 6132 41006
rect 6196 40594 6224 41386
rect 6748 40730 6776 42162
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 6736 40724 6788 40730
rect 6736 40666 6788 40672
rect 6184 40588 6236 40594
rect 6184 40530 6236 40536
rect 6196 40050 6224 40530
rect 6184 40044 6236 40050
rect 6184 39986 6236 39992
rect 6092 39840 6144 39846
rect 6092 39782 6144 39788
rect 5908 39296 5960 39302
rect 5908 39238 5960 39244
rect 5920 38826 5948 39238
rect 6104 39030 6132 39782
rect 6196 39642 6224 39986
rect 6644 39976 6696 39982
rect 6644 39918 6696 39924
rect 6656 39642 6684 39918
rect 6184 39636 6236 39642
rect 6184 39578 6236 39584
rect 6644 39636 6696 39642
rect 6644 39578 6696 39584
rect 6368 39500 6420 39506
rect 6368 39442 6420 39448
rect 6092 39024 6144 39030
rect 6092 38966 6144 38972
rect 5908 38820 5960 38826
rect 5908 38762 5960 38768
rect 5264 38752 5316 38758
rect 5264 38694 5316 38700
rect 5276 38418 5304 38694
rect 5264 38412 5316 38418
rect 5264 38354 5316 38360
rect 5276 38010 5304 38354
rect 5264 38004 5316 38010
rect 5264 37946 5316 37952
rect 5448 37868 5500 37874
rect 5448 37810 5500 37816
rect 5460 37330 5488 37810
rect 5920 37346 5948 38762
rect 6000 37664 6052 37670
rect 6000 37606 6052 37612
rect 6184 37664 6236 37670
rect 6184 37606 6236 37612
rect 5736 37330 5948 37346
rect 6012 37330 6040 37606
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5736 37324 5960 37330
rect 5736 37318 5908 37324
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5356 36168 5408 36174
rect 5356 36110 5408 36116
rect 5368 35834 5396 36110
rect 5552 36038 5580 36790
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5356 35828 5408 35834
rect 5356 35770 5408 35776
rect 5552 35018 5580 35974
rect 5540 35012 5592 35018
rect 5540 34954 5592 34960
rect 5356 34944 5408 34950
rect 5356 34886 5408 34892
rect 5172 34604 5224 34610
rect 5172 34546 5224 34552
rect 5184 34202 5212 34546
rect 5172 34196 5224 34202
rect 5172 34138 5224 34144
rect 5184 34082 5212 34138
rect 5092 34054 5212 34082
rect 5092 33658 5120 34054
rect 5172 33992 5224 33998
rect 5172 33934 5224 33940
rect 5080 33652 5132 33658
rect 5080 33594 5132 33600
rect 5184 32910 5212 33934
rect 5172 32904 5224 32910
rect 5172 32846 5224 32852
rect 5184 32502 5212 32846
rect 5172 32496 5224 32502
rect 5172 32438 5224 32444
rect 5184 31822 5212 32438
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 5368 31754 5396 34886
rect 5736 34474 5764 37318
rect 5908 37266 5960 37272
rect 6000 37324 6052 37330
rect 6000 37266 6052 37272
rect 5908 37188 5960 37194
rect 5908 37130 5960 37136
rect 5920 35834 5948 37130
rect 6196 36582 6224 37606
rect 6276 37460 6328 37466
rect 6276 37402 6328 37408
rect 6184 36576 6236 36582
rect 6184 36518 6236 36524
rect 6196 36174 6224 36518
rect 6184 36168 6236 36174
rect 6184 36110 6236 36116
rect 5908 35828 5960 35834
rect 5908 35770 5960 35776
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 6012 35630 6040 35770
rect 6000 35624 6052 35630
rect 6000 35566 6052 35572
rect 5816 35488 5868 35494
rect 5816 35430 5868 35436
rect 5828 34950 5856 35430
rect 6196 35154 6224 36110
rect 6288 35834 6316 37402
rect 6380 36854 6408 39442
rect 6748 38010 6776 40666
rect 7484 40594 7512 40870
rect 7472 40588 7524 40594
rect 7472 40530 7524 40536
rect 6920 38344 6972 38350
rect 6920 38286 6972 38292
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6748 37466 6776 37946
rect 6828 37800 6880 37806
rect 6828 37742 6880 37748
rect 6840 37618 6868 37742
rect 6932 37738 6960 38286
rect 7012 38276 7064 38282
rect 7012 38218 7064 38224
rect 6920 37732 6972 37738
rect 6920 37674 6972 37680
rect 6840 37590 6960 37618
rect 6736 37460 6788 37466
rect 6736 37402 6788 37408
rect 6368 36848 6420 36854
rect 6420 36808 6500 36836
rect 6368 36790 6420 36796
rect 6276 35828 6328 35834
rect 6276 35770 6328 35776
rect 6184 35148 6236 35154
rect 6184 35090 6236 35096
rect 5816 34944 5868 34950
rect 5816 34886 5868 34892
rect 5724 34468 5776 34474
rect 5644 34428 5724 34456
rect 5644 33590 5672 34428
rect 5724 34410 5776 34416
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 5736 33658 5764 33934
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 5632 33584 5684 33590
rect 5632 33526 5684 33532
rect 5540 33380 5592 33386
rect 5540 33322 5592 33328
rect 5276 31726 5396 31754
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 5184 29850 5212 30670
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 5276 28626 5304 31726
rect 5552 30122 5580 33322
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5644 32910 5672 33254
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5736 31754 5764 32710
rect 5644 31726 5764 31754
rect 5540 30116 5592 30122
rect 5540 30058 5592 30064
rect 5552 29306 5580 30058
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 5644 29186 5672 31726
rect 5828 29646 5856 34886
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 6104 33522 6132 33798
rect 6092 33516 6144 33522
rect 6092 33458 6144 33464
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 5908 32768 5960 32774
rect 5908 32710 5960 32716
rect 5920 31890 5948 32710
rect 6104 32434 6132 32846
rect 6288 32434 6316 35770
rect 6368 33448 6420 33454
rect 6368 33390 6420 33396
rect 6380 33114 6408 33390
rect 6368 33108 6420 33114
rect 6368 33050 6420 33056
rect 6472 32570 6500 36808
rect 6552 36100 6604 36106
rect 6552 36042 6604 36048
rect 6564 35290 6592 36042
rect 6932 36038 6960 37590
rect 7024 37466 7052 38218
rect 7472 37868 7524 37874
rect 7472 37810 7524 37816
rect 7104 37664 7156 37670
rect 7104 37606 7156 37612
rect 7012 37460 7064 37466
rect 7012 37402 7064 37408
rect 7116 37262 7144 37606
rect 7484 37466 7512 37810
rect 7472 37460 7524 37466
rect 7472 37402 7524 37408
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7012 36236 7064 36242
rect 7012 36178 7064 36184
rect 7024 36106 7052 36178
rect 7012 36100 7064 36106
rect 7012 36042 7064 36048
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6932 35630 6960 35974
rect 7012 35692 7064 35698
rect 7012 35634 7064 35640
rect 7104 35692 7156 35698
rect 7104 35634 7156 35640
rect 6920 35624 6972 35630
rect 6920 35566 6972 35572
rect 6920 35488 6972 35494
rect 6920 35430 6972 35436
rect 6932 35290 6960 35430
rect 6552 35284 6604 35290
rect 6552 35226 6604 35232
rect 6920 35284 6972 35290
rect 6920 35226 6972 35232
rect 7024 35170 7052 35634
rect 6932 35142 7052 35170
rect 6932 34950 6960 35142
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 6932 33522 6960 34886
rect 7116 34354 7144 35634
rect 7564 34604 7616 34610
rect 7564 34546 7616 34552
rect 7024 34326 7144 34354
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 7024 33402 7052 34326
rect 7392 33998 7420 34342
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 7380 33992 7432 33998
rect 7380 33934 7432 33940
rect 6828 33380 6880 33386
rect 6828 33322 6880 33328
rect 6932 33374 7052 33402
rect 6840 32570 6868 33322
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 6736 32564 6788 32570
rect 6736 32506 6788 32512
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6092 32428 6144 32434
rect 6276 32428 6328 32434
rect 6092 32370 6144 32376
rect 6196 32388 6276 32416
rect 6196 32026 6224 32388
rect 6276 32370 6328 32376
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6472 31890 6500 32506
rect 6748 32026 6776 32506
rect 6828 32224 6880 32230
rect 6828 32166 6880 32172
rect 6736 32020 6788 32026
rect 6736 31962 6788 31968
rect 5908 31884 5960 31890
rect 5908 31826 5960 31832
rect 6460 31884 6512 31890
rect 6460 31826 6512 31832
rect 6840 31754 6868 32166
rect 6828 31748 6880 31754
rect 6472 31708 6828 31736
rect 6472 31278 6500 31708
rect 6828 31690 6880 31696
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5920 29646 5948 30126
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6380 29850 6408 29990
rect 6368 29844 6420 29850
rect 6368 29786 6420 29792
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5908 29640 5960 29646
rect 5908 29582 5960 29588
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6276 29640 6328 29646
rect 6276 29582 6328 29588
rect 5644 29158 5764 29186
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 5276 28218 5304 28562
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5264 28212 5316 28218
rect 5264 28154 5316 28160
rect 4856 28104 4936 28132
rect 4804 28086 4856 28092
rect 4804 28008 4856 28014
rect 4804 27950 4856 27956
rect 1768 27872 1820 27878
rect 1768 27814 1820 27820
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1780 18902 1808 27814
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4816 27674 4844 27950
rect 5460 27674 5488 28358
rect 5644 28150 5672 28358
rect 5632 28144 5684 28150
rect 5632 28086 5684 28092
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 5448 27668 5500 27674
rect 5448 27610 5500 27616
rect 5552 26994 5580 28018
rect 5644 27674 5672 28086
rect 5736 28082 5764 29158
rect 5828 28529 5856 29582
rect 5920 29306 5948 29582
rect 6104 29306 6132 29582
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 6092 29300 6144 29306
rect 6092 29242 6144 29248
rect 6000 28960 6052 28966
rect 6000 28902 6052 28908
rect 6012 28626 6040 28902
rect 6000 28620 6052 28626
rect 6000 28562 6052 28568
rect 5814 28520 5870 28529
rect 6012 28490 6040 28562
rect 5814 28455 5816 28464
rect 5868 28455 5870 28464
rect 6000 28484 6052 28490
rect 5816 28426 5868 28432
rect 6000 28426 6052 28432
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5632 27668 5684 27674
rect 5632 27610 5684 27616
rect 5828 27554 5856 28426
rect 6196 28218 6224 29582
rect 6288 28642 6316 29582
rect 6288 28614 6408 28642
rect 6380 28422 6408 28614
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6380 28082 6408 28358
rect 6472 28121 6500 31214
rect 6550 30424 6606 30433
rect 6550 30359 6606 30368
rect 6564 30326 6592 30359
rect 6932 30326 6960 33374
rect 7116 33114 7144 33934
rect 7576 33658 7604 34546
rect 7564 33652 7616 33658
rect 7564 33594 7616 33600
rect 7668 33538 7696 42894
rect 7840 42696 7892 42702
rect 7840 42638 7892 42644
rect 7852 41414 7880 42638
rect 7760 41386 7880 41414
rect 7760 36242 7788 41386
rect 7748 36236 7800 36242
rect 7748 36178 7800 36184
rect 7840 36032 7892 36038
rect 7840 35974 7892 35980
rect 7852 35698 7880 35974
rect 7840 35692 7892 35698
rect 7840 35634 7892 35640
rect 7392 33510 7696 33538
rect 7104 33108 7156 33114
rect 7104 33050 7156 33056
rect 7116 32570 7144 33050
rect 7288 32904 7340 32910
rect 7288 32846 7340 32852
rect 7196 32836 7248 32842
rect 7196 32778 7248 32784
rect 7208 32570 7236 32778
rect 7300 32570 7328 32846
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 7196 32564 7248 32570
rect 7196 32506 7248 32512
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7392 32298 7420 33510
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7380 32292 7432 32298
rect 7380 32234 7432 32240
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 7116 31906 7144 31962
rect 7024 31878 7144 31906
rect 7024 31822 7052 31878
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 6644 30320 6696 30326
rect 6644 30262 6696 30268
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6656 29714 6684 30262
rect 6736 30252 6788 30258
rect 6736 30194 6788 30200
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6656 29170 6684 29650
rect 6748 29170 6776 30194
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 6656 29034 6684 29106
rect 6644 29028 6696 29034
rect 6644 28970 6696 28976
rect 6748 28762 6776 29106
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 6826 28656 6882 28665
rect 6826 28591 6882 28600
rect 6840 28558 6868 28591
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6564 28218 6592 28494
rect 6552 28212 6604 28218
rect 6552 28154 6604 28160
rect 6458 28112 6514 28121
rect 6368 28076 6420 28082
rect 6458 28047 6514 28056
rect 6368 28018 6420 28024
rect 6564 27674 6592 28154
rect 6840 28082 6868 28494
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 6552 27668 6604 27674
rect 6552 27610 6604 27616
rect 5644 27526 5856 27554
rect 5644 27402 5672 27526
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 6932 27062 6960 27814
rect 7024 27470 7052 31758
rect 7668 31754 7696 32302
rect 7668 31726 7788 31754
rect 7104 30116 7156 30122
rect 7104 30058 7156 30064
rect 7116 29578 7144 30058
rect 7104 29572 7156 29578
rect 7104 29514 7156 29520
rect 7116 28150 7144 29514
rect 7760 29322 7788 31726
rect 7852 31278 7880 35634
rect 7944 31754 7972 43318
rect 8116 43104 8168 43110
rect 8116 43046 8168 43052
rect 8128 42770 8156 43046
rect 8024 42764 8076 42770
rect 8024 42706 8076 42712
rect 8116 42764 8168 42770
rect 8116 42706 8168 42712
rect 8036 41206 8064 42706
rect 8220 42702 8248 43930
rect 9324 43382 9352 44270
rect 8852 43376 8904 43382
rect 8852 43318 8904 43324
rect 9312 43376 9364 43382
rect 9312 43318 9364 43324
rect 8300 43308 8352 43314
rect 8300 43250 8352 43256
rect 8484 43308 8536 43314
rect 8484 43250 8536 43256
rect 8760 43308 8812 43314
rect 8760 43250 8812 43256
rect 8312 42770 8340 43250
rect 8300 42764 8352 42770
rect 8300 42706 8352 42712
rect 8208 42696 8260 42702
rect 8208 42638 8260 42644
rect 8312 42378 8340 42706
rect 8312 42350 8432 42378
rect 8496 42362 8524 43250
rect 8300 42220 8352 42226
rect 8300 42162 8352 42168
rect 8312 41818 8340 42162
rect 8404 42022 8432 42350
rect 8484 42356 8536 42362
rect 8484 42298 8536 42304
rect 8496 42226 8524 42298
rect 8484 42220 8536 42226
rect 8484 42162 8536 42168
rect 8392 42016 8444 42022
rect 8392 41958 8444 41964
rect 8772 41818 8800 43250
rect 8864 42362 8892 43318
rect 9036 42628 9088 42634
rect 9036 42570 9088 42576
rect 8852 42356 8904 42362
rect 8852 42298 8904 42304
rect 8300 41812 8352 41818
rect 8300 41754 8352 41760
rect 8760 41812 8812 41818
rect 8760 41754 8812 41760
rect 8024 41200 8076 41206
rect 8024 41142 8076 41148
rect 8036 40526 8064 41142
rect 8864 41138 8892 42298
rect 8852 41132 8904 41138
rect 8852 41074 8904 41080
rect 8116 41064 8168 41070
rect 8116 41006 8168 41012
rect 8024 40520 8076 40526
rect 8024 40462 8076 40468
rect 8036 40118 8064 40462
rect 8128 40186 8156 41006
rect 8760 40724 8812 40730
rect 8760 40666 8812 40672
rect 8668 40588 8720 40594
rect 8668 40530 8720 40536
rect 8576 40520 8628 40526
rect 8576 40462 8628 40468
rect 8208 40384 8260 40390
rect 8208 40326 8260 40332
rect 8300 40384 8352 40390
rect 8300 40326 8352 40332
rect 8392 40384 8444 40390
rect 8392 40326 8444 40332
rect 8116 40180 8168 40186
rect 8116 40122 8168 40128
rect 8024 40112 8076 40118
rect 8024 40054 8076 40060
rect 8116 39840 8168 39846
rect 8116 39782 8168 39788
rect 8024 39636 8076 39642
rect 8024 39578 8076 39584
rect 8036 39370 8064 39578
rect 8128 39438 8156 39782
rect 8220 39574 8248 40326
rect 8208 39568 8260 39574
rect 8208 39510 8260 39516
rect 8116 39432 8168 39438
rect 8116 39374 8168 39380
rect 8024 39364 8076 39370
rect 8024 39306 8076 39312
rect 8116 39296 8168 39302
rect 8116 39238 8168 39244
rect 8024 33448 8076 33454
rect 8024 33390 8076 33396
rect 8036 32910 8064 33390
rect 8128 33114 8156 39238
rect 8220 39030 8248 39510
rect 8312 39438 8340 40326
rect 8404 39438 8432 40326
rect 8588 40186 8616 40462
rect 8680 40186 8708 40530
rect 8576 40180 8628 40186
rect 8576 40122 8628 40128
rect 8668 40180 8720 40186
rect 8668 40122 8720 40128
rect 8772 40066 8800 40666
rect 8588 40050 8800 40066
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 8576 40044 8800 40050
rect 8628 40038 8800 40044
rect 8576 39986 8628 39992
rect 8300 39432 8352 39438
rect 8300 39374 8352 39380
rect 8392 39432 8444 39438
rect 8392 39374 8444 39380
rect 8208 39024 8260 39030
rect 8208 38966 8260 38972
rect 8404 38962 8432 39374
rect 8496 39302 8524 39986
rect 8588 39642 8616 39986
rect 8576 39636 8628 39642
rect 8576 39578 8628 39584
rect 9048 39438 9076 42570
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 9140 42294 9168 42502
rect 9128 42288 9180 42294
rect 9128 42230 9180 42236
rect 9128 41540 9180 41546
rect 9128 41482 9180 41488
rect 8944 39432 8996 39438
rect 8944 39374 8996 39380
rect 9036 39432 9088 39438
rect 9036 39374 9088 39380
rect 8484 39296 8536 39302
rect 8484 39238 8536 39244
rect 8496 39098 8524 39238
rect 8484 39092 8536 39098
rect 8484 39034 8536 39040
rect 8392 38956 8444 38962
rect 8392 38898 8444 38904
rect 8208 38752 8260 38758
rect 8208 38694 8260 38700
rect 8220 38350 8248 38694
rect 8208 38344 8260 38350
rect 8208 38286 8260 38292
rect 8956 38010 8984 39374
rect 9036 39296 9088 39302
rect 9036 39238 9088 39244
rect 9048 38010 9076 39238
rect 9140 38010 9168 41482
rect 9312 41472 9364 41478
rect 9312 41414 9364 41420
rect 9404 41472 9456 41478
rect 9404 41414 9456 41420
rect 10060 41414 10088 44678
rect 10152 44538 10180 45426
rect 11520 45280 11572 45286
rect 11520 45222 11572 45228
rect 11532 45082 11560 45222
rect 11520 45076 11572 45082
rect 11520 45018 11572 45024
rect 10508 44804 10560 44810
rect 10508 44746 10560 44752
rect 10140 44532 10192 44538
rect 10140 44474 10192 44480
rect 10520 44266 10548 44746
rect 11716 44538 11744 45426
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 11980 44940 12032 44946
rect 11980 44882 12032 44888
rect 11704 44532 11756 44538
rect 11704 44474 11756 44480
rect 11244 44464 11296 44470
rect 11244 44406 11296 44412
rect 10692 44396 10744 44402
rect 10692 44338 10744 44344
rect 10508 44260 10560 44266
rect 10508 44202 10560 44208
rect 10704 43994 10732 44338
rect 10692 43988 10744 43994
rect 10692 43930 10744 43936
rect 10692 43240 10744 43246
rect 10692 43182 10744 43188
rect 10600 42696 10652 42702
rect 10600 42638 10652 42644
rect 10612 42294 10640 42638
rect 10600 42288 10652 42294
rect 10600 42230 10652 42236
rect 10612 42106 10640 42230
rect 9324 41274 9352 41414
rect 9416 41386 9628 41414
rect 9312 41268 9364 41274
rect 9312 41210 9364 41216
rect 9220 40384 9272 40390
rect 9220 40326 9272 40332
rect 9232 39982 9260 40326
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 9404 38888 9456 38894
rect 9404 38830 9456 38836
rect 9416 38554 9444 38830
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 9220 38344 9272 38350
rect 9220 38286 9272 38292
rect 9232 38010 9260 38286
rect 8944 38004 8996 38010
rect 8944 37946 8996 37952
rect 9036 38004 9088 38010
rect 9036 37946 9088 37952
rect 9128 38004 9180 38010
rect 9128 37946 9180 37952
rect 9220 38004 9272 38010
rect 9220 37946 9272 37952
rect 9128 37800 9180 37806
rect 9404 37800 9456 37806
rect 9180 37760 9260 37788
rect 9128 37742 9180 37748
rect 8668 37664 8720 37670
rect 8668 37606 8720 37612
rect 8680 37262 8708 37606
rect 8668 37256 8720 37262
rect 8668 37198 8720 37204
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 8312 35698 8340 36518
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8392 36100 8444 36106
rect 8392 36042 8444 36048
rect 8300 35692 8352 35698
rect 8300 35634 8352 35640
rect 8404 35630 8432 36042
rect 8956 35698 8984 36178
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 8576 34604 8628 34610
rect 8576 34546 8628 34552
rect 8588 33658 8616 34546
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8760 34400 8812 34406
rect 8760 34342 8812 34348
rect 8772 33998 8800 34342
rect 8864 34202 8892 34478
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8956 34066 8984 35634
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 9128 33856 9180 33862
rect 9128 33798 9180 33804
rect 9140 33658 9168 33798
rect 8576 33652 8628 33658
rect 8576 33594 8628 33600
rect 9128 33652 9180 33658
rect 9128 33594 9180 33600
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 9232 33046 9260 37760
rect 9404 37742 9456 37748
rect 9312 36032 9364 36038
rect 9312 35974 9364 35980
rect 9324 35290 9352 35974
rect 9416 35834 9444 37742
rect 9496 36780 9548 36786
rect 9496 36722 9548 36728
rect 9508 36038 9536 36722
rect 9600 36174 9628 41386
rect 9968 41386 10088 41414
rect 10428 42078 10640 42106
rect 9772 40180 9824 40186
rect 9772 40122 9824 40128
rect 9784 39642 9812 40122
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 9772 36304 9824 36310
rect 9772 36246 9824 36252
rect 9588 36168 9640 36174
rect 9588 36110 9640 36116
rect 9496 36032 9548 36038
rect 9496 35974 9548 35980
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9312 35284 9364 35290
rect 9312 35226 9364 35232
rect 9416 33454 9444 35770
rect 9508 35766 9536 35974
rect 9496 35760 9548 35766
rect 9496 35702 9548 35708
rect 9508 35018 9536 35702
rect 9600 35494 9628 36110
rect 9784 36038 9812 36246
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9772 36032 9824 36038
rect 9772 35974 9824 35980
rect 9692 35630 9720 35974
rect 9784 35766 9812 35974
rect 9772 35760 9824 35766
rect 9772 35702 9824 35708
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9876 35290 9904 36110
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9496 35012 9548 35018
rect 9496 34954 9548 34960
rect 9968 34490 9996 41386
rect 10428 41206 10456 42078
rect 10704 42022 10732 43182
rect 11060 42628 11112 42634
rect 11060 42570 11112 42576
rect 11072 42362 11100 42570
rect 11256 42362 11284 44406
rect 11992 43790 12020 44882
rect 12164 44736 12216 44742
rect 12164 44678 12216 44684
rect 12176 44538 12204 44678
rect 12164 44532 12216 44538
rect 12164 44474 12216 44480
rect 12544 44334 12572 45358
rect 13556 45082 13584 45426
rect 13544 45076 13596 45082
rect 13544 45018 13596 45024
rect 12900 44940 12952 44946
rect 12900 44882 12952 44888
rect 12912 44538 12940 44882
rect 13268 44736 13320 44742
rect 13268 44678 13320 44684
rect 12900 44532 12952 44538
rect 12900 44474 12952 44480
rect 12532 44328 12584 44334
rect 12532 44270 12584 44276
rect 13176 44328 13228 44334
rect 13176 44270 13228 44276
rect 12440 44192 12492 44198
rect 12440 44134 12492 44140
rect 12452 43790 12480 44134
rect 11980 43784 12032 43790
rect 11980 43726 12032 43732
rect 12440 43784 12492 43790
rect 12440 43726 12492 43732
rect 11796 42764 11848 42770
rect 11796 42706 11848 42712
rect 11704 42560 11756 42566
rect 11704 42502 11756 42508
rect 11060 42356 11112 42362
rect 11060 42298 11112 42304
rect 11244 42356 11296 42362
rect 11244 42298 11296 42304
rect 10784 42288 10836 42294
rect 10784 42230 10836 42236
rect 10692 42016 10744 42022
rect 10692 41958 10744 41964
rect 10796 41818 10824 42230
rect 11072 42226 11100 42298
rect 11060 42220 11112 42226
rect 11060 42162 11112 42168
rect 10784 41812 10836 41818
rect 10784 41754 10836 41760
rect 11072 41546 11100 42162
rect 11520 42152 11572 42158
rect 11520 42094 11572 42100
rect 11152 42016 11204 42022
rect 11152 41958 11204 41964
rect 11164 41818 11192 41958
rect 11532 41818 11560 42094
rect 11716 41818 11744 42502
rect 11152 41812 11204 41818
rect 11152 41754 11204 41760
rect 11520 41812 11572 41818
rect 11520 41754 11572 41760
rect 11704 41812 11756 41818
rect 11704 41754 11756 41760
rect 11808 41750 11836 42706
rect 11888 42356 11940 42362
rect 11888 42298 11940 42304
rect 11796 41744 11848 41750
rect 11796 41686 11848 41692
rect 11900 41682 11928 42298
rect 11992 42226 12020 43726
rect 12544 43722 12572 44270
rect 13188 43858 13216 44270
rect 13280 44198 13308 44678
rect 13452 44328 13504 44334
rect 13452 44270 13504 44276
rect 13268 44192 13320 44198
rect 13268 44134 13320 44140
rect 13176 43852 13228 43858
rect 13176 43794 13228 43800
rect 12532 43716 12584 43722
rect 12532 43658 12584 43664
rect 12900 43716 12952 43722
rect 12900 43658 12952 43664
rect 12808 42696 12860 42702
rect 12808 42638 12860 42644
rect 11980 42220 12032 42226
rect 11980 42162 12032 42168
rect 12256 42016 12308 42022
rect 12256 41958 12308 41964
rect 11888 41676 11940 41682
rect 11888 41618 11940 41624
rect 10508 41540 10560 41546
rect 10508 41482 10560 41488
rect 11060 41540 11112 41546
rect 11060 41482 11112 41488
rect 10520 41274 10548 41482
rect 10508 41268 10560 41274
rect 10508 41210 10560 41216
rect 10416 41200 10468 41206
rect 10416 41142 10468 41148
rect 10048 40452 10100 40458
rect 10048 40394 10100 40400
rect 10060 39982 10088 40394
rect 10428 40186 10456 41142
rect 10416 40180 10468 40186
rect 10416 40122 10468 40128
rect 11072 39982 11100 41482
rect 11244 41472 11296 41478
rect 11244 41414 11296 41420
rect 11256 41206 11284 41414
rect 11900 41274 11928 41618
rect 12268 41614 12296 41958
rect 12820 41818 12848 42638
rect 12808 41812 12860 41818
rect 12808 41754 12860 41760
rect 12256 41608 12308 41614
rect 12256 41550 12308 41556
rect 12912 41414 12940 43658
rect 13176 43104 13228 43110
rect 13176 43046 13228 43052
rect 13188 42294 13216 43046
rect 13176 42288 13228 42294
rect 13176 42230 13228 42236
rect 12820 41386 12940 41414
rect 11888 41268 11940 41274
rect 11888 41210 11940 41216
rect 11244 41200 11296 41206
rect 11244 41142 11296 41148
rect 11980 41064 12032 41070
rect 11980 41006 12032 41012
rect 12164 41064 12216 41070
rect 12164 41006 12216 41012
rect 11796 40724 11848 40730
rect 11796 40666 11848 40672
rect 11152 40520 11204 40526
rect 11152 40462 11204 40468
rect 11164 40050 11192 40462
rect 11808 40458 11836 40666
rect 11796 40452 11848 40458
rect 11796 40394 11848 40400
rect 11888 40452 11940 40458
rect 11888 40394 11940 40400
rect 11900 40186 11928 40394
rect 11888 40180 11940 40186
rect 11888 40122 11940 40128
rect 11152 40044 11204 40050
rect 11152 39986 11204 39992
rect 10048 39976 10100 39982
rect 10048 39918 10100 39924
rect 11060 39976 11112 39982
rect 11060 39918 11112 39924
rect 10060 39506 10088 39918
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10048 39500 10100 39506
rect 10048 39442 10100 39448
rect 10796 39438 10824 39782
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 10048 38956 10100 38962
rect 10048 38898 10100 38904
rect 10060 38010 10088 38898
rect 10796 38418 10824 39374
rect 11520 39364 11572 39370
rect 11520 39306 11572 39312
rect 11532 39098 11560 39306
rect 11900 39098 11928 40122
rect 11520 39092 11572 39098
rect 11520 39034 11572 39040
rect 11888 39092 11940 39098
rect 11888 39034 11940 39040
rect 10784 38412 10836 38418
rect 10784 38354 10836 38360
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 10048 38004 10100 38010
rect 10048 37946 10100 37952
rect 10244 36038 10272 38218
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 11256 37942 11284 38150
rect 11244 37936 11296 37942
rect 11244 37878 11296 37884
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 11152 36780 11204 36786
rect 11152 36722 11204 36728
rect 10704 36378 10732 36722
rect 11060 36576 11112 36582
rect 11060 36518 11112 36524
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 11072 36242 11100 36518
rect 11060 36236 11112 36242
rect 11060 36178 11112 36184
rect 11164 36122 11192 36722
rect 11072 36106 11192 36122
rect 11060 36100 11192 36106
rect 11112 36094 11192 36100
rect 11060 36042 11112 36048
rect 10232 36032 10284 36038
rect 10232 35974 10284 35980
rect 11072 35630 11100 36042
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10704 35290 10732 35430
rect 10692 35284 10744 35290
rect 10692 35226 10744 35232
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 9968 34462 10088 34490
rect 9496 34400 9548 34406
rect 9496 34342 9548 34348
rect 9956 34400 10008 34406
rect 9956 34342 10008 34348
rect 9508 33658 9536 34342
rect 9968 33930 9996 34342
rect 9956 33924 10008 33930
rect 9956 33866 10008 33872
rect 9496 33652 9548 33658
rect 9496 33594 9548 33600
rect 9404 33448 9456 33454
rect 9404 33390 9456 33396
rect 9588 33312 9640 33318
rect 9588 33254 9640 33260
rect 9220 33040 9272 33046
rect 9220 32982 9272 32988
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 8036 32570 8064 32846
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 8392 32564 8444 32570
rect 8392 32506 8444 32512
rect 8404 31822 8432 32506
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 8392 31816 8444 31822
rect 8392 31758 8444 31764
rect 7944 31726 8064 31754
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7760 29294 7972 29322
rect 7944 28966 7972 29294
rect 7932 28960 7984 28966
rect 7932 28902 7984 28908
rect 7944 28762 7972 28902
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7944 28558 7972 28698
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7944 28234 7972 28494
rect 7852 28218 7972 28234
rect 7840 28212 7972 28218
rect 7892 28206 7972 28212
rect 7840 28154 7892 28160
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7116 27062 7144 28086
rect 6920 27056 6972 27062
rect 6920 26998 6972 27004
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 7116 26042 7144 26998
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 7760 25498 7788 25774
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 8036 24410 8064 31726
rect 8312 31346 8340 31758
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8312 30870 8340 31078
rect 8300 30864 8352 30870
rect 8300 30806 8352 30812
rect 8680 30394 8708 31282
rect 8956 30938 8984 31282
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8956 30734 8984 30874
rect 9048 30802 9076 31282
rect 9036 30796 9088 30802
rect 9036 30738 9088 30744
rect 8944 30728 8996 30734
rect 8944 30670 8996 30676
rect 8668 30388 8720 30394
rect 8668 30330 8720 30336
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 8300 28688 8352 28694
rect 8300 28630 8352 28636
rect 8312 28422 8340 28630
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8128 27985 8156 28018
rect 8114 27976 8170 27985
rect 8114 27911 8170 27920
rect 8128 26858 8156 27911
rect 8312 27674 8340 28358
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8404 27334 8432 27814
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8220 26994 8248 27270
rect 8496 27130 8524 28494
rect 8680 28490 8708 28562
rect 8942 28520 8998 28529
rect 8576 28484 8628 28490
rect 8576 28426 8628 28432
rect 8668 28484 8720 28490
rect 8942 28455 8944 28464
rect 8668 28426 8720 28432
rect 8996 28455 8998 28464
rect 8944 28426 8996 28432
rect 8588 27130 8616 28426
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28218 9076 28358
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 8852 27668 8904 27674
rect 8852 27610 8904 27616
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 8576 27124 8628 27130
rect 8576 27066 8628 27072
rect 8864 26994 8892 27610
rect 9048 27130 9076 27950
rect 9140 27674 9168 28698
rect 9232 28626 9260 32982
rect 9600 32502 9628 33254
rect 9588 32496 9640 32502
rect 9588 32438 9640 32444
rect 9496 32224 9548 32230
rect 9496 32166 9548 32172
rect 9508 31822 9536 32166
rect 9496 31816 9548 31822
rect 9496 31758 9548 31764
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 9324 31482 9352 31690
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9312 31476 9364 31482
rect 9312 31418 9364 31424
rect 9416 31210 9444 31622
rect 9692 31482 9720 31758
rect 9864 31680 9916 31686
rect 9864 31622 9916 31628
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9496 31340 9548 31346
rect 9496 31282 9548 31288
rect 9404 31204 9456 31210
rect 9404 31146 9456 31152
rect 9416 30938 9444 31146
rect 9312 30932 9364 30938
rect 9312 30874 9364 30880
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9220 28620 9272 28626
rect 9220 28562 9272 28568
rect 9232 28150 9260 28562
rect 9220 28144 9272 28150
rect 9220 28086 9272 28092
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 9232 27470 9260 28086
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9036 27124 9088 27130
rect 9036 27066 9088 27072
rect 9232 26994 9260 27406
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 8116 26852 8168 26858
rect 8116 26794 8168 26800
rect 8220 25702 8248 26930
rect 9324 25702 9352 30874
rect 9508 30802 9536 31282
rect 9876 31278 9904 31622
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9600 30734 9628 31214
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9600 30394 9628 30670
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 29028 9548 29034
rect 9496 28970 9548 28976
rect 9508 28626 9536 28970
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9416 27470 9444 28154
rect 9692 27470 9720 28358
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9416 26926 9444 27406
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 8208 25696 8260 25702
rect 8208 25638 8260 25644
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9324 25294 9352 25638
rect 9692 25498 9720 25774
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 9784 24070 9812 30670
rect 9876 30598 9904 31214
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9968 28082 9996 33866
rect 10060 32910 10088 34462
rect 10244 33969 10272 34546
rect 10230 33960 10286 33969
rect 10152 33918 10230 33946
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 10060 32434 10088 32846
rect 10152 32570 10180 33918
rect 10230 33895 10286 33904
rect 10876 33924 10928 33930
rect 10876 33866 10928 33872
rect 10888 33658 10916 33866
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 10980 33454 11008 33798
rect 11256 33658 11284 37878
rect 11992 36378 12020 41006
rect 12176 38894 12204 41006
rect 12256 40384 12308 40390
rect 12256 40326 12308 40332
rect 12268 40118 12296 40326
rect 12256 40112 12308 40118
rect 12256 40054 12308 40060
rect 12820 39982 12848 41386
rect 12440 39976 12492 39982
rect 12440 39918 12492 39924
rect 12808 39976 12860 39982
rect 12808 39918 12860 39924
rect 12992 39976 13044 39982
rect 12992 39918 13044 39924
rect 12452 39642 12480 39918
rect 12440 39636 12492 39642
rect 12440 39578 12492 39584
rect 12348 39024 12400 39030
rect 12348 38966 12400 38972
rect 12164 38888 12216 38894
rect 12164 38830 12216 38836
rect 11980 36372 12032 36378
rect 11980 36314 12032 36320
rect 11992 35630 12020 36314
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 12256 34944 12308 34950
rect 12256 34886 12308 34892
rect 11612 33856 11664 33862
rect 11612 33798 11664 33804
rect 11888 33856 11940 33862
rect 11888 33798 11940 33804
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 11624 33522 11652 33798
rect 11900 33522 11928 33798
rect 12162 33688 12218 33697
rect 12162 33623 12164 33632
rect 12216 33623 12218 33632
rect 12164 33594 12216 33600
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10968 33448 11020 33454
rect 10968 33390 11020 33396
rect 10232 32768 10284 32774
rect 10232 32710 10284 32716
rect 10244 32570 10272 32710
rect 10140 32564 10192 32570
rect 10140 32506 10192 32512
rect 10232 32564 10284 32570
rect 10232 32506 10284 32512
rect 10244 32434 10272 32506
rect 10048 32428 10100 32434
rect 10048 32370 10100 32376
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 10140 32292 10192 32298
rect 10140 32234 10192 32240
rect 10152 31958 10180 32234
rect 10324 32224 10376 32230
rect 10324 32166 10376 32172
rect 10336 32026 10364 32166
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10140 31952 10192 31958
rect 10140 31894 10192 31900
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 10060 31686 10088 31758
rect 10048 31680 10100 31686
rect 10048 31622 10100 31628
rect 10152 31498 10180 31894
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 10060 31470 10180 31498
rect 10244 31482 10272 31758
rect 10324 31748 10376 31754
rect 10324 31690 10376 31696
rect 10336 31482 10364 31690
rect 10232 31476 10284 31482
rect 10060 31414 10088 31470
rect 10232 31418 10284 31424
rect 10324 31476 10376 31482
rect 10324 31418 10376 31424
rect 10048 31408 10100 31414
rect 10048 31350 10100 31356
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 10244 30734 10272 31282
rect 10520 31142 10548 31282
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 10612 28558 10640 33390
rect 11072 33046 11100 33458
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11060 33040 11112 33046
rect 11060 32982 11112 32988
rect 11256 32774 11284 33390
rect 11716 32978 11744 33458
rect 11900 33114 11928 33458
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 11888 33108 11940 33114
rect 11888 33050 11940 33056
rect 11704 32972 11756 32978
rect 11704 32914 11756 32920
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11244 32768 11296 32774
rect 11244 32710 11296 32716
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10888 30870 10916 31282
rect 11256 30870 11284 32710
rect 11624 32026 11652 32846
rect 11612 32020 11664 32026
rect 11612 31962 11664 31968
rect 11992 31822 12020 33254
rect 12164 32428 12216 32434
rect 12164 32370 12216 32376
rect 12176 31822 12204 32370
rect 12268 32366 12296 34886
rect 12256 32360 12308 32366
rect 12256 32302 12308 32308
rect 12268 31890 12296 32302
rect 12360 32026 12388 38966
rect 12532 37936 12584 37942
rect 12532 37878 12584 37884
rect 12544 37466 12572 37878
rect 12820 37806 12848 39918
rect 13004 39098 13032 39918
rect 12992 39092 13044 39098
rect 12992 39034 13044 39040
rect 12808 37800 12860 37806
rect 12808 37742 12860 37748
rect 12532 37460 12584 37466
rect 12532 37402 12584 37408
rect 12808 37256 12860 37262
rect 12808 37198 12860 37204
rect 12820 36922 12848 37198
rect 12808 36916 12860 36922
rect 12808 36858 12860 36864
rect 12440 36848 12492 36854
rect 12440 36790 12492 36796
rect 12452 35222 12480 36790
rect 12900 36780 12952 36786
rect 12900 36722 12952 36728
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 12912 36242 12940 36722
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 12820 36038 12848 36110
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 12912 35834 12940 36178
rect 12992 36168 13044 36174
rect 12992 36110 13044 36116
rect 12900 35828 12952 35834
rect 12900 35770 12952 35776
rect 12532 35624 12584 35630
rect 12532 35566 12584 35572
rect 12440 35216 12492 35222
rect 12440 35158 12492 35164
rect 12440 34468 12492 34474
rect 12440 34410 12492 34416
rect 12452 34066 12480 34410
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12544 33504 12572 35566
rect 12900 34400 12952 34406
rect 12900 34342 12952 34348
rect 12912 33998 12940 34342
rect 12900 33992 12952 33998
rect 12900 33934 12952 33940
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 12820 33658 12848 33798
rect 12808 33652 12860 33658
rect 12808 33594 12860 33600
rect 12452 33476 12572 33504
rect 12452 32434 12480 33476
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 12728 32570 12756 32710
rect 12716 32564 12768 32570
rect 12716 32506 12768 32512
rect 12440 32428 12492 32434
rect 12440 32370 12492 32376
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 11980 31816 12032 31822
rect 11980 31758 12032 31764
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12346 31784 12402 31793
rect 12256 31748 12308 31754
rect 12346 31719 12402 31728
rect 12256 31690 12308 31696
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 10876 30864 10928 30870
rect 10876 30806 10928 30812
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10796 29170 10824 29446
rect 10888 29238 10916 30262
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10704 28762 10732 29106
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9968 25974 9996 28018
rect 10232 26240 10284 26246
rect 10232 26182 10284 26188
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 10244 25430 10272 26182
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10336 25362 10364 25638
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10612 24154 10640 28494
rect 10888 26382 10916 29174
rect 11072 28966 11100 30670
rect 11152 30592 11204 30598
rect 11152 30534 11204 30540
rect 11164 30326 11192 30534
rect 11152 30320 11204 30326
rect 11152 30262 11204 30268
rect 11256 29850 11284 30806
rect 11900 30734 11928 30874
rect 12268 30734 12296 31690
rect 12360 31346 12388 31719
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12440 31204 12492 31210
rect 12440 31146 12492 31152
rect 11888 30728 11940 30734
rect 12256 30728 12308 30734
rect 11888 30670 11940 30676
rect 12254 30696 12256 30705
rect 12308 30696 12310 30705
rect 12254 30631 12310 30640
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11348 30433 11376 30534
rect 11334 30424 11390 30433
rect 11334 30359 11390 30368
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11348 29306 11376 30194
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11440 29170 11468 29446
rect 12268 29170 12296 29650
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 11428 29164 11480 29170
rect 11428 29106 11480 29112
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11072 28626 11100 28902
rect 11256 28762 11284 29106
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11060 28008 11112 28014
rect 11060 27950 11112 27956
rect 11336 28008 11388 28014
rect 11336 27950 11388 27956
rect 11072 27674 11100 27950
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 11348 27538 11376 27950
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10888 25838 10916 26318
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 11256 25498 11284 26386
rect 11244 25492 11296 25498
rect 11244 25434 11296 25440
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10888 24954 10916 25162
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 10980 24206 11008 24278
rect 11072 24206 11100 24346
rect 11256 24274 11284 25434
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10968 24200 11020 24206
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 8588 23118 8616 23462
rect 9232 23118 9260 24006
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 8588 22710 8616 23054
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8956 22574 8984 22918
rect 9784 22778 9812 24006
rect 10244 23186 10272 24006
rect 10428 23866 10456 24142
rect 10612 24126 10732 24154
rect 10968 24142 11020 24148
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10612 23118 10640 24006
rect 10704 23866 10732 24126
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 8944 22568 8996 22574
rect 8944 22510 8996 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 10612 22094 10640 23054
rect 10980 22710 11008 24142
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11072 23322 11100 23802
rect 11256 23662 11284 24210
rect 11244 23656 11296 23662
rect 11242 23624 11244 23633
rect 11296 23624 11298 23633
rect 11242 23559 11298 23568
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10612 22066 10824 22094
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 10796 20942 10824 22066
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9784 20602 9812 20810
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19514 10732 19722
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 6932 17814 6960 18566
rect 9232 18426 9260 18566
rect 10244 18426 10272 18566
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 10060 17610 10088 18022
rect 10796 17610 10824 20878
rect 11256 20398 11284 23559
rect 11440 21146 11468 29106
rect 12452 28150 12480 31146
rect 12544 30410 12572 31282
rect 12544 30394 12664 30410
rect 12532 30388 12664 30394
rect 12584 30382 12664 30388
rect 12532 30330 12584 30336
rect 12532 30184 12584 30190
rect 12532 30126 12584 30132
rect 12544 29306 12572 30126
rect 12636 29850 12664 30382
rect 12728 30054 12756 32166
rect 12808 31952 12860 31958
rect 12808 31894 12860 31900
rect 12820 31278 12848 31894
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12912 31142 12940 32982
rect 13004 32910 13032 36110
rect 13096 36038 13124 36722
rect 13084 36032 13136 36038
rect 13084 35974 13136 35980
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 13004 32366 13032 32846
rect 12992 32360 13044 32366
rect 12992 32302 13044 32308
rect 13096 31754 13124 35974
rect 13176 35216 13228 35222
rect 13176 35158 13228 35164
rect 13188 34490 13216 35158
rect 13280 34746 13308 44134
rect 13360 43308 13412 43314
rect 13360 43250 13412 43256
rect 13372 41818 13400 43250
rect 13360 41812 13412 41818
rect 13360 41754 13412 41760
rect 13360 41472 13412 41478
rect 13360 41414 13412 41420
rect 13372 37670 13400 41414
rect 13360 37664 13412 37670
rect 13360 37606 13412 37612
rect 13372 36786 13400 37606
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 13268 34740 13320 34746
rect 13268 34682 13320 34688
rect 13280 34610 13308 34682
rect 13464 34626 13492 44270
rect 13740 44198 13768 45494
rect 13820 44872 13872 44878
rect 13820 44814 13872 44820
rect 13728 44192 13780 44198
rect 13728 44134 13780 44140
rect 13740 42702 13768 44134
rect 13832 43994 13860 44814
rect 13820 43988 13872 43994
rect 13820 43930 13872 43936
rect 13728 42696 13780 42702
rect 13728 42638 13780 42644
rect 13544 42560 13596 42566
rect 13544 42502 13596 42508
rect 13556 42226 13584 42502
rect 13544 42220 13596 42226
rect 13544 42162 13596 42168
rect 13740 42158 13768 42638
rect 13912 42628 13964 42634
rect 13912 42570 13964 42576
rect 13924 42362 13952 42570
rect 13912 42356 13964 42362
rect 13912 42298 13964 42304
rect 13728 42152 13780 42158
rect 13728 42094 13780 42100
rect 13636 41676 13688 41682
rect 13636 41618 13688 41624
rect 13648 40934 13676 41618
rect 13740 41478 13768 42094
rect 13728 41472 13780 41478
rect 13728 41414 13780 41420
rect 14016 41414 14044 45766
rect 14844 45554 14872 45902
rect 15936 45892 15988 45898
rect 15936 45834 15988 45840
rect 15948 45558 15976 45834
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 14660 45526 14872 45554
rect 15936 45552 15988 45558
rect 14464 45008 14516 45014
rect 14464 44950 14516 44956
rect 14476 44334 14504 44950
rect 14660 44538 14688 45526
rect 15936 45494 15988 45500
rect 16304 45552 16356 45558
rect 16304 45494 16356 45500
rect 16488 45552 16540 45558
rect 21836 45554 21864 45970
rect 23860 45966 23888 47681
rect 33060 46866 33088 47790
rect 41878 47681 41934 48481
rect 33060 46838 33180 46866
rect 24124 46028 24176 46034
rect 24124 45970 24176 45976
rect 22192 45960 22244 45966
rect 22192 45902 22244 45908
rect 23848 45960 23900 45966
rect 23848 45902 23900 45908
rect 22204 45626 22232 45902
rect 22192 45620 22244 45626
rect 22192 45562 22244 45568
rect 21836 45526 22048 45554
rect 16488 45494 16540 45500
rect 14740 45280 14792 45286
rect 14740 45222 14792 45228
rect 14752 44946 14780 45222
rect 14740 44940 14792 44946
rect 14740 44882 14792 44888
rect 15292 44940 15344 44946
rect 15292 44882 15344 44888
rect 14648 44532 14700 44538
rect 14648 44474 14700 44480
rect 14464 44328 14516 44334
rect 14464 44270 14516 44276
rect 14660 43738 14688 44474
rect 14752 43790 14780 44882
rect 14832 44532 14884 44538
rect 14832 44474 14884 44480
rect 14844 44266 14872 44474
rect 14832 44260 14884 44266
rect 14832 44202 14884 44208
rect 15304 43858 15332 44882
rect 15384 44396 15436 44402
rect 15384 44338 15436 44344
rect 15396 43994 15424 44338
rect 15384 43988 15436 43994
rect 15384 43930 15436 43936
rect 15292 43852 15344 43858
rect 15292 43794 15344 43800
rect 14476 43710 14688 43738
rect 14740 43784 14792 43790
rect 14740 43726 14792 43732
rect 14476 43654 14504 43710
rect 14464 43648 14516 43654
rect 14464 43590 14516 43596
rect 14556 43648 14608 43654
rect 14556 43590 14608 43596
rect 14568 42906 14596 43590
rect 14556 42900 14608 42906
rect 14556 42842 14608 42848
rect 14096 42560 14148 42566
rect 14096 42502 14148 42508
rect 14188 42560 14240 42566
rect 14188 42502 14240 42508
rect 14108 42362 14136 42502
rect 14096 42356 14148 42362
rect 14096 42298 14148 42304
rect 14200 42022 14228 42502
rect 14464 42288 14516 42294
rect 14464 42230 14516 42236
rect 14188 42016 14240 42022
rect 14188 41958 14240 41964
rect 14016 41386 14136 41414
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 13728 40520 13780 40526
rect 13728 40462 13780 40468
rect 13740 40186 13768 40462
rect 13912 40384 13964 40390
rect 13912 40326 13964 40332
rect 13728 40180 13780 40186
rect 13728 40122 13780 40128
rect 13924 39982 13952 40326
rect 13912 39976 13964 39982
rect 13912 39918 13964 39924
rect 13544 39840 13596 39846
rect 13544 39782 13596 39788
rect 13636 39840 13688 39846
rect 13636 39782 13688 39788
rect 13556 39642 13584 39782
rect 13544 39636 13596 39642
rect 13544 39578 13596 39584
rect 13648 39506 13676 39782
rect 13636 39500 13688 39506
rect 13636 39442 13688 39448
rect 13820 39296 13872 39302
rect 13820 39238 13872 39244
rect 13832 39098 13860 39238
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 13728 37120 13780 37126
rect 13728 37062 13780 37068
rect 13740 36802 13768 37062
rect 13740 36786 13860 36802
rect 13740 36780 13872 36786
rect 13740 36774 13820 36780
rect 13544 36712 13596 36718
rect 13544 36654 13596 36660
rect 13556 36174 13584 36654
rect 13740 36650 13768 36774
rect 13820 36722 13872 36728
rect 13728 36644 13780 36650
rect 13728 36586 13780 36592
rect 13636 36576 13688 36582
rect 13636 36518 13688 36524
rect 13648 36242 13676 36518
rect 13740 36378 13768 36586
rect 13728 36372 13780 36378
rect 13728 36314 13780 36320
rect 13820 36304 13872 36310
rect 13820 36246 13872 36252
rect 13636 36236 13688 36242
rect 13636 36178 13688 36184
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 13372 34610 13492 34626
rect 13268 34604 13320 34610
rect 13268 34546 13320 34552
rect 13360 34604 13492 34610
rect 13412 34598 13492 34604
rect 13360 34546 13412 34552
rect 13188 34462 13492 34490
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13176 32564 13228 32570
rect 13176 32506 13228 32512
rect 13188 32434 13216 32506
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13176 31952 13228 31958
rect 13174 31920 13176 31929
rect 13228 31920 13230 31929
rect 13174 31855 13230 31864
rect 13004 31726 13124 31754
rect 13004 31278 13032 31726
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 12808 31136 12860 31142
rect 12808 31078 12860 31084
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12820 30938 12848 31078
rect 12808 30932 12860 30938
rect 12808 30874 12860 30880
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 12820 30546 12848 30738
rect 12900 30728 12952 30734
rect 13004 30682 13032 31214
rect 12952 30676 13032 30682
rect 12900 30670 13032 30676
rect 12912 30654 13032 30670
rect 13096 30546 13124 31282
rect 13176 31136 13228 31142
rect 13176 31078 13228 31084
rect 13188 30802 13216 31078
rect 13176 30796 13228 30802
rect 13176 30738 13228 30744
rect 12820 30518 13124 30546
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 12912 28762 12940 29038
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12716 28688 12768 28694
rect 12530 28656 12586 28665
rect 12716 28630 12768 28636
rect 12530 28591 12586 28600
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 12452 27985 12480 28086
rect 12438 27976 12494 27985
rect 12544 27946 12572 28591
rect 12728 28150 12756 28630
rect 13096 28558 13124 29106
rect 13188 28937 13216 29106
rect 13280 28966 13308 32710
rect 13372 31482 13400 33934
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13464 30938 13492 34462
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13556 32978 13584 33934
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13556 32416 13584 32914
rect 13648 32774 13676 36178
rect 13832 35834 13860 36246
rect 13912 36168 13964 36174
rect 13912 36110 13964 36116
rect 13924 35834 13952 36110
rect 14004 36032 14056 36038
rect 14004 35974 14056 35980
rect 13820 35828 13872 35834
rect 13820 35770 13872 35776
rect 13912 35828 13964 35834
rect 13912 35770 13964 35776
rect 14016 35766 14044 35974
rect 14004 35760 14056 35766
rect 14004 35702 14056 35708
rect 14108 35612 14136 41386
rect 14200 41274 14228 41958
rect 14280 41676 14332 41682
rect 14280 41618 14332 41624
rect 14188 41268 14240 41274
rect 14188 41210 14240 41216
rect 14292 41138 14320 41618
rect 14280 41132 14332 41138
rect 14280 41074 14332 41080
rect 14476 40526 14504 42230
rect 14568 41614 14596 42842
rect 14740 42764 14792 42770
rect 14740 42706 14792 42712
rect 14648 42696 14700 42702
rect 14648 42638 14700 42644
rect 14556 41608 14608 41614
rect 14556 41550 14608 41556
rect 14568 41138 14596 41550
rect 14556 41132 14608 41138
rect 14556 41074 14608 41080
rect 14660 41002 14688 42638
rect 14752 41138 14780 42706
rect 15568 42696 15620 42702
rect 15568 42638 15620 42644
rect 15580 42362 15608 42638
rect 15844 42628 15896 42634
rect 15844 42570 15896 42576
rect 15752 42560 15804 42566
rect 15752 42502 15804 42508
rect 15568 42356 15620 42362
rect 15568 42298 15620 42304
rect 15292 42016 15344 42022
rect 15292 41958 15344 41964
rect 15304 41206 15332 41958
rect 15476 41540 15528 41546
rect 15476 41482 15528 41488
rect 15384 41472 15436 41478
rect 15384 41414 15436 41420
rect 15292 41200 15344 41206
rect 15292 41142 15344 41148
rect 14740 41132 14792 41138
rect 14740 41074 14792 41080
rect 14648 40996 14700 41002
rect 14648 40938 14700 40944
rect 14464 40520 14516 40526
rect 14464 40462 14516 40468
rect 14476 40118 14504 40462
rect 14648 40180 14700 40186
rect 14648 40122 14700 40128
rect 14464 40112 14516 40118
rect 14464 40054 14516 40060
rect 14188 39364 14240 39370
rect 14188 39306 14240 39312
rect 14200 39098 14228 39306
rect 14188 39092 14240 39098
rect 14188 39034 14240 39040
rect 14188 37800 14240 37806
rect 14188 37742 14240 37748
rect 14556 37800 14608 37806
rect 14556 37742 14608 37748
rect 14200 36922 14228 37742
rect 14188 36916 14240 36922
rect 14188 36858 14240 36864
rect 14568 36378 14596 37742
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14568 35698 14596 36314
rect 14556 35692 14608 35698
rect 14556 35634 14608 35640
rect 14016 35584 14136 35612
rect 13728 34672 13780 34678
rect 13728 34614 13780 34620
rect 13740 34202 13768 34614
rect 13820 34400 13872 34406
rect 13820 34342 13872 34348
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 13726 34096 13782 34105
rect 13726 34031 13782 34040
rect 13740 33998 13768 34031
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13832 33930 13860 34342
rect 13820 33924 13872 33930
rect 13820 33866 13872 33872
rect 13728 32904 13780 32910
rect 13728 32846 13780 32852
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 13636 32428 13688 32434
rect 13556 32388 13636 32416
rect 13636 32370 13688 32376
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13452 30932 13504 30938
rect 13452 30874 13504 30880
rect 13556 30870 13584 31758
rect 13636 31748 13688 31754
rect 13636 31690 13688 31696
rect 13544 30864 13596 30870
rect 13544 30806 13596 30812
rect 13648 30734 13676 31690
rect 13636 30728 13688 30734
rect 13636 30670 13688 30676
rect 13544 30592 13596 30598
rect 13740 30580 13768 32846
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 13820 31748 13872 31754
rect 13820 31690 13872 31696
rect 13832 31414 13860 31690
rect 13820 31408 13872 31414
rect 13820 31350 13872 31356
rect 13820 31204 13872 31210
rect 13820 31146 13872 31152
rect 13596 30552 13768 30580
rect 13544 30534 13596 30540
rect 13268 28960 13320 28966
rect 13174 28928 13230 28937
rect 13268 28902 13320 28908
rect 13174 28863 13230 28872
rect 13188 28558 13216 28863
rect 13280 28694 13308 28902
rect 13556 28762 13584 30534
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 13832 28694 13860 31146
rect 13924 30938 13952 32166
rect 13912 30932 13964 30938
rect 13912 30874 13964 30880
rect 13912 30660 13964 30666
rect 13912 30602 13964 30608
rect 13924 29306 13952 30602
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 13268 28688 13320 28694
rect 13268 28630 13320 28636
rect 13820 28688 13872 28694
rect 13820 28630 13872 28636
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 12716 28144 12768 28150
rect 12716 28086 12768 28092
rect 12438 27911 12494 27920
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 12820 27674 12848 27814
rect 12808 27668 12860 27674
rect 12808 27610 12860 27616
rect 12072 26920 12124 26926
rect 12072 26862 12124 26868
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 24818 11560 26726
rect 12084 26586 12112 26862
rect 13096 26586 13124 28494
rect 13464 28150 13492 28562
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13556 28150 13584 28426
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 13544 28144 13596 28150
rect 13544 28086 13596 28092
rect 13634 28112 13690 28121
rect 13464 27674 13492 28086
rect 13452 27668 13504 27674
rect 13452 27610 13504 27616
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11612 25968 11664 25974
rect 11612 25910 11664 25916
rect 11624 25226 11652 25910
rect 11808 25498 11836 26250
rect 12452 26042 12480 26386
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11624 24954 11652 25162
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11900 24818 11928 25638
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 12452 24274 12480 25978
rect 13464 25906 13492 27066
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13004 25498 13032 25842
rect 13360 25696 13412 25702
rect 13360 25638 13412 25644
rect 13372 25498 13400 25638
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13464 24954 13492 25842
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11532 23322 11560 23598
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11624 22642 11652 23054
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11624 22094 11652 22578
rect 11808 22438 11836 24142
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11900 22710 11928 24006
rect 12084 23866 12112 24142
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12452 23662 12480 24006
rect 12544 23866 12572 24006
rect 12636 23866 12664 24074
rect 12532 23860 12584 23866
rect 12532 23802 12584 23808
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12820 23662 12848 24210
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11624 22066 12020 22094
rect 11992 21486 12020 22066
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11440 20602 11468 21082
rect 11992 20942 12020 21422
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 11072 17746 11100 19722
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11532 18834 11560 19654
rect 11900 19514 11928 20266
rect 11992 19854 12020 20878
rect 12084 20534 12112 23530
rect 12912 23118 12940 24006
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13556 22710 13584 28086
rect 13634 28047 13636 28056
rect 13688 28047 13690 28056
rect 13636 28018 13688 28024
rect 13636 27872 13688 27878
rect 13636 27814 13688 27820
rect 13648 27402 13676 27814
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13636 27396 13688 27402
rect 13636 27338 13688 27344
rect 13648 25922 13676 27338
rect 13740 27130 13768 27474
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13648 25894 13768 25922
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13648 24750 13676 25094
rect 13740 24886 13768 25894
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13648 22778 13676 23598
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 12084 20058 12112 20470
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12084 19310 12112 19654
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17338 7144 17478
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 1584 15972 1636 15978
rect 1584 15914 1636 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 7024 15026 7052 16594
rect 7208 16574 7236 17546
rect 10796 17270 10824 17546
rect 11440 17270 11468 18022
rect 11716 17882 11744 18158
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7300 16658 7328 16934
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7116 16546 7236 16574
rect 7116 16046 7144 16546
rect 10796 16522 10824 17206
rect 11532 17202 11560 17682
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 12176 16574 12204 22374
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 13096 21622 13124 21830
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12268 20398 12296 20810
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19514 12480 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 13096 19446 13124 20334
rect 13556 20262 13584 21286
rect 13832 21146 13860 28358
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13832 20602 13860 21082
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18970 12480 19314
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12360 17746 12388 18022
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17270 12296 17478
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12084 16546 12204 16574
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16182 9536 16390
rect 9692 16250 9720 16458
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7024 14618 7052 14962
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14498 7144 15982
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15706 8340 15846
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8956 15502 8984 15982
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8404 15026 8432 15438
rect 9692 15434 9720 16186
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 10690 15736 10746 15745
rect 10690 15671 10692 15680
rect 10744 15671 10746 15680
rect 10692 15642 10744 15648
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8772 14618 8800 14894
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 7024 14470 7144 14498
rect 8944 14476 8996 14482
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 1584 12708 1636 12714
rect 1584 12650 1636 12656
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1596 2650 1624 12650
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 6932 9178 6960 13398
rect 7024 13394 7052 14470
rect 8944 14418 8996 14424
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7300 14074 7328 14282
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7208 13530 7236 13874
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 8956 13394 8984 14418
rect 9692 14346 9720 15370
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 7024 12918 7052 13330
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9232 12986 9260 13194
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 9968 12646 9996 13194
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12434 9996 12582
rect 10152 12434 10180 14962
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14618 10272 14758
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10690 14376 10746 14385
rect 10690 14311 10746 14320
rect 10704 14278 10732 14311
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 11256 13734 11284 15982
rect 11426 15464 11482 15473
rect 11426 15399 11428 15408
rect 11480 15399 11482 15408
rect 11428 15370 11480 15376
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14550 11836 14962
rect 11978 14920 12034 14929
rect 11978 14855 12034 14864
rect 11992 14618 12020 14855
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 13852 11468 14418
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11532 14074 11560 14214
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11440 13824 11560 13852
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 13530 11376 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11348 12850 11376 13126
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 9784 12406 9996 12434
rect 10060 12406 10180 12434
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 6932 7002 6960 7278
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6458 5764 6734
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6380 6458 6408 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 7300 6390 7328 6666
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5710 3832 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1872 4826 1900 5102
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2700 4554 2728 5306
rect 3252 5030 3280 5646
rect 4172 5370 4200 5646
rect 5460 5642 5488 6326
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 5920 5914 5948 6190
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6932 5778 6960 6190
rect 7300 5914 7328 6326
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 5460 5234 5488 5578
rect 6932 5370 6960 5714
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4690 3280 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 3068 4282 3096 4558
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3252 4146 3280 4626
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3602 3280 4082
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3618 4660 4014
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 4540 3590 4660 3618
rect 4540 3194 4568 3590
rect 5460 3534 5488 5170
rect 7300 4214 7328 5850
rect 7576 5642 7604 7142
rect 9784 6798 9812 12406
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 8220 6254 8248 6734
rect 9508 6458 9536 6734
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9600 6322 9628 6598
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8588 5914 8616 6190
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 9600 5846 9628 6258
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 9600 5302 9628 5782
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4622 8340 4966
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5552 3602 5580 4014
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3528 5500 3534
rect 5500 3476 5580 3482
rect 5448 3470 5580 3476
rect 5460 3454 5580 3470
rect 5552 3194 5580 3454
rect 6012 3194 6040 3878
rect 6196 3194 6224 4082
rect 7300 3466 7328 4150
rect 7668 4146 7696 4422
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7760 3738 7788 3946
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8036 3466 8064 4014
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3738 8248 3878
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6932 2990 6960 3334
rect 7668 3058 7696 3402
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2774 6960 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 6932 2746 7236 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 7208 2514 7236 2746
rect 8312 2514 8340 4558
rect 8496 2650 8524 4626
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4010 8984 4422
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 9324 3738 9352 4558
rect 9600 4162 9628 5238
rect 9692 4622 9720 5578
rect 9784 5574 9812 6734
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4214 9720 4558
rect 9508 4134 9628 4162
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9508 3126 9536 4134
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3738 9628 4014
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9600 3058 9628 3538
rect 9784 3534 9812 5510
rect 10060 5370 10088 12406
rect 11440 11762 11468 13126
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11082 11468 11698
rect 11532 11121 11560 13824
rect 11624 12986 11652 14214
rect 11808 13394 11836 14486
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11900 13274 11928 14214
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11808 13246 11928 13274
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12646 11652 12786
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 11778 11652 12106
rect 11716 11898 11744 12922
rect 11808 12102 11836 13246
rect 11992 12850 12020 13874
rect 12084 12918 12112 16546
rect 13464 16250 13492 19994
rect 13556 19446 13584 20198
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 14016 18154 14044 35584
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 14108 32978 14136 33254
rect 14096 32972 14148 32978
rect 14096 32914 14148 32920
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 14108 31210 14136 31962
rect 14200 31754 14228 34546
rect 14280 34400 14332 34406
rect 14280 34342 14332 34348
rect 14292 33386 14320 34342
rect 14568 34202 14596 34682
rect 14660 34202 14688 40122
rect 15396 39982 15424 41414
rect 15384 39976 15436 39982
rect 15384 39918 15436 39924
rect 15396 39506 15424 39918
rect 15384 39500 15436 39506
rect 15384 39442 15436 39448
rect 15108 39432 15160 39438
rect 15108 39374 15160 39380
rect 15120 39098 15148 39374
rect 15108 39092 15160 39098
rect 15108 39034 15160 39040
rect 15396 38418 15424 39442
rect 15384 38412 15436 38418
rect 15384 38354 15436 38360
rect 15396 38026 15424 38354
rect 15212 38010 15424 38026
rect 15200 38004 15424 38010
rect 15252 37998 15424 38004
rect 15200 37946 15252 37952
rect 15488 37942 15516 41482
rect 15764 41274 15792 42502
rect 15856 42090 15884 42570
rect 15844 42084 15896 42090
rect 15844 42026 15896 42032
rect 15752 41268 15804 41274
rect 15752 41210 15804 41216
rect 15948 41154 15976 45494
rect 16212 45280 16264 45286
rect 16212 45222 16264 45228
rect 16224 44946 16252 45222
rect 16316 45082 16344 45494
rect 16304 45076 16356 45082
rect 16304 45018 16356 45024
rect 16212 44940 16264 44946
rect 16212 44882 16264 44888
rect 16500 43858 16528 45494
rect 22020 45490 22048 45526
rect 24136 45490 24164 45970
rect 33152 45966 33180 46838
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 41892 45966 41920 47681
rect 27896 45960 27948 45966
rect 27896 45902 27948 45908
rect 33140 45960 33192 45966
rect 33140 45902 33192 45908
rect 41880 45960 41932 45966
rect 41880 45902 41932 45908
rect 24952 45824 25004 45830
rect 24952 45766 25004 45772
rect 27528 45824 27580 45830
rect 27528 45766 27580 45772
rect 16856 45484 16908 45490
rect 16856 45426 16908 45432
rect 18420 45484 18472 45490
rect 18420 45426 18472 45432
rect 22008 45484 22060 45490
rect 22008 45426 22060 45432
rect 23388 45484 23440 45490
rect 23388 45426 23440 45432
rect 23940 45484 23992 45490
rect 23940 45426 23992 45432
rect 24124 45484 24176 45490
rect 24124 45426 24176 45432
rect 16580 45348 16632 45354
rect 16580 45290 16632 45296
rect 16592 44792 16620 45290
rect 16672 44804 16724 44810
rect 16592 44764 16672 44792
rect 16672 44746 16724 44752
rect 16684 44402 16712 44746
rect 16868 44742 16896 45426
rect 17316 45416 17368 45422
rect 17316 45358 17368 45364
rect 17040 45280 17092 45286
rect 17040 45222 17092 45228
rect 16856 44736 16908 44742
rect 16856 44678 16908 44684
rect 16672 44396 16724 44402
rect 16672 44338 16724 44344
rect 16672 44192 16724 44198
rect 16672 44134 16724 44140
rect 16488 43852 16540 43858
rect 16488 43794 16540 43800
rect 16684 43790 16712 44134
rect 16672 43784 16724 43790
rect 16672 43726 16724 43732
rect 16672 43240 16724 43246
rect 16672 43182 16724 43188
rect 16684 42906 16712 43182
rect 16672 42900 16724 42906
rect 16672 42842 16724 42848
rect 16488 42628 16540 42634
rect 16488 42570 16540 42576
rect 16500 41614 16528 42570
rect 16488 41608 16540 41614
rect 16488 41550 16540 41556
rect 16028 41540 16080 41546
rect 16028 41482 16080 41488
rect 16040 41274 16068 41482
rect 16028 41268 16080 41274
rect 16028 41210 16080 41216
rect 15672 41126 15976 41154
rect 15476 37936 15528 37942
rect 15476 37878 15528 37884
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 15212 37738 15240 37810
rect 15200 37732 15252 37738
rect 15200 37674 15252 37680
rect 15212 36106 15240 37674
rect 15200 36100 15252 36106
rect 15200 36042 15252 36048
rect 14740 35692 14792 35698
rect 14740 35634 14792 35640
rect 14556 34196 14608 34202
rect 14556 34138 14608 34144
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 14292 33114 14320 33322
rect 14280 33108 14332 33114
rect 14280 33050 14332 33056
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14292 31793 14320 31826
rect 14384 31822 14412 33934
rect 14476 33522 14504 33934
rect 14660 33674 14688 34138
rect 14568 33658 14688 33674
rect 14556 33652 14688 33658
rect 14608 33646 14688 33652
rect 14556 33594 14608 33600
rect 14648 33584 14700 33590
rect 14648 33526 14700 33532
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14476 32910 14504 33458
rect 14660 33114 14688 33526
rect 14648 33108 14700 33114
rect 14648 33050 14700 33056
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 14752 31890 14780 35634
rect 15016 33856 15068 33862
rect 15068 33816 15148 33844
rect 15016 33798 15068 33804
rect 14924 33516 14976 33522
rect 15120 33504 15148 33816
rect 14976 33476 15148 33504
rect 14924 33458 14976 33464
rect 15120 32978 15148 33476
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15212 33046 15240 33390
rect 15200 33040 15252 33046
rect 15200 32982 15252 32988
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15108 32836 15160 32842
rect 15108 32778 15160 32784
rect 15120 32570 15148 32778
rect 15212 32570 15240 32846
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15304 32502 15332 33390
rect 15488 32910 15516 37878
rect 15672 37874 15700 41126
rect 15844 41064 15896 41070
rect 15844 41006 15896 41012
rect 15856 38010 15884 41006
rect 16120 40724 16172 40730
rect 16120 40666 16172 40672
rect 15936 40588 15988 40594
rect 15936 40530 15988 40536
rect 15948 40050 15976 40530
rect 16028 40384 16080 40390
rect 16028 40326 16080 40332
rect 15936 40044 15988 40050
rect 15936 39986 15988 39992
rect 16040 39982 16068 40326
rect 16132 40050 16160 40666
rect 16120 40044 16172 40050
rect 16120 39986 16172 39992
rect 16212 40044 16264 40050
rect 16212 39986 16264 39992
rect 16028 39976 16080 39982
rect 16028 39918 16080 39924
rect 16224 39098 16252 39986
rect 16212 39092 16264 39098
rect 16212 39034 16264 39040
rect 16396 38956 16448 38962
rect 16396 38898 16448 38904
rect 15936 38276 15988 38282
rect 15936 38218 15988 38224
rect 15948 38010 15976 38218
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15936 38004 15988 38010
rect 15936 37946 15988 37952
rect 15660 37868 15712 37874
rect 15660 37810 15712 37816
rect 15856 37262 15884 37946
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 16040 36378 16068 36722
rect 16028 36372 16080 36378
rect 16028 36314 16080 36320
rect 15660 36100 15712 36106
rect 15660 36042 15712 36048
rect 15672 35630 15700 36042
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15752 34400 15804 34406
rect 15752 34342 15804 34348
rect 15764 34202 15792 34342
rect 16040 34202 16068 36314
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 15752 34196 15804 34202
rect 15752 34138 15804 34144
rect 16028 34196 16080 34202
rect 16028 34138 16080 34144
rect 15672 34048 15700 34138
rect 15672 34020 15976 34048
rect 15752 33924 15804 33930
rect 15752 33866 15804 33872
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 14832 32020 14884 32026
rect 14832 31962 14884 31968
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14372 31816 14424 31822
rect 14278 31784 14334 31793
rect 14188 31748 14240 31754
rect 14372 31758 14424 31764
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 14278 31719 14334 31728
rect 14188 31690 14240 31696
rect 14096 31204 14148 31210
rect 14096 31146 14148 31152
rect 14096 30660 14148 30666
rect 14096 30602 14148 30608
rect 14108 30190 14136 30602
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 14384 28994 14412 31758
rect 14660 31482 14688 31758
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14844 31346 14872 31962
rect 15488 31793 15516 32846
rect 15764 32434 15792 33866
rect 15948 33318 15976 34020
rect 16132 33998 16160 34342
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16120 33992 16172 33998
rect 16120 33934 16172 33940
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16040 33658 16068 33934
rect 16028 33652 16080 33658
rect 16028 33594 16080 33600
rect 16224 33522 16252 33934
rect 16408 33522 16436 38898
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16592 37874 16620 38694
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16684 35834 16712 36518
rect 16764 36236 16816 36242
rect 16764 36178 16816 36184
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 16672 34196 16724 34202
rect 16672 34138 16724 34144
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 16396 33516 16448 33522
rect 16396 33458 16448 33464
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 15672 32026 15700 32370
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15474 31784 15530 31793
rect 15856 31754 15884 33254
rect 15948 32570 15976 33254
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 16224 32434 16252 32846
rect 16316 32570 16344 33390
rect 16304 32564 16356 32570
rect 16304 32506 16356 32512
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 15474 31719 15530 31728
rect 15764 31726 15884 31754
rect 14740 31340 14792 31346
rect 14292 28966 14412 28994
rect 14660 31300 14740 31328
rect 14292 28150 14320 28966
rect 14464 28960 14516 28966
rect 14464 28902 14516 28908
rect 14476 28558 14504 28902
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14384 28014 14412 28358
rect 14476 28014 14504 28494
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14108 26994 14136 27814
rect 14292 27674 14320 27814
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 14556 27396 14608 27402
rect 14556 27338 14608 27344
rect 14568 27130 14596 27338
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14108 23050 14136 24142
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14188 21548 14240 21554
rect 14292 21536 14320 24278
rect 14660 23662 14688 31300
rect 14740 31282 14792 31288
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 15488 31278 15516 31719
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 14740 31136 14792 31142
rect 14740 31078 14792 31084
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 14752 27062 14780 31078
rect 15488 30938 15516 31078
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15292 30728 15344 30734
rect 14830 30696 14886 30705
rect 15292 30670 15344 30676
rect 14830 30631 14832 30640
rect 14884 30631 14886 30640
rect 14832 30602 14884 30608
rect 15304 30326 15332 30670
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14936 29238 14964 29582
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15212 29306 15240 29446
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15304 29238 15332 30262
rect 15580 29646 15608 31282
rect 15660 31136 15712 31142
rect 15660 31078 15712 31084
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14844 28150 14872 28358
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14936 27962 14964 29174
rect 15396 29170 15424 29446
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15028 28014 15056 29106
rect 15212 28762 15240 29106
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15396 28014 15424 29106
rect 15672 29102 15700 31078
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 14844 27934 14964 27962
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 14844 25226 14872 27934
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14936 26994 14964 27814
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14844 24954 14872 25162
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14936 24818 14964 25298
rect 15212 25294 15240 25638
rect 15304 25498 15332 26250
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15120 24410 15148 24754
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15212 24206 15240 25230
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 14648 23656 14700 23662
rect 15304 23633 15332 25434
rect 14648 23598 14700 23604
rect 15290 23624 15346 23633
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14476 21690 14504 22578
rect 14660 22094 14688 23598
rect 15290 23559 15346 23568
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14844 22234 14872 22986
rect 14936 22778 14964 22986
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 15304 22556 15332 23559
rect 15672 22778 15700 29038
rect 15764 28082 15792 31726
rect 16224 31346 16252 32370
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 15856 30394 15884 30670
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 16224 30054 16252 30534
rect 16304 30184 16356 30190
rect 16304 30126 16356 30132
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16316 29646 16344 30126
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16316 29306 16344 29582
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16408 28626 16436 33458
rect 16500 33114 16528 33458
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16684 32366 16712 34138
rect 16776 33114 16804 36178
rect 16868 34746 16896 44678
rect 17052 44538 17080 45222
rect 17328 44538 17356 45358
rect 18236 45280 18288 45286
rect 18236 45222 18288 45228
rect 18248 45082 18276 45222
rect 18236 45076 18288 45082
rect 18236 45018 18288 45024
rect 17868 44804 17920 44810
rect 17920 44764 18092 44792
rect 17868 44746 17920 44752
rect 17040 44532 17092 44538
rect 17040 44474 17092 44480
rect 17316 44532 17368 44538
rect 17316 44474 17368 44480
rect 17500 44396 17552 44402
rect 17500 44338 17552 44344
rect 17132 44328 17184 44334
rect 17132 44270 17184 44276
rect 17316 44328 17368 44334
rect 17316 44270 17368 44276
rect 17144 42566 17172 44270
rect 17328 43722 17356 44270
rect 17316 43716 17368 43722
rect 17316 43658 17368 43664
rect 17316 43104 17368 43110
rect 17316 43046 17368 43052
rect 17328 42906 17356 43046
rect 17316 42900 17368 42906
rect 17316 42842 17368 42848
rect 17512 42634 17540 44338
rect 18064 44266 18092 44764
rect 18052 44260 18104 44266
rect 18052 44202 18104 44208
rect 18064 42702 18092 44202
rect 18432 43994 18460 45426
rect 22376 45280 22428 45286
rect 22376 45222 22428 45228
rect 22192 44940 22244 44946
rect 22192 44882 22244 44888
rect 21180 44872 21232 44878
rect 21180 44814 21232 44820
rect 20628 44804 20680 44810
rect 20628 44746 20680 44752
rect 19064 44736 19116 44742
rect 19064 44678 19116 44684
rect 18880 44396 18932 44402
rect 18880 44338 18932 44344
rect 18892 43994 18920 44338
rect 18420 43988 18472 43994
rect 18420 43930 18472 43936
rect 18880 43988 18932 43994
rect 18880 43930 18932 43936
rect 18880 43852 18932 43858
rect 18880 43794 18932 43800
rect 18420 43648 18472 43654
rect 18420 43590 18472 43596
rect 18052 42696 18104 42702
rect 18052 42638 18104 42644
rect 17500 42628 17552 42634
rect 17500 42570 17552 42576
rect 17132 42560 17184 42566
rect 17132 42502 17184 42508
rect 17144 42362 17172 42502
rect 17132 42356 17184 42362
rect 17132 42298 17184 42304
rect 17316 42152 17368 42158
rect 17316 42094 17368 42100
rect 17328 41818 17356 42094
rect 17316 41812 17368 41818
rect 17316 41754 17368 41760
rect 17316 41200 17368 41206
rect 17316 41142 17368 41148
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 16960 39914 16988 40054
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 16948 39908 17000 39914
rect 16948 39850 17000 39856
rect 17144 39642 17172 39986
rect 17132 39636 17184 39642
rect 17132 39578 17184 39584
rect 17040 39296 17092 39302
rect 17040 39238 17092 39244
rect 17052 38962 17080 39238
rect 17040 38956 17092 38962
rect 17040 38898 17092 38904
rect 17052 36922 17080 38898
rect 17328 38350 17356 41142
rect 17512 40594 17540 42570
rect 17592 42560 17644 42566
rect 17592 42502 17644 42508
rect 17604 42226 17632 42502
rect 18064 42294 18092 42638
rect 18052 42288 18104 42294
rect 18052 42230 18104 42236
rect 17592 42220 17644 42226
rect 17592 42162 17644 42168
rect 18328 41676 18380 41682
rect 18328 41618 18380 41624
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 17500 40588 17552 40594
rect 17500 40530 17552 40536
rect 17684 40384 17736 40390
rect 17684 40326 17736 40332
rect 17696 40186 17724 40326
rect 17684 40180 17736 40186
rect 17684 40122 17736 40128
rect 17592 39840 17644 39846
rect 17592 39782 17644 39788
rect 17604 39098 17632 39782
rect 17684 39432 17736 39438
rect 17684 39374 17736 39380
rect 17592 39092 17644 39098
rect 17592 39034 17644 39040
rect 17408 38888 17460 38894
rect 17408 38830 17460 38836
rect 17420 38418 17448 38830
rect 17592 38820 17644 38826
rect 17592 38762 17644 38768
rect 17408 38412 17460 38418
rect 17408 38354 17460 38360
rect 17316 38344 17368 38350
rect 17316 38286 17368 38292
rect 17604 37670 17632 38762
rect 17696 38554 17724 39374
rect 17880 39030 17908 40666
rect 17868 39024 17920 39030
rect 17868 38966 17920 38972
rect 17684 38548 17736 38554
rect 17684 38490 17736 38496
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17592 37664 17644 37670
rect 17592 37606 17644 37612
rect 17604 37108 17632 37606
rect 17696 37466 17724 37810
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 17788 37262 17816 38150
rect 17972 38010 18000 41414
rect 18340 41206 18368 41618
rect 18328 41200 18380 41206
rect 18328 41142 18380 41148
rect 18328 39840 18380 39846
rect 18328 39782 18380 39788
rect 18340 39574 18368 39782
rect 18328 39568 18380 39574
rect 18328 39510 18380 39516
rect 18236 38344 18288 38350
rect 18236 38286 18288 38292
rect 18144 38208 18196 38214
rect 18144 38150 18196 38156
rect 17960 38004 18012 38010
rect 17960 37946 18012 37952
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17604 37080 17816 37108
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 17788 36242 17816 37080
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 17776 36236 17828 36242
rect 17776 36178 17828 36184
rect 16960 35630 16988 36178
rect 17788 35630 17816 36178
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 17960 36100 18012 36106
rect 17960 36042 18012 36048
rect 17868 36032 17920 36038
rect 17868 35974 17920 35980
rect 17880 35834 17908 35974
rect 17868 35828 17920 35834
rect 17868 35770 17920 35776
rect 17972 35766 18000 36042
rect 17960 35760 18012 35766
rect 17960 35702 18012 35708
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 17776 35624 17828 35630
rect 17776 35566 17828 35572
rect 18064 35290 18092 36110
rect 18052 35284 18104 35290
rect 18052 35226 18104 35232
rect 18156 35154 18184 38150
rect 18248 37126 18276 38286
rect 18432 37618 18460 43590
rect 18788 42696 18840 42702
rect 18788 42638 18840 42644
rect 18512 42560 18564 42566
rect 18512 42502 18564 42508
rect 18696 42560 18748 42566
rect 18696 42502 18748 42508
rect 18524 41818 18552 42502
rect 18708 42226 18736 42502
rect 18696 42220 18748 42226
rect 18696 42162 18748 42168
rect 18800 41818 18828 42638
rect 18512 41812 18564 41818
rect 18512 41754 18564 41760
rect 18788 41812 18840 41818
rect 18788 41754 18840 41760
rect 18788 41608 18840 41614
rect 18788 41550 18840 41556
rect 18800 41274 18828 41550
rect 18788 41268 18840 41274
rect 18788 41210 18840 41216
rect 18892 41154 18920 43794
rect 19076 43654 19104 44678
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19616 44192 19668 44198
rect 19616 44134 19668 44140
rect 19628 43790 19656 44134
rect 19616 43784 19668 43790
rect 19616 43726 19668 43732
rect 20444 43716 20496 43722
rect 20444 43658 20496 43664
rect 19064 43648 19116 43654
rect 19064 43590 19116 43596
rect 20076 43648 20128 43654
rect 20076 43590 20128 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19156 43104 19208 43110
rect 19156 43046 19208 43052
rect 19168 42158 19196 43046
rect 19340 42696 19392 42702
rect 19340 42638 19392 42644
rect 19156 42152 19208 42158
rect 19156 42094 19208 42100
rect 18972 42016 19024 42022
rect 18972 41958 19024 41964
rect 18984 41478 19012 41958
rect 18972 41472 19024 41478
rect 18972 41414 19024 41420
rect 18708 41138 18920 41154
rect 18696 41132 18920 41138
rect 18748 41126 18920 41132
rect 18696 41074 18748 41080
rect 18708 40730 18736 41074
rect 18696 40724 18748 40730
rect 18696 40666 18748 40672
rect 19168 40594 19196 42094
rect 19352 41818 19380 42638
rect 19984 42560 20036 42566
rect 19984 42502 20036 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19800 42356 19852 42362
rect 19800 42298 19852 42304
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19812 41750 19840 42298
rect 19996 42158 20024 42502
rect 19984 42152 20036 42158
rect 19984 42094 20036 42100
rect 20088 41818 20116 43590
rect 20076 41812 20128 41818
rect 20076 41754 20128 41760
rect 19800 41744 19852 41750
rect 19800 41686 19852 41692
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 20456 41206 20484 43658
rect 20640 42158 20668 44746
rect 21192 44334 21220 44814
rect 21180 44328 21232 44334
rect 21180 44270 21232 44276
rect 20812 43308 20864 43314
rect 20812 43250 20864 43256
rect 20628 42152 20680 42158
rect 20628 42094 20680 42100
rect 20536 42016 20588 42022
rect 20536 41958 20588 41964
rect 20548 41818 20576 41958
rect 20536 41812 20588 41818
rect 20536 41754 20588 41760
rect 20444 41200 20496 41206
rect 20444 41142 20496 41148
rect 19156 40588 19208 40594
rect 19156 40530 19208 40536
rect 20168 40520 20220 40526
rect 20168 40462 20220 40468
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 18788 39840 18840 39846
rect 18788 39782 18840 39788
rect 18800 39030 18828 39782
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19156 39296 19208 39302
rect 19156 39238 19208 39244
rect 18788 39024 18840 39030
rect 18788 38966 18840 38972
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 18616 38554 18644 38898
rect 18604 38548 18656 38554
rect 18604 38490 18656 38496
rect 19168 38418 19196 39238
rect 19444 38962 19472 39374
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19996 39098 20024 39306
rect 20180 39098 20208 40462
rect 20352 39568 20404 39574
rect 20352 39510 20404 39516
rect 20260 39296 20312 39302
rect 20260 39238 20312 39244
rect 20272 39098 20300 39238
rect 20364 39098 20392 39510
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20260 39092 20312 39098
rect 20260 39034 20312 39040
rect 20352 39092 20404 39098
rect 20352 39034 20404 39040
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 20456 38842 20484 41142
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20548 39794 20576 40870
rect 20640 40118 20668 42094
rect 20720 41608 20772 41614
rect 20720 41550 20772 41556
rect 20628 40112 20680 40118
rect 20628 40054 20680 40060
rect 20640 39930 20668 40054
rect 20732 40050 20760 41550
rect 20720 40044 20772 40050
rect 20720 39986 20772 39992
rect 20640 39902 20760 39930
rect 20548 39766 20668 39794
rect 20364 38826 20484 38842
rect 20352 38820 20484 38826
rect 20404 38814 20484 38820
rect 20352 38762 20404 38768
rect 19156 38412 19208 38418
rect 19156 38354 19208 38360
rect 18788 38344 18840 38350
rect 18788 38286 18840 38292
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 18340 37590 18460 37618
rect 18236 37120 18288 37126
rect 18236 37062 18288 37068
rect 18144 35148 18196 35154
rect 18144 35090 18196 35096
rect 18236 35080 18288 35086
rect 18236 35022 18288 35028
rect 18248 34746 18276 35022
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 18052 34740 18104 34746
rect 18052 34682 18104 34688
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 16856 33856 16908 33862
rect 16856 33798 16908 33804
rect 16868 33658 16896 33798
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16776 31754 16804 33050
rect 17052 32570 17080 34342
rect 17132 33992 17184 33998
rect 17132 33934 17184 33940
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17144 33697 17172 33934
rect 17224 33924 17276 33930
rect 17224 33866 17276 33872
rect 17130 33688 17186 33697
rect 17236 33658 17264 33866
rect 17130 33623 17186 33632
rect 17224 33652 17276 33658
rect 17224 33594 17276 33600
rect 17328 33590 17356 33934
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 17684 33924 17736 33930
rect 17684 33866 17736 33872
rect 17316 33584 17368 33590
rect 17316 33526 17368 33532
rect 17132 32836 17184 32842
rect 17132 32778 17184 32784
rect 17040 32564 17092 32570
rect 17040 32506 17092 32512
rect 17052 32434 17080 32506
rect 17144 32434 17172 32778
rect 17408 32768 17460 32774
rect 17408 32710 17460 32716
rect 17420 32570 17448 32710
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 16684 31726 16804 31754
rect 16488 30932 16540 30938
rect 16488 30874 16540 30880
rect 16500 30734 16528 30874
rect 16684 30802 16712 31726
rect 16672 30796 16724 30802
rect 16672 30738 16724 30744
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16488 30592 16540 30598
rect 16540 30540 16620 30546
rect 16488 30534 16620 30540
rect 16500 30518 16620 30534
rect 16592 30258 16620 30518
rect 16684 30394 16712 30602
rect 16672 30388 16724 30394
rect 16672 30330 16724 30336
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16592 28937 16620 30194
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16578 28928 16634 28937
rect 16578 28863 16634 28872
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15856 24410 15884 24754
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15384 22568 15436 22574
rect 15212 22528 15384 22556
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14660 22066 14780 22094
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14660 21690 14688 21966
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14240 21508 14320 21536
rect 14188 21490 14240 21496
rect 14200 20942 14228 21490
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14108 19990 14136 20878
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20398 14504 20742
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14476 19514 14504 20334
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19514 14596 19790
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14108 18970 14136 19314
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16658 14320 16934
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 16250 14136 16526
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12176 15162 12204 15438
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12176 14618 12204 14962
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11992 12374 12020 12786
rect 12268 12442 12296 14962
rect 12360 13530 12388 15438
rect 13096 15162 13124 15438
rect 13188 15162 13216 15506
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13464 15094 13492 16186
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15638 13584 15846
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12544 14618 12572 14962
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13530 12572 13874
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11624 11750 11744 11778
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11518 11112 11574 11121
rect 11428 11076 11480 11082
rect 11518 11047 11574 11056
rect 11428 11018 11480 11024
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11058 10296 11114 10305
rect 11058 10231 11060 10240
rect 11112 10231 11114 10240
rect 11060 10202 11112 10208
rect 11256 9518 11284 10406
rect 11532 10130 11560 11047
rect 11624 10674 11652 11630
rect 11716 11558 11744 11750
rect 11704 11552 11756 11558
rect 11808 11529 11836 12038
rect 11900 11750 11928 12106
rect 12360 12084 12388 12786
rect 12544 12646 12572 12786
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12452 12374 12480 12582
rect 12544 12481 12572 12582
rect 12530 12472 12586 12481
rect 12530 12407 12586 12416
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12532 12232 12584 12238
rect 12636 12220 12664 13126
rect 12584 12192 12664 12220
rect 12532 12174 12584 12180
rect 12532 12096 12584 12102
rect 12360 12064 12532 12084
rect 12584 12064 12586 12073
rect 12360 12056 12530 12064
rect 12530 11999 12586 12008
rect 12164 11756 12216 11762
rect 11900 11722 12164 11750
rect 11704 11494 11756 11500
rect 11794 11520 11850 11529
rect 11716 11370 11744 11494
rect 11794 11455 11850 11464
rect 11716 11342 11836 11370
rect 11808 10674 11836 11342
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 7750 11284 9454
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11440 8362 11468 9386
rect 11532 9042 11560 9522
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11624 7954 11652 10610
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 9586 11744 10542
rect 11808 10470 11836 10610
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11900 10282 11928 11722
rect 12164 11698 12216 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11808 10254 11928 10282
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11808 9450 11836 10254
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11808 8974 11836 9386
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11716 8634 11744 8842
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11716 8090 11744 8570
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6798 11376 7142
rect 11624 7002 11652 7890
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7002 11744 7346
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11808 6662 11836 7754
rect 11900 6866 11928 9998
rect 11992 9722 12020 9998
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 9382 12020 9522
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 7818 12020 9114
rect 12084 8090 12112 11630
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12176 10198 12204 11290
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10810 12572 10950
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12268 10266 12296 10406
rect 12360 10266 12388 10542
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12544 9926 12572 10746
rect 12636 10606 12664 12192
rect 12728 11898 12756 13262
rect 12912 13258 12940 14758
rect 13188 14362 13216 14962
rect 13188 14334 13308 14362
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 13326 13124 13874
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12238 12940 13194
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12986 13124 13126
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12728 10810 12756 11834
rect 12820 11762 12848 12038
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12912 11642 12940 12038
rect 12820 11614 12940 11642
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 10266 12664 10542
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12268 9058 12296 9862
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9489 12388 9522
rect 12346 9480 12402 9489
rect 12346 9415 12402 9424
rect 12176 9030 12296 9058
rect 12176 8430 12204 9030
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8430 12296 8910
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10060 4826 10088 5306
rect 10336 5234 10364 6054
rect 11992 5914 12020 7754
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12084 7410 12112 7482
rect 12268 7410 12296 7686
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12084 6780 12112 7346
rect 12164 6792 12216 6798
rect 12084 6752 12164 6780
rect 12164 6734 12216 6740
rect 12176 6254 12204 6734
rect 12360 6730 12388 9415
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 6746 12480 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 7886 12572 8434
rect 12636 8022 12664 10202
rect 12820 9926 12848 11614
rect 13004 11014 13032 12650
rect 13096 12442 13124 12786
rect 13188 12442 13216 14214
rect 13280 13841 13308 14334
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 14006 13400 14214
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13266 13832 13322 13841
rect 13266 13767 13322 13776
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13096 11626 13124 12378
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 13096 10130 13124 10542
rect 13280 10441 13308 13767
rect 13372 12986 13400 13942
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13372 12434 13400 12786
rect 13372 12406 13492 12434
rect 13464 12102 13492 12406
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13372 11150 13400 12038
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13266 10432 13322 10441
rect 13266 10367 13322 10376
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12728 9625 12756 9862
rect 12714 9616 12770 9625
rect 12820 9586 12848 9862
rect 12714 9551 12770 9560
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 12912 9518 12940 9998
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 9512 12952 9518
rect 13004 9489 13032 9522
rect 12900 9454 12952 9460
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13004 9110 13032 9415
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13096 8838 13124 10066
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13280 8090 13308 10367
rect 13372 9586 13400 10610
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 9178 13400 9522
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12544 7546 12572 7822
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12728 6934 12756 7822
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12348 6724 12400 6730
rect 12452 6718 12572 6746
rect 12348 6666 12400 6672
rect 12256 6656 12308 6662
rect 12360 6633 12388 6666
rect 12256 6598 12308 6604
rect 12346 6624 12402 6633
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12268 5846 12296 6598
rect 12346 6559 12402 6568
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 10416 5704 10468 5710
rect 12544 5681 12572 6718
rect 10416 5646 10468 5652
rect 12530 5672 12586 5681
rect 10428 5370 10456 5646
rect 10968 5636 11020 5642
rect 13096 5642 13124 7414
rect 13188 7206 13216 7754
rect 13280 7546 13308 7890
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6866 13216 7142
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13280 6390 13308 7482
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13372 6458 13400 7210
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13464 6186 13492 12038
rect 13556 10470 13584 15574
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13648 14550 13676 15370
rect 13832 15094 13860 15438
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13832 14618 13860 14826
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 13326 13676 14486
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13832 13870 13860 13942
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 12646 13768 13194
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 12209 13768 12310
rect 13726 12200 13782 12209
rect 13726 12135 13782 12144
rect 13924 11898 13952 16050
rect 14278 15872 14334 15881
rect 14278 15807 14334 15816
rect 14292 15706 14320 15807
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 14016 13870 14044 15370
rect 14476 15162 14504 16594
rect 14752 16182 14780 22066
rect 15212 21486 15240 22528
rect 15384 22510 15436 22516
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15764 21690 15792 21898
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15120 19990 15148 21422
rect 15212 20398 15240 21422
rect 15948 20602 15976 28494
rect 16040 28150 16068 28562
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16040 27674 16068 28086
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 16684 27538 16712 29038
rect 17144 28558 17172 32370
rect 17236 32230 17264 32506
rect 17604 32298 17632 33866
rect 17696 33386 17724 33866
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17684 33380 17736 33386
rect 17684 33322 17736 33328
rect 17696 33114 17724 33322
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17592 32292 17644 32298
rect 17592 32234 17644 32240
rect 17224 32224 17276 32230
rect 17224 32166 17276 32172
rect 17788 32026 17816 33458
rect 17880 32910 17908 34478
rect 18064 33998 18092 34682
rect 18340 33998 18368 37590
rect 18800 37466 18828 38286
rect 19260 38010 19288 38286
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 20456 37466 20484 38814
rect 18788 37460 18840 37466
rect 18788 37402 18840 37408
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 18420 36712 18472 36718
rect 18420 36654 18472 36660
rect 18432 35154 18460 36654
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 18432 34542 18460 35090
rect 18420 34536 18472 34542
rect 18420 34478 18472 34484
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18064 33658 18092 33934
rect 18144 33856 18196 33862
rect 18144 33798 18196 33804
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 18156 33522 18184 33798
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 17880 32570 17908 32846
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 17788 31482 17816 31962
rect 18064 31929 18092 31962
rect 18156 31958 18184 33458
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18248 32570 18276 32710
rect 18236 32564 18288 32570
rect 18236 32506 18288 32512
rect 18432 32434 18460 33050
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18144 31952 18196 31958
rect 18050 31920 18106 31929
rect 18144 31894 18196 31900
rect 18050 31855 18106 31864
rect 18236 31884 18288 31890
rect 18236 31826 18288 31832
rect 17776 31476 17828 31482
rect 17776 31418 17828 31424
rect 18248 30938 18276 31826
rect 18340 31346 18368 32370
rect 18432 31822 18460 32370
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18236 30932 18288 30938
rect 18156 30892 18236 30920
rect 17684 30388 17736 30394
rect 17684 30330 17736 30336
rect 17696 29102 17724 30330
rect 18156 30326 18184 30892
rect 18236 30874 18288 30880
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 18248 29238 18276 30602
rect 18236 29232 18288 29238
rect 18236 29174 18288 29180
rect 17684 29096 17736 29102
rect 17684 29038 17736 29044
rect 17696 28558 17724 29038
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17684 28552 17736 28558
rect 17684 28494 17736 28500
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 28218 17632 28358
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17132 28008 17184 28014
rect 17132 27950 17184 27956
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16316 26382 16344 27270
rect 17144 26450 17172 27950
rect 18144 27396 18196 27402
rect 18144 27338 18196 27344
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17972 26568 18000 26726
rect 18052 26580 18104 26586
rect 17972 26540 18052 26568
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 16132 25498 16160 25638
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16224 24954 16252 25774
rect 16684 25498 16712 26318
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 17052 26042 17080 26250
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16776 24954 16804 25842
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17052 24954 17080 25434
rect 17144 25362 17172 26386
rect 17972 25770 18000 26540
rect 18052 26522 18104 26528
rect 18156 26382 18184 27338
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 17960 25764 18012 25770
rect 17960 25706 18012 25712
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 18156 25242 18184 26318
rect 18340 25498 18368 31282
rect 18432 26586 18460 31758
rect 18524 29646 18552 37198
rect 19260 36922 19288 37198
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 20076 36848 20128 36854
rect 20076 36790 20128 36796
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19444 35834 19472 36110
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19156 35488 19208 35494
rect 19156 35430 19208 35436
rect 19168 35290 19196 35430
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19444 34746 19472 35022
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34746 20024 34886
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 19616 34400 19668 34406
rect 19616 34342 19668 34348
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 18788 33312 18840 33318
rect 18788 33254 18840 33260
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18800 32434 18828 33254
rect 18892 32910 18920 33254
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 18972 32768 19024 32774
rect 18972 32710 19024 32716
rect 18984 32570 19012 32710
rect 19076 32570 19104 32778
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 19168 31890 19196 33390
rect 19260 32978 19288 33934
rect 19628 33930 19656 34342
rect 19616 33924 19668 33930
rect 19616 33866 19668 33872
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20088 33658 20116 36790
rect 20352 36780 20404 36786
rect 20352 36722 20404 36728
rect 20364 36360 20392 36722
rect 20456 36718 20484 37402
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20444 36372 20496 36378
rect 20364 36332 20444 36360
rect 20364 35834 20392 36332
rect 20444 36314 20496 36320
rect 20352 35828 20404 35834
rect 20352 35770 20404 35776
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20456 34746 20484 35770
rect 20444 34740 20496 34746
rect 20444 34682 20496 34688
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20272 34202 20300 34546
rect 20260 34196 20312 34202
rect 20260 34138 20312 34144
rect 20076 33652 20128 33658
rect 20076 33594 20128 33600
rect 20272 33522 20300 34138
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 19248 32972 19300 32978
rect 19248 32914 19300 32920
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19260 31754 19288 32914
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20536 32224 20588 32230
rect 20536 32166 20588 32172
rect 20548 32026 20576 32166
rect 20536 32020 20588 32026
rect 20536 31962 20588 31968
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19168 31726 19288 31754
rect 19338 31784 19394 31793
rect 19168 31278 19196 31726
rect 19338 31719 19394 31728
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18524 29306 18552 29582
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18800 29170 18828 30194
rect 19168 30190 19196 31214
rect 19352 30938 19380 31719
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18524 28762 18552 28902
rect 18512 28756 18564 28762
rect 18512 28698 18564 28704
rect 18800 28558 18828 29106
rect 18984 28762 19012 29106
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 18788 28552 18840 28558
rect 18788 28494 18840 28500
rect 19076 28014 19104 28562
rect 19168 28558 19196 30126
rect 19352 29850 19380 30602
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 30326 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19996 30190 20024 31826
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 20088 31414 20116 31622
rect 20076 31408 20128 31414
rect 20076 31350 20128 31356
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19996 29646 20024 30126
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19156 28552 19208 28558
rect 19156 28494 19208 28500
rect 19168 28082 19196 28494
rect 19260 28422 19288 29106
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 19444 28490 19472 28970
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19260 28150 19288 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18432 26042 18460 26522
rect 19260 26382 19288 28086
rect 20272 28082 20300 28902
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19352 26042 19380 27270
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20640 27062 20668 39766
rect 20732 39370 20760 39902
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20824 37942 20852 43250
rect 21192 43110 21220 44270
rect 22204 43994 22232 44882
rect 22388 44538 22416 45222
rect 22652 44804 22704 44810
rect 22652 44746 22704 44752
rect 22376 44532 22428 44538
rect 22376 44474 22428 44480
rect 22664 44470 22692 44746
rect 22652 44464 22704 44470
rect 22572 44424 22652 44452
rect 22192 43988 22244 43994
rect 22192 43930 22244 43936
rect 21180 43104 21232 43110
rect 21180 43046 21232 43052
rect 21192 42702 21220 43046
rect 22572 42702 22600 44424
rect 22652 44406 22704 44412
rect 23400 44198 23428 45426
rect 23480 45416 23532 45422
rect 23480 45358 23532 45364
rect 23492 44742 23520 45358
rect 23572 45008 23624 45014
rect 23572 44950 23624 44956
rect 23480 44736 23532 44742
rect 23480 44678 23532 44684
rect 23492 44538 23520 44678
rect 23480 44532 23532 44538
rect 23480 44474 23532 44480
rect 23388 44192 23440 44198
rect 23388 44134 23440 44140
rect 22652 43648 22704 43654
rect 22652 43590 22704 43596
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 22560 42696 22612 42702
rect 22560 42638 22612 42644
rect 21192 41614 21220 42638
rect 21548 42628 21600 42634
rect 21548 42570 21600 42576
rect 21560 42362 21588 42570
rect 21548 42356 21600 42362
rect 21548 42298 21600 42304
rect 22284 42220 22336 42226
rect 22284 42162 22336 42168
rect 22296 42022 22324 42162
rect 22192 42016 22244 42022
rect 22192 41958 22244 41964
rect 22284 42016 22336 42022
rect 22284 41958 22336 41964
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 21456 41540 21508 41546
rect 21456 41482 21508 41488
rect 21468 41274 21496 41482
rect 21180 41268 21232 41274
rect 21180 41210 21232 41216
rect 21456 41268 21508 41274
rect 21456 41210 21508 41216
rect 20904 40384 20956 40390
rect 20904 40326 20956 40332
rect 20916 40118 20944 40326
rect 21192 40186 21220 41210
rect 22204 41206 22232 41958
rect 22192 41200 22244 41206
rect 22192 41142 22244 41148
rect 22572 41070 22600 42638
rect 22664 42226 22692 43590
rect 22836 42764 22888 42770
rect 22836 42706 22888 42712
rect 22848 42226 22876 42706
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 22836 42220 22888 42226
rect 22836 42162 22888 42168
rect 23112 42220 23164 42226
rect 23112 42162 23164 42168
rect 22928 42152 22980 42158
rect 22928 42094 22980 42100
rect 22836 42016 22888 42022
rect 22836 41958 22888 41964
rect 22744 41540 22796 41546
rect 22744 41482 22796 41488
rect 22560 41064 22612 41070
rect 22560 41006 22612 41012
rect 22652 40928 22704 40934
rect 22652 40870 22704 40876
rect 22664 40730 22692 40870
rect 22652 40724 22704 40730
rect 22652 40666 22704 40672
rect 21180 40180 21232 40186
rect 21180 40122 21232 40128
rect 20904 40112 20956 40118
rect 20904 40054 20956 40060
rect 20904 39976 20956 39982
rect 20904 39918 20956 39924
rect 20916 39642 20944 39918
rect 21088 39840 21140 39846
rect 21088 39782 21140 39788
rect 20904 39636 20956 39642
rect 20904 39578 20956 39584
rect 20916 39098 20944 39578
rect 21100 39302 21128 39782
rect 21192 39302 21220 40122
rect 21548 39840 21600 39846
rect 21548 39782 21600 39788
rect 21088 39296 21140 39302
rect 21088 39238 21140 39244
rect 21180 39296 21232 39302
rect 21180 39238 21232 39244
rect 21100 39098 21128 39238
rect 20904 39092 20956 39098
rect 20904 39034 20956 39040
rect 21088 39092 21140 39098
rect 21088 39034 21140 39040
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20996 38956 21048 38962
rect 20996 38898 21048 38904
rect 20916 38758 20944 38898
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20812 37936 20864 37942
rect 20812 37878 20864 37884
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20824 36922 20852 37130
rect 21008 37126 21036 38898
rect 21192 38826 21220 39238
rect 21560 39098 21588 39782
rect 21640 39500 21692 39506
rect 21640 39442 21692 39448
rect 21652 39098 21680 39442
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 22008 39364 22060 39370
rect 22008 39306 22060 39312
rect 22020 39098 22048 39306
rect 21548 39092 21600 39098
rect 21548 39034 21600 39040
rect 21640 39092 21692 39098
rect 21640 39034 21692 39040
rect 22008 39092 22060 39098
rect 22008 39034 22060 39040
rect 21180 38820 21232 38826
rect 21180 38762 21232 38768
rect 22296 38418 22324 39374
rect 22664 39370 22692 40666
rect 22756 40186 22784 41482
rect 22848 41138 22876 41958
rect 22940 41546 22968 42094
rect 23124 41614 23152 42162
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 23308 41818 23336 42094
rect 23296 41812 23348 41818
rect 23296 41754 23348 41760
rect 23112 41608 23164 41614
rect 23112 41550 23164 41556
rect 23204 41608 23256 41614
rect 23204 41550 23256 41556
rect 22928 41540 22980 41546
rect 22928 41482 22980 41488
rect 23216 41138 23244 41550
rect 23308 41206 23336 41754
rect 23400 41682 23428 44134
rect 23492 43790 23520 44474
rect 23584 43858 23612 44950
rect 23664 44872 23716 44878
rect 23664 44814 23716 44820
rect 23676 43994 23704 44814
rect 23756 44804 23808 44810
rect 23756 44746 23808 44752
rect 23664 43988 23716 43994
rect 23664 43930 23716 43936
rect 23572 43852 23624 43858
rect 23572 43794 23624 43800
rect 23480 43784 23532 43790
rect 23480 43726 23532 43732
rect 23768 43722 23796 44746
rect 23952 44538 23980 45426
rect 24032 45280 24084 45286
rect 24032 45222 24084 45228
rect 24044 45082 24072 45222
rect 24032 45076 24084 45082
rect 24032 45018 24084 45024
rect 24136 44878 24164 45426
rect 24124 44872 24176 44878
rect 24124 44814 24176 44820
rect 24400 44872 24452 44878
rect 24400 44814 24452 44820
rect 23940 44532 23992 44538
rect 24136 44520 24164 44814
rect 24216 44532 24268 44538
rect 24136 44492 24216 44520
rect 23940 44474 23992 44480
rect 24216 44474 24268 44480
rect 23756 43716 23808 43722
rect 23756 43658 23808 43664
rect 24412 42770 24440 44814
rect 24964 44690 24992 45766
rect 25872 45552 25924 45558
rect 25872 45494 25924 45500
rect 25136 45280 25188 45286
rect 25136 45222 25188 45228
rect 25504 45280 25556 45286
rect 25504 45222 25556 45228
rect 25148 44810 25176 45222
rect 25136 44804 25188 44810
rect 25188 44764 25268 44792
rect 25136 44746 25188 44752
rect 24964 44662 25176 44690
rect 25148 44266 25176 44662
rect 25136 44260 25188 44266
rect 25136 44202 25188 44208
rect 25240 42906 25268 44764
rect 25320 44192 25372 44198
rect 25320 44134 25372 44140
rect 25332 43790 25360 44134
rect 25320 43784 25372 43790
rect 25320 43726 25372 43732
rect 25228 42900 25280 42906
rect 25228 42842 25280 42848
rect 24400 42764 24452 42770
rect 24400 42706 24452 42712
rect 24032 42696 24084 42702
rect 24032 42638 24084 42644
rect 23480 42560 23532 42566
rect 23480 42502 23532 42508
rect 23848 42560 23900 42566
rect 23848 42502 23900 42508
rect 23388 41676 23440 41682
rect 23388 41618 23440 41624
rect 23492 41614 23520 42502
rect 23860 42362 23888 42502
rect 24044 42362 24072 42638
rect 23848 42356 23900 42362
rect 23848 42298 23900 42304
rect 24032 42356 24084 42362
rect 24032 42298 24084 42304
rect 23572 42288 23624 42294
rect 23572 42230 23624 42236
rect 23480 41608 23532 41614
rect 23480 41550 23532 41556
rect 23492 41274 23520 41550
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23296 41200 23348 41206
rect 23296 41142 23348 41148
rect 22836 41132 22888 41138
rect 22836 41074 22888 41080
rect 23204 41132 23256 41138
rect 23204 41074 23256 41080
rect 23480 41132 23532 41138
rect 23480 41074 23532 41080
rect 22744 40180 22796 40186
rect 22744 40122 22796 40128
rect 23492 40050 23520 41074
rect 23584 40202 23612 42230
rect 23940 41676 23992 41682
rect 23940 41618 23992 41624
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 23676 40526 23704 41006
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23584 40174 23796 40202
rect 23480 40044 23532 40050
rect 23480 39986 23532 39992
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 22652 39364 22704 39370
rect 22652 39306 22704 39312
rect 22284 38412 22336 38418
rect 22284 38354 22336 38360
rect 21456 38344 21508 38350
rect 21456 38286 21508 38292
rect 21468 38010 21496 38286
rect 21456 38004 21508 38010
rect 21456 37946 21508 37952
rect 21468 37330 21496 37946
rect 21456 37324 21508 37330
rect 21456 37266 21508 37272
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 21468 36854 21496 37266
rect 22284 37120 22336 37126
rect 22284 37062 22336 37068
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 21456 36848 21508 36854
rect 21456 36790 21508 36796
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20916 35698 20944 35974
rect 20904 35692 20956 35698
rect 20904 35634 20956 35640
rect 20996 34536 21048 34542
rect 20996 34478 21048 34484
rect 21008 32978 21036 34478
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21100 33810 21128 34342
rect 21178 33960 21234 33969
rect 21178 33895 21180 33904
rect 21232 33895 21234 33904
rect 21180 33866 21232 33872
rect 21100 33782 21220 33810
rect 20996 32972 21048 32978
rect 20996 32914 21048 32920
rect 21088 32360 21140 32366
rect 21088 32302 21140 32308
rect 21100 32026 21128 32302
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21192 31890 21220 33782
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21284 32842 21312 33254
rect 21272 32836 21324 32842
rect 21272 32778 21324 32784
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20824 30326 20852 31282
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 21192 29714 21220 31826
rect 21284 31822 21312 32370
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 21284 31482 21312 31758
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 21376 30138 21404 36654
rect 21468 36242 21496 36790
rect 21548 36576 21600 36582
rect 21548 36518 21600 36524
rect 21560 36310 21588 36518
rect 21548 36304 21600 36310
rect 21548 36246 21600 36252
rect 22296 36242 22324 37062
rect 21456 36236 21508 36242
rect 21456 36178 21508 36184
rect 22284 36236 22336 36242
rect 22284 36178 22336 36184
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21284 30110 21404 30138
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21284 28966 21312 30110
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 21284 28626 21312 28902
rect 21376 28762 21404 29106
rect 21468 28762 21496 35974
rect 22376 35624 22428 35630
rect 22376 35566 22428 35572
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 21560 34746 21588 35430
rect 22388 35290 22416 35566
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22480 35154 22508 37062
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22100 35012 22152 35018
rect 22100 34954 22152 34960
rect 21548 34740 21600 34746
rect 21548 34682 21600 34688
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 22020 34202 22048 34342
rect 22008 34196 22060 34202
rect 22008 34138 22060 34144
rect 22112 34066 22140 34954
rect 22664 34610 22692 39306
rect 23388 39296 23440 39302
rect 23388 39238 23440 39244
rect 23400 38826 23428 39238
rect 23480 38888 23532 38894
rect 23480 38830 23532 38836
rect 23572 38888 23624 38894
rect 23572 38830 23624 38836
rect 23388 38820 23440 38826
rect 23388 38762 23440 38768
rect 22836 38752 22888 38758
rect 22836 38694 22888 38700
rect 22848 38418 22876 38694
rect 22836 38412 22888 38418
rect 22836 38354 22888 38360
rect 23400 37874 23428 38762
rect 23492 38554 23520 38830
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23584 38010 23612 38830
rect 23572 38004 23624 38010
rect 23572 37946 23624 37952
rect 23676 37874 23704 39782
rect 23768 38962 23796 40174
rect 23756 38956 23808 38962
rect 23756 38898 23808 38904
rect 23388 37868 23440 37874
rect 23388 37810 23440 37816
rect 23480 37868 23532 37874
rect 23480 37810 23532 37816
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23492 37262 23520 37810
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22940 36922 22968 37062
rect 22928 36916 22980 36922
rect 22928 36858 22980 36864
rect 23676 36854 23704 37810
rect 23664 36848 23716 36854
rect 23664 36790 23716 36796
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 36378 23060 36722
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 23296 36236 23348 36242
rect 23296 36178 23348 36184
rect 23308 35630 23336 36178
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23308 35154 23336 35566
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 22652 34604 22704 34610
rect 22652 34546 22704 34552
rect 22284 34128 22336 34134
rect 22284 34070 22336 34076
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 22008 33856 22060 33862
rect 22008 33798 22060 33804
rect 21652 33658 21680 33798
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 21560 31482 21588 33526
rect 22020 32774 22048 33798
rect 22296 32842 22324 34070
rect 22284 32836 22336 32842
rect 22284 32778 22336 32784
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21824 32360 21876 32366
rect 21824 32302 21876 32308
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21836 31278 21864 32302
rect 22192 31952 22244 31958
rect 22192 31894 22244 31900
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 31414 22140 31622
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 21824 31272 21876 31278
rect 21824 31214 21876 31220
rect 21836 30938 21864 31214
rect 21548 30932 21600 30938
rect 21548 30874 21600 30880
rect 21824 30932 21876 30938
rect 21824 30874 21876 30880
rect 21560 29102 21588 30874
rect 22204 30326 22232 31894
rect 22296 31482 22324 32778
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22572 30666 22600 31622
rect 22560 30660 22612 30666
rect 22560 30602 22612 30608
rect 22192 30320 22244 30326
rect 22192 30262 22244 30268
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 21364 28756 21416 28762
rect 21364 28698 21416 28704
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21560 28082 21588 29038
rect 21744 28558 21772 29446
rect 22112 29238 22140 29446
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21744 28218 21772 28494
rect 21732 28212 21784 28218
rect 21732 28154 21784 28160
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21560 27674 21588 28018
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20628 27056 20680 27062
rect 20680 27004 20760 27010
rect 20628 26998 20760 27004
rect 20640 26982 20760 26998
rect 20824 26994 20852 27406
rect 20628 26920 20680 26926
rect 20548 26880 20628 26908
rect 20548 26450 20576 26880
rect 20628 26862 20680 26868
rect 20732 26738 20760 26982
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 21364 26852 21416 26858
rect 21364 26794 21416 26800
rect 20640 26710 20760 26738
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 26042 19472 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 18064 25226 18184 25242
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 18052 25220 18196 25226
rect 18104 25214 18144 25220
rect 18052 25162 18104 25168
rect 18144 25162 18196 25168
rect 17604 24954 17632 25162
rect 18340 24954 18368 25434
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 17592 24948 17644 24954
rect 17592 24890 17644 24896
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18616 24750 18644 25774
rect 17224 24744 17276 24750
rect 17224 24686 17276 24692
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23730 16712 24006
rect 16776 23866 16804 24346
rect 17236 23866 17264 24686
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17604 23866 17632 24074
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23866 18184 24006
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 16040 21622 16068 23054
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22778 16436 22918
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16592 22234 16620 22646
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16592 21690 16620 22170
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15108 19984 15160 19990
rect 15108 19926 15160 19932
rect 15120 19378 15148 19926
rect 15396 19786 15424 20198
rect 15948 19922 15976 20538
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15212 18834 15240 19450
rect 15488 19446 15516 19858
rect 16040 19786 16068 21558
rect 16684 21554 16712 22374
rect 16776 21554 16804 23122
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16868 22098 16896 23054
rect 17236 23050 17264 23802
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17788 23322 17816 23666
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 18156 23118 18184 23802
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17880 22778 17908 22986
rect 18432 22778 18460 24686
rect 18708 24410 18736 25842
rect 19352 24954 19380 25842
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19444 25294 19472 25774
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25498 19564 25638
rect 20272 25498 20300 26250
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 17236 21350 17264 22510
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17420 20942 17448 22034
rect 17880 21486 17908 22510
rect 18064 22234 18092 22578
rect 18432 22506 18460 22714
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 18156 22030 18184 22374
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17776 20868 17828 20874
rect 17776 20810 17828 20816
rect 17788 20602 17816 20810
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17880 20398 17908 21422
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 20602 18092 21286
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 16132 19514 16160 20334
rect 18340 20330 18368 21422
rect 18708 21146 18736 24142
rect 19444 23866 19472 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20272 24954 20300 25434
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22778 18920 22918
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 19076 21690 19104 21898
rect 19260 21894 19288 22986
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21690 19288 21830
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18708 20602 18736 21082
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15488 18834 15516 19382
rect 16040 19242 16068 19450
rect 16776 19446 16804 19790
rect 17696 19514 17724 19790
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15948 18766 15976 19110
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 15120 18358 15148 18566
rect 16776 18426 16804 19246
rect 17972 18902 18000 20266
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18064 18970 18092 19246
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18340 18766 18368 19246
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18432 18612 18460 20334
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19514 18736 19654
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18340 18584 18460 18612
rect 18340 18426 18368 18584
rect 18984 18426 19012 18634
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 18340 18222 18368 18362
rect 19168 18290 19196 18906
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15580 17678 15608 18022
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17338 15700 17478
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14844 16114 14872 16594
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14830 15872 14886 15881
rect 14830 15807 14886 15816
rect 14554 15600 14610 15609
rect 14554 15535 14610 15544
rect 14568 15162 14596 15535
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14618 14136 14962
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14292 14074 14320 14826
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14004 13864 14056 13870
rect 14002 13832 14004 13841
rect 14056 13832 14058 13841
rect 14002 13767 14058 13776
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14002 12608 14058 12617
rect 14002 12543 14058 12552
rect 14016 12442 14044 12543
rect 14108 12442 14136 14010
rect 14278 13968 14334 13977
rect 14278 13903 14280 13912
rect 14332 13903 14334 13912
rect 14280 13874 14332 13880
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14200 12322 14228 13806
rect 14384 12322 14412 14758
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14568 13938 14596 14214
rect 14660 13938 14688 15302
rect 14738 14240 14794 14249
rect 14738 14175 14794 14184
rect 14752 14074 14780 14175
rect 14740 14068 14792 14074
rect 14844 14056 14872 15807
rect 14936 15570 14964 16118
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14844 14028 14964 14056
rect 14740 14010 14792 14016
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13394 14780 13670
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14844 12986 14872 13874
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14936 12866 14964 14028
rect 14660 12838 14964 12866
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12434 14596 12718
rect 14016 12294 14228 12322
rect 14292 12294 14412 12322
rect 14476 12406 14596 12434
rect 14016 12238 14044 12294
rect 14292 12238 14320 12294
rect 14476 12238 14504 12406
rect 14660 12238 14688 12838
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13648 10742 13676 11698
rect 13832 11665 13860 11698
rect 14016 11694 14044 12174
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14004 11688 14056 11694
rect 13818 11656 13874 11665
rect 14004 11630 14056 11636
rect 13818 11591 13874 11600
rect 13820 11552 13872 11558
rect 13740 11512 13820 11540
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13740 10538 13768 11512
rect 14016 11506 14044 11630
rect 13820 11494 13872 11500
rect 13924 11478 14044 11506
rect 13818 10840 13874 10849
rect 13818 10775 13874 10784
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13740 9674 13768 10474
rect 13832 10470 13860 10775
rect 13924 10606 13952 11478
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13556 9646 13768 9674
rect 13556 9586 13584 9646
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13924 9518 13952 10542
rect 14108 10033 14136 11018
rect 14200 10130 14228 11698
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14292 10062 14320 12174
rect 14384 11898 14412 12174
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14476 11762 14504 12038
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 11286 14504 11698
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14280 10056 14332 10062
rect 14094 10024 14150 10033
rect 14280 9998 14332 10004
rect 14094 9959 14150 9968
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13832 9178 13860 9454
rect 14108 9382 14136 9959
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14016 9042 14044 9318
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8838 13860 8910
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13740 8566 13768 8774
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 14384 8498 14412 9454
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13740 7546 13768 8026
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 13542 6896 13598 6905
rect 13542 6831 13598 6840
rect 13556 6662 13584 6831
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13372 5778 13400 6122
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 12530 5607 12586 5616
rect 13084 5636 13136 5642
rect 10968 5578 11020 5584
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10612 4690 10640 5170
rect 10980 5166 11008 5578
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 3602 10640 4626
rect 10980 4214 11008 5102
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4690 12020 4966
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11992 4214 12020 4490
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3602 11560 3878
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 11992 3466 12020 4150
rect 12544 4078 12572 5607
rect 13084 5578 13136 5584
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 4282 12664 5170
rect 13096 4758 13124 5578
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4758 13216 5102
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13556 4622 13584 6598
rect 13832 6322 13860 6666
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13648 5710 13676 6258
rect 14108 6254 14136 6734
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 5846 14136 6054
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14016 5710 14044 5782
rect 14292 5710 14320 7414
rect 14476 7410 14504 11222
rect 14568 11218 14596 11766
rect 14660 11354 14688 12174
rect 14752 11898 14780 12174
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11778 14872 12582
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14936 12102 14964 12378
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14752 11750 14872 11778
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10470 14596 11154
rect 14752 11150 14780 11750
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14832 11144 14884 11150
rect 14936 11132 14964 12038
rect 15028 11898 15056 16050
rect 15120 15706 15148 16526
rect 15304 16250 15332 17138
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15108 15700 15160 15706
rect 15488 15688 15516 17138
rect 15856 16522 15884 17138
rect 15948 16658 15976 17206
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 17512 17190 17724 17218
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16132 16658 16160 16934
rect 16408 16658 16436 17002
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 15844 16516 15896 16522
rect 15896 16476 15976 16504
rect 15844 16458 15896 16464
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15580 16114 15608 16390
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15108 15642 15160 15648
rect 15304 15660 15516 15688
rect 15304 15570 15332 15660
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 15162 15240 15438
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 14618 15332 15370
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14657 15608 14758
rect 15566 14648 15622 14657
rect 15292 14612 15344 14618
rect 15566 14583 15622 14592
rect 15292 14554 15344 14560
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15120 14278 15148 14350
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15304 14074 15332 14554
rect 15580 14482 15608 14583
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15396 13954 15424 14214
rect 15672 14090 15700 15574
rect 15764 15570 15792 15846
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15764 14346 15792 14962
rect 15856 14618 15884 15438
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15304 13926 15424 13954
rect 15580 14062 15700 14090
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12442 15148 13330
rect 15212 12850 15240 13806
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15198 12744 15254 12753
rect 15198 12679 15254 12688
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15212 12374 15240 12679
rect 15304 12442 15332 13926
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12782 15516 13262
rect 15476 12776 15528 12782
rect 15396 12736 15476 12764
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15120 11744 15148 12106
rect 15212 12073 15240 12174
rect 15198 12064 15254 12073
rect 15198 11999 15254 12008
rect 15028 11716 15148 11744
rect 15028 11393 15056 11716
rect 15014 11384 15070 11393
rect 15014 11319 15070 11328
rect 14884 11104 14964 11132
rect 14832 11086 14884 11092
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14660 10062 14688 10406
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9586 14596 9862
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14660 9042 14688 9590
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8430 14596 8842
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14384 6254 14412 6734
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14384 5914 14412 6190
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 13648 5370 13676 5646
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13924 5302 13952 5646
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 14384 5030 14412 5850
rect 14568 5760 14596 8366
rect 14660 6798 14688 8774
rect 14752 7410 14780 11086
rect 14844 10742 14872 11086
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14844 9382 14872 10678
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14844 8566 14872 9114
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14936 8362 14964 10610
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7546 14872 7686
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14752 6322 14780 7346
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 6322 14872 7210
rect 14936 6798 14964 7346
rect 15028 6934 15056 11319
rect 15212 11234 15240 11999
rect 15396 11898 15424 12736
rect 15476 12718 15528 12724
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15488 12102 15516 12378
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15290 11792 15346 11801
rect 15290 11727 15292 11736
rect 15344 11727 15346 11736
rect 15292 11698 15344 11704
rect 15212 11206 15332 11234
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10606 15240 11086
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15304 9654 15332 11206
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15396 10985 15424 11086
rect 15382 10976 15438 10985
rect 15382 10911 15438 10920
rect 15396 10470 15424 10911
rect 15488 10742 15516 11086
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15580 10266 15608 14062
rect 15764 13938 15792 14282
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15672 12782 15700 13874
rect 15660 12776 15712 12782
rect 15658 12744 15660 12753
rect 15712 12744 15714 12753
rect 15658 12679 15714 12688
rect 15658 12608 15714 12617
rect 15658 12543 15714 12552
rect 15672 12374 15700 12543
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15672 9110 15700 11086
rect 15764 10742 15792 13874
rect 15856 13841 15884 14554
rect 15948 14278 15976 16476
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16040 15502 16068 15914
rect 16132 15881 16160 15982
rect 16118 15872 16174 15881
rect 16118 15807 16174 15816
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16040 14414 16068 15438
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15842 13832 15898 13841
rect 15842 13767 15898 13776
rect 15948 13190 15976 13874
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15856 10606 15884 12922
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11286 15976 12174
rect 16040 11370 16068 14350
rect 16316 13734 16344 15030
rect 16500 14482 16528 17138
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16868 16794 16896 17070
rect 17512 17066 17540 17190
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17604 16794 17632 17070
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17052 16114 17080 16186
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16776 15502 16804 15846
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16684 15026 16712 15370
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16776 14906 16804 15438
rect 16684 14878 16804 14906
rect 16684 14482 16712 14878
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14550 16804 14758
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13938 16436 14214
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16132 12306 16160 12582
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16212 12232 16264 12238
rect 16132 12180 16212 12186
rect 16132 12174 16264 12180
rect 16132 12158 16252 12174
rect 16132 11558 16160 12158
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16040 11342 16160 11370
rect 16224 11354 16252 12038
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10810 15976 11086
rect 16132 11082 16160 11342
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16316 10674 16344 13670
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16132 10130 16160 10406
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 9722 16252 9998
rect 16316 9722 16344 10406
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 15750 9616 15806 9625
rect 15750 9551 15806 9560
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 8634 15700 9046
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15120 6322 15148 8434
rect 15488 7954 15516 8434
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15488 7546 15516 7890
rect 15764 7562 15792 9551
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8430 15884 8910
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 8634 15976 8774
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15672 7534 15792 7562
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15212 6390 15240 6802
rect 15672 6798 15700 7534
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15764 7206 15792 7414
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6798 15792 7142
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15672 6662 15700 6734
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15304 6458 15332 6598
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15474 6352 15530 6361
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15292 6316 15344 6322
rect 15948 6322 15976 6938
rect 16040 6866 16068 9658
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16224 8974 16252 9522
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16316 7206 16344 9658
rect 16408 9450 16436 13874
rect 16500 12986 16528 14418
rect 16684 13977 16712 14418
rect 16670 13968 16726 13977
rect 16670 13903 16726 13912
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16592 13326 16620 13806
rect 16684 13462 16712 13806
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12986 16712 13194
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16684 12850 16712 12922
rect 16776 12918 16804 13126
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11665 16528 12174
rect 16486 11656 16542 11665
rect 16486 11591 16542 11600
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16592 11014 16620 11154
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 10282 16620 10542
rect 16500 10254 16620 10282
rect 16500 9625 16528 10254
rect 16684 10130 16712 12582
rect 16868 11370 16896 15982
rect 17052 15162 17080 16050
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14482 16988 14894
rect 17040 14816 17092 14822
rect 17038 14784 17040 14793
rect 17092 14784 17094 14793
rect 17038 14719 17094 14728
rect 17144 14521 17172 16390
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17236 15337 17264 16050
rect 17420 15502 17448 16050
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17408 15360 17460 15366
rect 17222 15328 17278 15337
rect 17408 15302 17460 15308
rect 17222 15263 17278 15272
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17130 14512 17186 14521
rect 16948 14476 17000 14482
rect 17130 14447 17186 14456
rect 16948 14418 17000 14424
rect 17040 14408 17092 14414
rect 17144 14396 17172 14447
rect 17328 14414 17356 15098
rect 17420 14618 17448 15302
rect 17512 15094 17540 16594
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17604 14929 17632 15506
rect 17696 15065 17724 17190
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 17788 15910 17816 17070
rect 17880 16046 17908 17070
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 18064 15706 18092 16390
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17684 14952 17736 14958
rect 17590 14920 17646 14929
rect 17684 14894 17736 14900
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17590 14855 17646 14864
rect 17592 14816 17644 14822
rect 17590 14784 17592 14793
rect 17644 14784 17646 14793
rect 17590 14719 17646 14728
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17092 14368 17172 14396
rect 17316 14408 17368 14414
rect 17040 14350 17092 14356
rect 17316 14350 17368 14356
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17052 13734 17080 14350
rect 17512 13870 17540 14350
rect 17316 13864 17368 13870
rect 17314 13832 17316 13841
rect 17500 13864 17552 13870
rect 17368 13832 17370 13841
rect 17500 13806 17552 13812
rect 17314 13767 17370 13776
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17224 13728 17276 13734
rect 17512 13716 17540 13806
rect 17604 13734 17632 14719
rect 17224 13670 17276 13676
rect 17328 13688 17540 13716
rect 17592 13728 17644 13734
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17052 12374 17080 12582
rect 17236 12434 17264 13670
rect 17144 12406 17264 12434
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 11762 16988 12174
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16776 11342 16896 11370
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16486 9616 16542 9625
rect 16684 9586 16712 9862
rect 16486 9551 16542 9560
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16580 9512 16632 9518
rect 16632 9460 16712 9466
rect 16580 9454 16712 9460
rect 16396 9444 16448 9450
rect 16592 9438 16712 9454
rect 16396 9386 16448 9392
rect 16408 9042 16436 9386
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8566 16528 8910
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16592 7886 16620 9318
rect 16684 9092 16712 9438
rect 16776 9364 16804 11342
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10266 16896 11086
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9674 16896 10066
rect 16960 10062 16988 11698
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17052 10305 17080 10678
rect 17038 10296 17094 10305
rect 17038 10231 17094 10240
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16868 9646 16988 9674
rect 16856 9376 16908 9382
rect 16776 9336 16856 9364
rect 16856 9318 16908 9324
rect 16764 9104 16816 9110
rect 16684 9064 16764 9092
rect 16764 9046 16816 9052
rect 16670 8936 16726 8945
rect 16670 8871 16672 8880
rect 16724 8871 16726 8880
rect 16672 8842 16724 8848
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8362 16804 8774
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16486 6896 16542 6905
rect 16028 6860 16080 6866
rect 16486 6831 16542 6840
rect 16028 6802 16080 6808
rect 16040 6322 16068 6802
rect 16500 6798 16528 6831
rect 16868 6798 16896 9318
rect 16960 8820 16988 9646
rect 17144 9178 17172 12406
rect 17328 12306 17356 13688
rect 17592 13670 17644 13676
rect 17696 12617 17724 14894
rect 17788 14074 17816 14894
rect 17880 14414 17908 15642
rect 18156 15434 18184 16390
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17958 14648 18014 14657
rect 17958 14583 18014 14592
rect 17972 14482 18000 14583
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17880 13920 17908 14350
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17788 13892 17908 13920
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17316 11212 17368 11218
rect 17236 11172 17316 11200
rect 17236 11121 17264 11172
rect 17316 11154 17368 11160
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17222 11112 17278 11121
rect 17222 11047 17278 11056
rect 17224 11008 17276 11014
rect 17408 11008 17460 11014
rect 17224 10950 17276 10956
rect 17328 10968 17408 10996
rect 17236 10810 17264 10950
rect 17328 10849 17356 10968
rect 17408 10950 17460 10956
rect 17314 10840 17370 10849
rect 17224 10804 17276 10810
rect 17314 10775 17370 10784
rect 17224 10746 17276 10752
rect 17512 10674 17540 11154
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17236 10441 17264 10474
rect 17222 10432 17278 10441
rect 17222 10367 17278 10376
rect 17222 9616 17278 9625
rect 17278 9560 17356 9568
rect 17222 9551 17224 9560
rect 17276 9540 17356 9560
rect 17224 9522 17276 9528
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17222 8936 17278 8945
rect 17132 8900 17184 8906
rect 17222 8871 17278 8880
rect 17132 8842 17184 8848
rect 17040 8832 17092 8838
rect 16960 8792 17040 8820
rect 16960 8430 16988 8792
rect 17040 8774 17092 8780
rect 17144 8498 17172 8842
rect 17236 8838 17264 8871
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 15474 6287 15476 6296
rect 15292 6258 15344 6264
rect 15528 6287 15530 6296
rect 15936 6316 15988 6322
rect 15476 6258 15528 6264
rect 15936 6258 15988 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 14752 6118 14780 6258
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14648 5772 14700 5778
rect 14568 5732 14648 5760
rect 14648 5714 14700 5720
rect 14844 5370 14872 6258
rect 15120 5574 15148 6258
rect 15304 5778 15332 6258
rect 15948 6118 15976 6258
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15396 5914 15424 6054
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5574 15240 5646
rect 16040 5642 16068 6258
rect 16224 5710 16252 6734
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 5710 16528 6258
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5914 16988 6190
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 12544 3074 12572 4014
rect 13004 3738 13032 4082
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12176 3058 12572 3074
rect 12728 3058 12756 3334
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 12164 3052 12572 3058
rect 12216 3046 12572 3052
rect 12716 3052 12768 3058
rect 12164 2994 12216 3000
rect 12716 2994 12768 3000
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10520 2650 10548 2858
rect 12084 2650 12112 2926
rect 12820 2922 12848 3470
rect 12912 3194 12940 3538
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13556 2990 13584 4422
rect 13648 4078 13676 4626
rect 14108 4146 14136 4966
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 3058 13676 4014
rect 14108 3602 14136 4082
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14292 3602 14320 4014
rect 15212 4010 15240 5510
rect 15580 5302 15608 5578
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15580 4214 15608 5238
rect 17052 5234 17080 7278
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17328 6798 17356 9540
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17420 8974 17448 9386
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7546 17448 8230
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 6662 17448 6734
rect 17408 6656 17460 6662
rect 17130 6624 17186 6633
rect 17408 6598 17460 6604
rect 17130 6559 17186 6568
rect 17144 6322 17172 6559
rect 17420 6322 17448 6598
rect 17512 6390 17540 10610
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8838 17632 9318
rect 17788 9178 17816 13892
rect 17972 13326 18000 14282
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17880 10130 17908 12786
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11354 18000 11494
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17960 11144 18012 11150
rect 17958 11112 17960 11121
rect 18012 11112 18014 11121
rect 17958 11047 18014 11056
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10470 18000 10950
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17880 10033 17908 10066
rect 18064 10062 18092 15030
rect 18156 14618 18184 15370
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 11082 18184 14418
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12850 18276 13194
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18340 12714 18368 15302
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11218 18276 12038
rect 18432 11898 18460 16594
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 15162 18552 16526
rect 18708 16454 18736 17070
rect 18800 16794 18828 18158
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18984 16590 19012 17002
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 16114 18736 16390
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18602 15736 18658 15745
rect 18602 15671 18658 15680
rect 18616 15162 18644 15671
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18524 14006 18552 14962
rect 18616 14249 18644 14962
rect 18602 14240 18658 14249
rect 18602 14175 18658 14184
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18524 12102 18552 13942
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12238 18644 12786
rect 18708 12782 18736 16050
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18800 12986 18828 13942
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18340 11257 18368 11494
rect 18326 11248 18382 11257
rect 18236 11212 18288 11218
rect 18326 11183 18382 11192
rect 18236 11154 18288 11160
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18052 10056 18104 10062
rect 17866 10024 17922 10033
rect 18052 9998 18104 10004
rect 17866 9959 17922 9968
rect 18064 9586 18092 9998
rect 18156 9674 18184 11018
rect 18156 9646 18276 9674
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 9178 18092 9522
rect 18248 9450 18276 9646
rect 18432 9489 18460 11834
rect 18616 11778 18644 12174
rect 18524 11750 18644 11778
rect 18524 10538 18552 11750
rect 18604 11688 18656 11694
rect 18656 11648 18736 11676
rect 18604 11630 18656 11636
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18616 10985 18644 11018
rect 18602 10976 18658 10985
rect 18602 10911 18658 10920
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18418 9480 18474 9489
rect 18236 9444 18288 9450
rect 18418 9415 18474 9424
rect 18236 9386 18288 9392
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17604 8498 17632 8774
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17604 5778 17632 8434
rect 17684 7880 17736 7886
rect 17736 7840 17816 7868
rect 17684 7822 17736 7828
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7546 17724 7686
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17788 7002 17816 7840
rect 17972 7410 18000 9046
rect 18156 7886 18184 9318
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18340 7410 18368 7686
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 7002 18000 7210
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18340 6905 18368 7346
rect 18326 6896 18382 6905
rect 18326 6831 18382 6840
rect 18524 6798 18552 9522
rect 18616 9217 18644 10911
rect 18708 10810 18736 11648
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18602 9208 18658 9217
rect 18602 9143 18658 9152
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 17696 6458 17724 6734
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 18248 5914 18276 6734
rect 18432 6254 18460 6734
rect 18524 6390 18552 6734
rect 18604 6724 18656 6730
rect 18708 6712 18736 9386
rect 18800 8090 18828 12582
rect 18892 10674 18920 14350
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 13734 19012 14214
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11898 19012 12038
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18984 11393 19012 11562
rect 18970 11384 19026 11393
rect 19076 11354 19104 18090
rect 19260 17270 19288 21422
rect 19444 20058 19472 23666
rect 19812 23254 19840 23666
rect 20088 23322 20116 23666
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19800 23248 19852 23254
rect 19800 23190 19852 23196
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22438 20024 23122
rect 20272 23118 20300 24074
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21486 20024 22374
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19628 19990 19656 20402
rect 19996 20398 20024 21422
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 19996 19922 20024 20334
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 17338 20024 19654
rect 20088 19514 20116 20470
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20364 17338 20392 24686
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19248 17128 19300 17134
rect 19300 17088 19380 17116
rect 19248 17070 19300 17076
rect 19352 15366 19380 17088
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19444 16250 19472 16934
rect 20272 16794 20300 16934
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 19536 15450 19564 15846
rect 19798 15736 19854 15745
rect 19444 15422 19564 15450
rect 19720 15694 19798 15722
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19168 14521 19196 14826
rect 19248 14544 19300 14550
rect 19154 14512 19210 14521
rect 19248 14486 19300 14492
rect 19154 14447 19210 14456
rect 19168 14414 19196 14447
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19168 13870 19196 14350
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12918 19196 13262
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 11830 19196 12718
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 18970 11319 19026 11328
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19168 11234 19196 11766
rect 18984 11206 19196 11234
rect 18984 11121 19012 11206
rect 18970 11112 19026 11121
rect 18970 11047 19026 11056
rect 19154 11112 19210 11121
rect 19154 11047 19156 11056
rect 18984 10792 19012 11047
rect 19208 11047 19210 11056
rect 19156 11018 19208 11024
rect 19064 11008 19116 11014
rect 19116 10956 19196 10962
rect 19064 10950 19196 10956
rect 19076 10934 19196 10950
rect 19168 10810 19196 10934
rect 19156 10804 19208 10810
rect 18984 10764 19104 10792
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18880 10532 18932 10538
rect 18880 10474 18932 10480
rect 18892 9518 18920 10474
rect 18984 9926 19012 10610
rect 19076 10470 19104 10764
rect 19156 10746 19208 10752
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 9654 19012 9862
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18800 7002 18828 8026
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18656 6684 18736 6712
rect 18604 6666 18656 6672
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18616 6118 18644 6666
rect 18892 6254 18920 9454
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18984 7478 19012 8366
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 19076 6361 19104 10202
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9382 19196 9862
rect 19156 9376 19208 9382
rect 19260 9364 19288 14486
rect 19444 14362 19472 15422
rect 19720 15366 19748 15694
rect 19798 15671 19854 15680
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19522 15056 19578 15065
rect 19996 15026 20024 15302
rect 19522 14991 19578 15000
rect 19984 15020 20036 15026
rect 19536 14396 19564 14991
rect 19984 14962 20036 14968
rect 20088 14958 20116 15302
rect 20180 15026 20208 15846
rect 20456 15586 20484 26318
rect 20548 24750 20576 26386
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20640 22710 20668 26710
rect 21376 26450 21404 26794
rect 21560 26450 21588 27610
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 21548 26444 21600 26450
rect 21548 26386 21600 26392
rect 21376 26042 21404 26386
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 26042 21680 26250
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21640 26036 21692 26042
rect 21640 25978 21692 25984
rect 22020 24818 22048 28562
rect 22664 27470 22692 34546
rect 23112 32564 23164 32570
rect 23112 32506 23164 32512
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22756 32026 22784 32166
rect 22848 32026 22876 32370
rect 22744 32020 22796 32026
rect 22744 31962 22796 31968
rect 22836 32020 22888 32026
rect 22836 31962 22888 31968
rect 23124 31890 23152 32506
rect 23308 32042 23336 35090
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34746 23428 35022
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23492 32910 23520 33934
rect 23952 33590 23980 41618
rect 24412 41070 24440 42706
rect 25240 42634 25268 42842
rect 25228 42628 25280 42634
rect 25228 42570 25280 42576
rect 25044 42220 25096 42226
rect 25044 42162 25096 42168
rect 25056 41478 25084 42162
rect 25044 41472 25096 41478
rect 25044 41414 25096 41420
rect 25240 41206 25268 42570
rect 25516 42566 25544 45222
rect 25688 44736 25740 44742
rect 25688 44678 25740 44684
rect 25700 44334 25728 44678
rect 25884 44402 25912 45494
rect 26700 45416 26752 45422
rect 26700 45358 26752 45364
rect 26424 45280 26476 45286
rect 26424 45222 26476 45228
rect 26240 44872 26292 44878
rect 26240 44814 26292 44820
rect 25872 44396 25924 44402
rect 25872 44338 25924 44344
rect 25688 44328 25740 44334
rect 25688 44270 25740 44276
rect 26252 43858 26280 44814
rect 26436 44470 26464 45222
rect 26516 44804 26568 44810
rect 26516 44746 26568 44752
rect 26528 44538 26556 44746
rect 26712 44538 26740 45358
rect 27160 45280 27212 45286
rect 27160 45222 27212 45228
rect 26516 44532 26568 44538
rect 26516 44474 26568 44480
rect 26700 44532 26752 44538
rect 26700 44474 26752 44480
rect 27172 44470 27200 45222
rect 27540 44470 27568 45766
rect 27908 45626 27936 45902
rect 41972 45892 42024 45898
rect 41972 45834 42024 45840
rect 29092 45824 29144 45830
rect 29092 45766 29144 45772
rect 32036 45824 32088 45830
rect 32036 45766 32088 45772
rect 27896 45620 27948 45626
rect 27896 45562 27948 45568
rect 26424 44464 26476 44470
rect 26424 44406 26476 44412
rect 27160 44464 27212 44470
rect 27160 44406 27212 44412
rect 27528 44464 27580 44470
rect 27528 44406 27580 44412
rect 26516 44396 26568 44402
rect 26516 44338 26568 44344
rect 26528 44198 26556 44338
rect 26976 44328 27028 44334
rect 26976 44270 27028 44276
rect 26516 44192 26568 44198
rect 26516 44134 26568 44140
rect 26988 43858 27016 44270
rect 27908 44198 27936 45562
rect 28080 45552 28132 45558
rect 28080 45494 28132 45500
rect 28092 45082 28120 45494
rect 28540 45484 28592 45490
rect 28540 45426 28592 45432
rect 28080 45076 28132 45082
rect 28080 45018 28132 45024
rect 28552 44810 28580 45426
rect 29104 44946 29132 45766
rect 29644 45416 29696 45422
rect 29644 45358 29696 45364
rect 29920 45416 29972 45422
rect 29920 45358 29972 45364
rect 29656 45082 29684 45358
rect 29644 45076 29696 45082
rect 29644 45018 29696 45024
rect 29092 44940 29144 44946
rect 29092 44882 29144 44888
rect 28540 44804 28592 44810
rect 28540 44746 28592 44752
rect 28080 44736 28132 44742
rect 28080 44678 28132 44684
rect 28092 44538 28120 44678
rect 28080 44532 28132 44538
rect 28080 44474 28132 44480
rect 28552 44402 28580 44746
rect 28540 44396 28592 44402
rect 28540 44338 28592 44344
rect 27896 44192 27948 44198
rect 27896 44134 27948 44140
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 26976 43852 27028 43858
rect 26976 43794 27028 43800
rect 26252 42770 26280 43794
rect 28552 43654 28580 44338
rect 29932 43858 29960 45358
rect 30012 45280 30064 45286
rect 30012 45222 30064 45228
rect 30024 45082 30052 45222
rect 30012 45076 30064 45082
rect 30012 45018 30064 45024
rect 29920 43852 29972 43858
rect 29920 43794 29972 43800
rect 31852 43852 31904 43858
rect 31852 43794 31904 43800
rect 27712 43648 27764 43654
rect 27712 43590 27764 43596
rect 28540 43648 28592 43654
rect 28540 43590 28592 43596
rect 26792 43308 26844 43314
rect 26792 43250 26844 43256
rect 26884 43308 26936 43314
rect 26884 43250 26936 43256
rect 26240 42764 26292 42770
rect 26240 42706 26292 42712
rect 26700 42764 26752 42770
rect 26700 42706 26752 42712
rect 26712 42566 26740 42706
rect 25504 42560 25556 42566
rect 25504 42502 25556 42508
rect 26148 42560 26200 42566
rect 26148 42502 26200 42508
rect 26700 42560 26752 42566
rect 26700 42502 26752 42508
rect 25320 41268 25372 41274
rect 25320 41210 25372 41216
rect 25228 41200 25280 41206
rect 25228 41142 25280 41148
rect 24400 41064 24452 41070
rect 24400 41006 24452 41012
rect 24676 41064 24728 41070
rect 24676 41006 24728 41012
rect 24124 40384 24176 40390
rect 24124 40326 24176 40332
rect 24136 38894 24164 40326
rect 24412 39506 24440 41006
rect 24492 40928 24544 40934
rect 24544 40876 24624 40882
rect 24492 40870 24624 40876
rect 24504 40854 24624 40870
rect 24596 39982 24624 40854
rect 24688 40730 24716 41006
rect 24676 40724 24728 40730
rect 24676 40666 24728 40672
rect 25332 40662 25360 41210
rect 25320 40656 25372 40662
rect 25320 40598 25372 40604
rect 24584 39976 24636 39982
rect 24584 39918 24636 39924
rect 24400 39500 24452 39506
rect 24400 39442 24452 39448
rect 24596 39030 24624 39918
rect 24676 39364 24728 39370
rect 24676 39306 24728 39312
rect 24688 39098 24716 39306
rect 24676 39092 24728 39098
rect 24676 39034 24728 39040
rect 24584 39024 24636 39030
rect 24584 38966 24636 38972
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 24136 37874 24164 38830
rect 24768 38820 24820 38826
rect 24768 38762 24820 38768
rect 24400 38208 24452 38214
rect 24400 38150 24452 38156
rect 24412 38010 24440 38150
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 36922 24440 37198
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24780 36786 24808 38762
rect 25044 37800 25096 37806
rect 25044 37742 25096 37748
rect 25136 37800 25188 37806
rect 25136 37742 25188 37748
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24872 36786 24900 37062
rect 25056 36854 25084 37742
rect 25148 36922 25176 37742
rect 25228 37256 25280 37262
rect 25228 37198 25280 37204
rect 25136 36916 25188 36922
rect 25136 36858 25188 36864
rect 25044 36848 25096 36854
rect 25044 36790 25096 36796
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24872 36174 24900 36722
rect 25240 36242 25268 37198
rect 25228 36236 25280 36242
rect 25228 36178 25280 36184
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24412 35834 24440 35974
rect 24400 35828 24452 35834
rect 24400 35770 24452 35776
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24044 34746 24072 35022
rect 24584 34944 24636 34950
rect 24636 34892 24716 34898
rect 24584 34886 24716 34892
rect 24596 34870 24716 34886
rect 24032 34740 24084 34746
rect 24032 34682 24084 34688
rect 24688 34610 24716 34870
rect 24780 34746 24808 35974
rect 25240 35494 25268 36178
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 24768 34740 24820 34746
rect 24768 34682 24820 34688
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24398 34096 24454 34105
rect 24398 34031 24454 34040
rect 24412 33658 24440 34031
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 23940 33584 23992 33590
rect 23940 33526 23992 33532
rect 23952 33386 23980 33526
rect 23940 33380 23992 33386
rect 23940 33322 23992 33328
rect 24504 32978 24532 34478
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24596 33114 24624 33934
rect 24688 33454 24716 34546
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25240 33658 25268 33798
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24676 33448 24728 33454
rect 24676 33390 24728 33396
rect 24780 33114 24808 33458
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 24492 32972 24544 32978
rect 24492 32914 24544 32920
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23308 32014 23520 32042
rect 23388 31952 23440 31958
rect 23216 31900 23388 31906
rect 23216 31894 23440 31900
rect 23216 31890 23428 31894
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 23204 31884 23428 31890
rect 23256 31878 23428 31884
rect 23204 31826 23256 31832
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22848 29306 22876 30126
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22848 28558 22876 29242
rect 22940 28762 22968 29582
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22204 27130 22232 27406
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22480 25838 22508 26998
rect 22664 26994 22692 27406
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22848 25922 22876 26862
rect 23032 26518 23060 28358
rect 23124 27606 23152 31826
rect 23308 28626 23336 31878
rect 23492 31770 23520 32014
rect 23400 31742 23520 31770
rect 23584 31754 23612 32166
rect 24504 31958 24532 32914
rect 24584 32836 24636 32842
rect 24584 32778 24636 32784
rect 24492 31952 24544 31958
rect 24492 31894 24544 31900
rect 24216 31884 24268 31890
rect 24216 31826 24268 31832
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23572 31748 23624 31754
rect 23296 28620 23348 28626
rect 23400 28608 23428 31742
rect 23572 31690 23624 31696
rect 23676 31482 23704 31758
rect 24124 31680 24176 31686
rect 24124 31622 24176 31628
rect 24136 31482 24164 31622
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 24124 31476 24176 31482
rect 24124 31418 24176 31424
rect 24136 30394 24164 31418
rect 24228 31278 24256 31826
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 24216 30592 24268 30598
rect 24216 30534 24268 30540
rect 24124 30388 24176 30394
rect 24124 30330 24176 30336
rect 24228 30258 24256 30534
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24596 30122 24624 32778
rect 24780 32502 24808 33050
rect 25056 32910 25084 33594
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24780 31414 24808 31622
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24780 30734 24808 31078
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 24584 30116 24636 30122
rect 24584 30058 24636 30064
rect 24400 29572 24452 29578
rect 24400 29514 24452 29520
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23480 28620 23532 28626
rect 23400 28580 23480 28608
rect 23296 28562 23348 28568
rect 23480 28562 23532 28568
rect 23492 28014 23520 28562
rect 23768 28218 23796 29106
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 23940 28552 23992 28558
rect 23940 28494 23992 28500
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23124 27130 23152 27542
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23492 26926 23520 27950
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 26042 23060 26182
rect 23020 26036 23072 26042
rect 23020 25978 23072 25984
rect 22848 25894 22968 25922
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24206 21956 24686
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21928 23662 21956 24142
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 22296 23202 22324 25774
rect 22848 25498 22876 25774
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22388 24954 22416 25094
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22388 23322 22416 24278
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22204 23174 22324 23202
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22778 20760 23054
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20640 22250 20668 22646
rect 20548 22234 20668 22250
rect 20536 22228 20668 22234
rect 20588 22222 20668 22228
rect 20536 22170 20588 22176
rect 20824 22094 20852 22918
rect 20824 22066 20944 22094
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20602 20760 20878
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18970 20852 19246
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20640 18426 20668 18634
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20272 15558 20484 15586
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14550 19656 14758
rect 19616 14544 19668 14550
rect 20272 14498 20300 15558
rect 20548 15026 20576 15642
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20640 15026 20668 15574
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 19616 14486 19668 14492
rect 20180 14470 20300 14498
rect 19616 14408 19668 14414
rect 19536 14368 19616 14396
rect 19352 14334 19472 14362
rect 19984 14408 20036 14414
rect 19668 14368 19984 14396
rect 19616 14350 19668 14356
rect 19984 14350 20036 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19352 13394 19380 14334
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12374 19380 13126
rect 19444 12986 19472 14214
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19536 12753 19564 12786
rect 19522 12744 19578 12753
rect 19522 12679 19578 12688
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11626 19380 12038
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19444 11234 19472 12242
rect 19536 12238 19564 12582
rect 19996 12458 20024 14350
rect 20088 14006 20116 14350
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20180 12986 20208 14470
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20272 13258 20300 14214
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20272 12850 20300 13194
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19904 12430 20024 12458
rect 19904 12238 19932 12430
rect 20088 12345 20116 12718
rect 20074 12336 20130 12345
rect 20074 12271 20130 12280
rect 19524 12232 19576 12238
rect 19708 12232 19760 12238
rect 19524 12174 19576 12180
rect 19706 12200 19708 12209
rect 19892 12232 19944 12238
rect 19760 12200 19762 12209
rect 19892 12174 19944 12180
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19706 12135 19762 12144
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19524 11892 19576 11898
rect 19576 11852 19656 11880
rect 19524 11834 19576 11840
rect 19628 11529 19656 11852
rect 19996 11778 20024 12174
rect 20168 12096 20220 12102
rect 20074 12064 20130 12073
rect 20168 12038 20220 12044
rect 20074 11999 20130 12008
rect 20088 11898 20116 11999
rect 20180 11898 20208 12038
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 19708 11756 19760 11762
rect 19996 11750 20116 11778
rect 19708 11698 19760 11704
rect 19720 11665 19748 11698
rect 19706 11656 19762 11665
rect 19706 11591 19762 11600
rect 19984 11552 20036 11558
rect 19614 11520 19670 11529
rect 19984 11494 20036 11500
rect 19614 11455 19670 11464
rect 19444 11206 19656 11234
rect 19628 11150 19656 11206
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19352 10810 19380 11086
rect 19536 10996 19564 11086
rect 19444 10968 19564 10996
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19352 9636 19380 10474
rect 19444 10198 19472 10968
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10198 20024 11494
rect 20088 10266 20116 11750
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19432 10192 19484 10198
rect 19430 10160 19432 10169
rect 19984 10192 20036 10198
rect 19484 10160 19486 10169
rect 19984 10134 20036 10140
rect 19430 10095 19486 10104
rect 19984 9920 20036 9926
rect 20036 9880 20116 9908
rect 19984 9862 20036 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19616 9716 19668 9722
rect 19522 9688 19578 9697
rect 19352 9608 19472 9636
rect 19616 9658 19668 9664
rect 19800 9716 19852 9722
rect 20088 9704 20116 9880
rect 19996 9676 20116 9704
rect 19852 9664 19932 9674
rect 19800 9658 19932 9664
rect 19522 9623 19578 9632
rect 19340 9512 19392 9518
rect 19444 9500 19472 9608
rect 19392 9472 19472 9500
rect 19340 9454 19392 9460
rect 19340 9376 19392 9382
rect 19260 9336 19340 9364
rect 19156 9318 19208 9324
rect 19340 9318 19392 9324
rect 19338 9208 19394 9217
rect 19338 9143 19394 9152
rect 19352 7818 19380 9143
rect 19444 7954 19472 9472
rect 19536 8974 19564 9623
rect 19628 9353 19656 9658
rect 19812 9646 19932 9658
rect 19614 9344 19670 9353
rect 19614 9279 19670 9288
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19904 8888 19932 9646
rect 19996 9586 20024 9676
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20076 9512 20128 9518
rect 19982 9480 20038 9489
rect 20038 9460 20076 9466
rect 20038 9454 20128 9460
rect 20038 9438 20116 9454
rect 19982 9415 20038 9424
rect 19996 9042 20024 9415
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 9217 20116 9318
rect 20074 9208 20130 9217
rect 20074 9143 20130 9152
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 20076 8900 20128 8906
rect 19904 8860 20024 8888
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19062 6352 19118 6361
rect 19168 6322 19196 6598
rect 19062 6287 19118 6296
rect 19156 6316 19208 6322
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 19076 6186 19104 6287
rect 19156 6258 19208 6264
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 19260 5914 19288 6734
rect 19352 6322 19380 7414
rect 19444 6390 19472 7890
rect 19536 7750 19564 8026
rect 19628 8022 19656 8366
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19904 7954 19932 8502
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7546 20024 8860
rect 20076 8842 20128 8848
rect 20088 8634 20116 8842
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20088 8090 20116 8570
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19996 7426 20024 7482
rect 19904 7398 20024 7426
rect 19904 6866 19932 7398
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19996 6322 20024 7278
rect 20180 7206 20208 11698
rect 20272 7410 20300 12174
rect 20364 10198 20392 14758
rect 20456 14618 20484 14758
rect 20444 14612 20496 14618
rect 20640 14600 20668 14962
rect 20732 14890 20760 15438
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20824 15162 20852 15370
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20824 14822 20852 14962
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20812 14612 20864 14618
rect 20640 14572 20760 14600
rect 20444 14554 20496 14560
rect 20444 14408 20496 14414
rect 20732 14362 20760 14572
rect 20916 14600 20944 22066
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21468 20602 21496 21490
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21284 19922 21312 20538
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21088 19304 21140 19310
rect 21192 19281 21220 19382
rect 21088 19246 21140 19252
rect 21178 19272 21234 19281
rect 21100 18766 21128 19246
rect 21178 19207 21234 19216
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 18970 21496 19178
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 21560 18426 21588 19654
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18902 21680 19110
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21744 18426 21772 20334
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21836 18358 21864 19314
rect 21928 19281 21956 19790
rect 21914 19272 21970 19281
rect 21914 19207 21970 19216
rect 21928 18902 21956 19207
rect 21916 18896 21968 18902
rect 21916 18838 21968 18844
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21100 15706 21128 16050
rect 21192 15706 21220 18158
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21928 17746 21956 18090
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 17134 21864 17478
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21638 15600 21694 15609
rect 21744 15570 21772 15846
rect 21836 15638 21864 15914
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21638 15535 21640 15544
rect 21692 15535 21694 15544
rect 21732 15564 21784 15570
rect 21640 15506 21692 15512
rect 21732 15506 21784 15512
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20864 14572 20944 14600
rect 20812 14554 20864 14560
rect 20444 14350 20496 14356
rect 20456 14074 20484 14350
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20640 14334 20760 14362
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 12850 20576 14282
rect 20640 13190 20668 14334
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 11898 20484 12650
rect 20548 12646 20576 12786
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20536 12232 20588 12238
rect 20640 12209 20668 12310
rect 20536 12174 20588 12180
rect 20626 12200 20682 12209
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 11393 20484 11698
rect 20442 11384 20498 11393
rect 20442 11319 20498 11328
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20456 10146 20484 11319
rect 20548 10810 20576 12174
rect 20626 12135 20682 12144
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11830 20668 12038
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20640 11665 20668 11766
rect 20732 11762 20760 13874
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20824 12850 20852 13262
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20824 12238 20852 12786
rect 20916 12442 20944 12786
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20626 11656 20682 11665
rect 20626 11591 20682 11600
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20456 10118 20668 10146
rect 20352 10056 20404 10062
rect 20350 10024 20352 10033
rect 20444 10058 20496 10064
rect 20404 10024 20406 10033
rect 20444 10000 20496 10006
rect 20350 9959 20406 9968
rect 20350 9888 20406 9897
rect 20350 9823 20406 9832
rect 20364 9178 20392 9823
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20350 8256 20406 8265
rect 20350 8191 20406 8200
rect 20364 7750 20392 8191
rect 20456 7886 20484 10000
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9722 20576 9862
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 8906 20576 9318
rect 20640 8974 20668 10118
rect 20824 10062 20852 12174
rect 21008 11801 21036 14962
rect 21836 14482 21864 15370
rect 21928 15094 21956 15438
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 20994 11792 21050 11801
rect 20994 11727 21050 11736
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20732 9897 20760 9998
rect 20718 9888 20774 9897
rect 20718 9823 20774 9832
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20640 8566 20668 8910
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20364 7478 20392 7686
rect 20548 7546 20576 7686
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17590 5672 17646 5681
rect 17408 5636 17460 5642
rect 17590 5607 17592 5616
rect 17408 5578 17460 5584
rect 17644 5607 17646 5616
rect 17592 5578 17644 5584
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13740 3194 13768 3470
rect 14568 3194 14596 3878
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 14844 2990 14872 3946
rect 16132 3534 16160 4490
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 4146 16620 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16316 3738 16344 4082
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16868 3602 16896 4490
rect 17420 3942 17448 5578
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16132 2990 16160 3334
rect 17420 3126 17448 3878
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17604 3176 17632 3470
rect 17972 3398 18000 4558
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18064 3602 18092 4014
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18156 3534 18184 5034
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18708 3942 18736 4694
rect 19168 4622 19196 5102
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 4214 18828 4422
rect 19168 4282 19196 4558
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 19444 3992 19472 6054
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5386 20024 6258
rect 19996 5370 20116 5386
rect 19996 5364 20128 5370
rect 19996 5358 20076 5364
rect 20076 5306 20128 5312
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 19996 4486 20024 5238
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4146 20024 4422
rect 20180 4282 20208 7142
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20272 6458 20300 6734
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20456 6390 20484 6734
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 20824 5914 20852 9998
rect 21008 9926 21036 11727
rect 21192 11694 21220 12378
rect 21376 12306 21404 12650
rect 21744 12374 21772 14282
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12986 21956 13330
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 22020 8634 22048 19858
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22112 17882 22140 18226
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22204 16130 22232 23174
rect 22388 22778 22416 23258
rect 22480 23186 22508 23598
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22778 22508 22918
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22468 22568 22520 22574
rect 22468 22510 22520 22516
rect 22296 16250 22324 22510
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22388 22030 22416 22442
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22480 20398 22508 22510
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22388 19446 22416 20334
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22480 19174 22508 19654
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22480 18714 22508 19110
rect 22388 18686 22508 18714
rect 22560 18692 22612 18698
rect 22388 18630 22416 18686
rect 22560 18634 22612 18640
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 18057 22508 18566
rect 22466 18048 22522 18057
rect 22466 17983 22522 17992
rect 22572 17678 22600 18634
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22664 17626 22692 23054
rect 22756 22778 22784 23666
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22940 22094 22968 25894
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23584 24954 23612 25842
rect 23756 25696 23808 25702
rect 23756 25638 23808 25644
rect 23768 25362 23796 25638
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 23526 23428 24142
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 23032 22574 23060 23122
rect 23400 23118 23428 23462
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23124 22098 23152 22510
rect 22848 22066 22968 22094
rect 23112 22092 23164 22098
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20602 22784 20742
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22756 18426 22784 18770
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22756 17746 22784 18362
rect 22744 17740 22796 17746
rect 22744 17682 22796 17688
rect 22664 17598 22784 17626
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22388 16250 22416 17138
rect 22664 16697 22692 17478
rect 22650 16688 22706 16697
rect 22650 16623 22706 16632
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22204 16102 22324 16130
rect 22100 15496 22152 15502
rect 22098 15464 22100 15473
rect 22152 15464 22154 15473
rect 22098 15399 22154 15408
rect 22296 13462 22324 16102
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15745 22416 16050
rect 22374 15736 22430 15745
rect 22374 15671 22430 15680
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22388 15008 22416 15506
rect 22480 15502 22508 15642
rect 22756 15638 22784 17598
rect 22744 15632 22796 15638
rect 22744 15574 22796 15580
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22652 15496 22704 15502
rect 22742 15464 22798 15473
rect 22704 15444 22742 15450
rect 22652 15438 22742 15444
rect 22572 15162 22600 15438
rect 22664 15422 22742 15438
rect 22742 15399 22798 15408
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 15162 22784 15302
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22468 15020 22520 15026
rect 22388 14980 22468 15008
rect 22468 14962 22520 14968
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22112 12986 22140 13262
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 8090 21864 8366
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 22112 7886 22140 10406
rect 22204 9926 22232 13194
rect 22388 12889 22416 13262
rect 22374 12880 22430 12889
rect 22374 12815 22430 12824
rect 22480 12646 22508 14962
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14618 22600 14758
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22650 13832 22706 13841
rect 22650 13767 22706 13776
rect 22664 13394 22692 13767
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22204 9586 22232 9862
rect 22388 9654 22416 11086
rect 22480 10674 22508 12582
rect 22848 12442 22876 22066
rect 23952 22094 23980 28494
rect 24228 28218 24256 28630
rect 24412 28558 24440 29514
rect 24780 29102 24808 30670
rect 25044 30592 25096 30598
rect 25044 30534 25096 30540
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24872 29306 24900 29582
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 25056 29238 25084 30534
rect 25044 29232 25096 29238
rect 25044 29174 25096 29180
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 24780 28506 24808 29038
rect 24860 28552 24912 28558
rect 24780 28500 24860 28506
rect 24780 28494 24912 28500
rect 24780 28478 24900 28494
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24688 27538 24716 27950
rect 24676 27532 24728 27538
rect 24676 27474 24728 27480
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24412 27130 24440 27270
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24596 26874 24624 27406
rect 24780 27062 24808 28478
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24124 26852 24176 26858
rect 24596 26846 24808 26874
rect 24124 26794 24176 26800
rect 24136 26382 24164 26794
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24044 26042 24072 26318
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 24136 25362 24164 26318
rect 24676 26308 24728 26314
rect 24676 26250 24728 26256
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24688 25226 24716 26250
rect 24780 25838 24808 26846
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24780 25362 24808 25774
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24688 24410 24716 24754
rect 24780 24750 24808 25298
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22778 24808 23054
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 23952 22066 24072 22094
rect 23112 22034 23164 22040
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21690 23244 21966
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23216 21010 23244 21626
rect 23676 21486 23704 21830
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23308 21146 23336 21286
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 23308 20466 23336 21082
rect 23400 20942 23428 21422
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23204 19440 23256 19446
rect 23204 19382 23256 19388
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23032 18426 23060 18634
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23216 17354 23244 19382
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23400 18834 23428 19314
rect 23584 18970 23612 19314
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23676 18834 23704 20946
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23768 20602 23796 20742
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23952 19514 23980 19722
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23400 18290 23428 18566
rect 23768 18426 23796 18566
rect 23952 18426 23980 19450
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23216 17326 23336 17354
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22940 16250 22968 17002
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 23020 16176 23072 16182
rect 23124 16164 23152 16526
rect 23216 16250 23244 17206
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23072 16136 23152 16164
rect 23020 16118 23072 16124
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 23020 15972 23072 15978
rect 23020 15914 23072 15920
rect 22940 15366 22968 15914
rect 23032 15706 23060 15914
rect 23124 15706 23152 16136
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 23032 13394 23060 15438
rect 23216 15026 23244 16050
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23216 14618 23244 14962
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22558 10976 22614 10985
rect 22558 10911 22614 10920
rect 22572 10810 22600 10911
rect 22664 10810 22692 11086
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22756 10266 22784 12038
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 10266 22876 10406
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22558 10024 22614 10033
rect 22558 9959 22560 9968
rect 22612 9959 22614 9968
rect 22560 9930 22612 9936
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22558 9616 22614 9625
rect 22192 9580 22244 9586
rect 22756 9586 22784 10202
rect 22558 9551 22614 9560
rect 22744 9580 22796 9586
rect 22192 9522 22244 9528
rect 22204 8906 22232 9522
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 9178 22508 9318
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22572 9110 22600 9551
rect 22744 9522 22796 9528
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22204 8430 22232 8842
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21100 7002 21128 7278
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21192 6798 21220 7210
rect 21468 7002 21496 7754
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20824 5166 20852 5850
rect 21192 5710 21220 6734
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4826 20392 4966
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20824 4690 20852 5102
rect 21284 4826 21312 5102
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 21560 4622 21588 7754
rect 22112 7410 22140 7822
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22204 5234 22232 8366
rect 22296 8294 22324 8910
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22940 7546 22968 12174
rect 23032 10742 23060 12786
rect 23216 12730 23244 12922
rect 23124 12702 23244 12730
rect 23124 12306 23152 12702
rect 23308 12628 23336 17326
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 16114 23428 16594
rect 23492 16590 23520 18022
rect 23952 17746 23980 18362
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23584 16182 23612 16526
rect 23676 16454 23704 17682
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23480 15496 23532 15502
rect 23386 15464 23442 15473
rect 23480 15438 23532 15444
rect 23386 15399 23388 15408
rect 23440 15399 23442 15408
rect 23388 15370 23440 15376
rect 23492 15094 23520 15438
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23400 12782 23428 14554
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23216 12600 23336 12628
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23216 11354 23244 12600
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23020 10736 23072 10742
rect 23020 10678 23072 10684
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 8974 23060 9318
rect 23216 8974 23244 11154
rect 23400 11082 23428 12718
rect 23584 11898 23612 15982
rect 23768 15978 23796 17546
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23676 15162 23704 15846
rect 24044 15706 24072 22066
rect 24136 16674 24164 22578
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24320 21486 24348 22374
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24780 21146 24808 22102
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20602 24256 20742
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24412 19786 24440 20878
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24688 20602 24716 20810
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24400 19780 24452 19786
rect 24400 19722 24452 19728
rect 24492 18896 24544 18902
rect 24320 18856 24492 18884
rect 24320 18850 24348 18856
rect 24228 18834 24348 18850
rect 24492 18838 24544 18844
rect 24216 18828 24348 18834
rect 24268 18822 24348 18828
rect 24216 18770 24268 18776
rect 24136 16646 24440 16674
rect 24122 15736 24178 15745
rect 24032 15700 24084 15706
rect 24308 15700 24360 15706
rect 24178 15680 24308 15688
rect 24122 15671 24308 15680
rect 24136 15660 24308 15671
rect 24032 15642 24084 15648
rect 24308 15642 24360 15648
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 23756 15496 23808 15502
rect 23808 15456 23980 15484
rect 23756 15438 23808 15444
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 12918 23796 14758
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23860 12850 23888 15302
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23860 12594 23888 12786
rect 23768 12566 23888 12594
rect 23768 12306 23796 12566
rect 23952 12434 23980 15456
rect 24136 15366 24164 15506
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24136 13462 24164 13738
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 24320 12850 24348 14010
rect 24412 13326 24440 16646
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24504 16046 24532 16526
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24504 15910 24532 15982
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24504 15434 24532 15846
rect 24688 15706 24716 16050
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24492 15428 24544 15434
rect 24676 15428 24728 15434
rect 24544 15388 24676 15416
rect 24492 15370 24544 15376
rect 24676 15370 24728 15376
rect 24688 13938 24716 15370
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 23860 12406 23980 12434
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23020 8968 23072 8974
rect 23204 8968 23256 8974
rect 23020 8910 23072 8916
rect 23124 8928 23204 8956
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22112 4690 22140 5102
rect 23124 5098 23152 8928
rect 23204 8910 23256 8916
rect 23308 8514 23336 10678
rect 23400 9586 23428 11018
rect 23768 10742 23796 12242
rect 23756 10736 23808 10742
rect 23756 10678 23808 10684
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23492 9722 23520 10542
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23400 9178 23428 9522
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 8634 23428 8774
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23308 8486 23428 8514
rect 23400 8362 23428 8486
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23294 8120 23350 8129
rect 23294 8055 23296 8064
rect 23348 8055 23350 8064
rect 23296 8026 23348 8032
rect 23308 5166 23336 8026
rect 23400 7206 23428 8298
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23492 6662 23520 9658
rect 23584 9654 23612 10610
rect 23676 9722 23704 10610
rect 23860 10130 23888 12406
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23952 10742 23980 11834
rect 24044 10810 24072 12786
rect 24412 12714 24440 13262
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 24492 12708 24544 12714
rect 24492 12650 24544 12656
rect 24504 11150 24532 12650
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23768 8906 23796 9522
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23952 8090 23980 9522
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24412 8634 24440 8910
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23860 7478 23888 7822
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23584 7002 23612 7278
rect 23860 7002 23888 7414
rect 24412 7342 24440 7686
rect 24596 7546 24624 13806
rect 24688 11218 24716 13874
rect 24780 11694 24808 15982
rect 24872 14074 24900 27950
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24964 24954 24992 25162
rect 24952 24948 25004 24954
rect 24952 24890 25004 24896
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24964 23186 24992 24550
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 25056 18884 25084 27270
rect 25332 24274 25360 40598
rect 25516 38350 25544 42502
rect 26160 42226 26188 42502
rect 26712 42362 26740 42502
rect 26700 42356 26752 42362
rect 26700 42298 26752 42304
rect 26332 42288 26384 42294
rect 26332 42230 26384 42236
rect 26148 42220 26200 42226
rect 26148 42162 26200 42168
rect 26148 41472 26200 41478
rect 26148 41414 26200 41420
rect 26160 40526 26188 41414
rect 26344 41256 26372 42230
rect 26700 42220 26752 42226
rect 26700 42162 26752 42168
rect 26712 42129 26740 42162
rect 26698 42120 26754 42129
rect 26804 42090 26832 43250
rect 26896 42294 26924 43250
rect 26976 43104 27028 43110
rect 26976 43046 27028 43052
rect 26884 42288 26936 42294
rect 26884 42230 26936 42236
rect 26698 42055 26754 42064
rect 26792 42084 26844 42090
rect 26792 42026 26844 42032
rect 26700 42016 26752 42022
rect 26700 41958 26752 41964
rect 26712 41818 26740 41958
rect 26700 41812 26752 41818
rect 26700 41754 26752 41760
rect 26252 41228 26372 41256
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 26252 40186 26280 41228
rect 26804 41206 26832 42026
rect 26988 41614 27016 43046
rect 27252 42152 27304 42158
rect 27252 42094 27304 42100
rect 27264 41818 27292 42094
rect 27252 41812 27304 41818
rect 27252 41754 27304 41760
rect 26976 41608 27028 41614
rect 26976 41550 27028 41556
rect 27252 41540 27304 41546
rect 27252 41482 27304 41488
rect 26792 41200 26844 41206
rect 26792 41142 26844 41148
rect 27264 41138 27292 41482
rect 26332 41132 26384 41138
rect 26332 41074 26384 41080
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 26344 40458 26372 41074
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 27160 40928 27212 40934
rect 27160 40870 27212 40876
rect 26528 40594 26556 40870
rect 26884 40656 26936 40662
rect 27172 40610 27200 40870
rect 26936 40604 27200 40610
rect 26884 40598 27200 40604
rect 26516 40588 26568 40594
rect 26896 40582 27200 40598
rect 26516 40530 26568 40536
rect 26332 40452 26384 40458
rect 26332 40394 26384 40400
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 25688 39296 25740 39302
rect 25688 39238 25740 39244
rect 25700 38418 25728 39238
rect 26252 38978 26280 40122
rect 26344 39846 26372 40394
rect 26792 40384 26844 40390
rect 26792 40326 26844 40332
rect 26884 40384 26936 40390
rect 26884 40326 26936 40332
rect 26332 39840 26384 39846
rect 26332 39782 26384 39788
rect 26516 39840 26568 39846
rect 26516 39782 26568 39788
rect 26424 39432 26476 39438
rect 26424 39374 26476 39380
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26344 39098 26372 39238
rect 26436 39098 26464 39374
rect 26332 39092 26384 39098
rect 26332 39034 26384 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 26252 38950 26372 38978
rect 26240 38752 26292 38758
rect 26240 38694 26292 38700
rect 25688 38412 25740 38418
rect 25688 38354 25740 38360
rect 26056 38412 26108 38418
rect 26056 38354 26108 38360
rect 25504 38344 25556 38350
rect 25504 38286 25556 38292
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25516 37874 25544 38150
rect 25504 37868 25556 37874
rect 25504 37810 25556 37816
rect 25516 36786 25544 37810
rect 25688 37664 25740 37670
rect 25688 37606 25740 37612
rect 25700 37330 25728 37606
rect 26068 37330 26096 38354
rect 25688 37324 25740 37330
rect 25688 37266 25740 37272
rect 26056 37324 26108 37330
rect 26056 37266 26108 37272
rect 26068 37194 26096 37266
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25792 35834 25820 36110
rect 25780 35828 25832 35834
rect 25780 35770 25832 35776
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25884 35154 25912 35430
rect 25872 35148 25924 35154
rect 25872 35090 25924 35096
rect 26068 34950 26096 37130
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 26160 35290 26188 36654
rect 26148 35284 26200 35290
rect 26148 35226 26200 35232
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 26252 34610 26280 38694
rect 26344 36174 26372 38950
rect 26528 38826 26556 39782
rect 26804 39506 26832 40326
rect 26896 39982 26924 40326
rect 27172 40050 27200 40582
rect 27344 40520 27396 40526
rect 27344 40462 27396 40468
rect 27356 40050 27384 40462
rect 27436 40384 27488 40390
rect 27436 40326 27488 40332
rect 27448 40186 27476 40326
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 27620 40112 27672 40118
rect 27620 40054 27672 40060
rect 27160 40044 27212 40050
rect 27160 39986 27212 39992
rect 27344 40044 27396 40050
rect 27344 39986 27396 39992
rect 26884 39976 26936 39982
rect 26884 39918 26936 39924
rect 27528 39908 27580 39914
rect 27528 39850 27580 39856
rect 27540 39642 27568 39850
rect 27528 39636 27580 39642
rect 27528 39578 27580 39584
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 27540 38962 27568 39578
rect 27632 39098 27660 40054
rect 27620 39092 27672 39098
rect 27620 39034 27672 39040
rect 27528 38956 27580 38962
rect 27528 38898 27580 38904
rect 26516 38820 26568 38826
rect 26516 38762 26568 38768
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 27528 38208 27580 38214
rect 27528 38150 27580 38156
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26436 35034 26464 38150
rect 27540 37466 27568 38150
rect 27528 37460 27580 37466
rect 27528 37402 27580 37408
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 27080 37233 27108 37266
rect 27066 37224 27122 37233
rect 27066 37159 27122 37168
rect 27436 37188 27488 37194
rect 27080 36854 27108 37159
rect 27436 37130 27488 37136
rect 27448 36922 27476 37130
rect 27436 36916 27488 36922
rect 27436 36858 27488 36864
rect 27068 36848 27120 36854
rect 27068 36790 27120 36796
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27356 36310 27384 36722
rect 27344 36304 27396 36310
rect 27342 36272 27344 36281
rect 27396 36272 27398 36281
rect 27342 36207 27398 36216
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27632 35698 27660 36042
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27620 35556 27672 35562
rect 27620 35498 27672 35504
rect 26436 35006 26648 35034
rect 26436 34678 26464 35006
rect 26620 34950 26648 35006
rect 26516 34944 26568 34950
rect 26516 34886 26568 34892
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26424 34672 26476 34678
rect 26424 34614 26476 34620
rect 26528 34610 26556 34886
rect 27632 34610 27660 35498
rect 27724 35034 27752 43590
rect 28552 42906 28580 43590
rect 29932 43450 29960 43794
rect 30840 43716 30892 43722
rect 30840 43658 30892 43664
rect 29920 43444 29972 43450
rect 29920 43386 29972 43392
rect 28540 42900 28592 42906
rect 28540 42842 28592 42848
rect 27988 42628 28040 42634
rect 27988 42570 28040 42576
rect 27804 40588 27856 40594
rect 27804 40530 27856 40536
rect 27816 38758 27844 40530
rect 27896 40044 27948 40050
rect 27896 39986 27948 39992
rect 27908 39642 27936 39986
rect 27896 39636 27948 39642
rect 27896 39578 27948 39584
rect 27804 38752 27856 38758
rect 27804 38694 27856 38700
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27816 36582 27844 37742
rect 28000 36854 28028 42570
rect 28552 42294 28580 42842
rect 30012 42628 30064 42634
rect 30012 42570 30064 42576
rect 28540 42288 28592 42294
rect 28540 42230 28592 42236
rect 29092 42152 29144 42158
rect 28814 42120 28870 42129
rect 29092 42094 29144 42100
rect 28814 42055 28870 42064
rect 28356 42016 28408 42022
rect 28356 41958 28408 41964
rect 28368 41682 28396 41958
rect 28356 41676 28408 41682
rect 28356 41618 28408 41624
rect 28368 41414 28396 41618
rect 28276 41386 28396 41414
rect 28276 41274 28304 41386
rect 28264 41268 28316 41274
rect 28264 41210 28316 41216
rect 28368 40934 28396 41386
rect 28828 41206 28856 42055
rect 29104 41818 29132 42094
rect 29092 41812 29144 41818
rect 29092 41754 29144 41760
rect 29828 41812 29880 41818
rect 29828 41754 29880 41760
rect 29840 41546 29868 41754
rect 29828 41540 29880 41546
rect 29828 41482 29880 41488
rect 29644 41472 29696 41478
rect 29644 41414 29696 41420
rect 29656 41313 29684 41414
rect 29642 41304 29698 41313
rect 29642 41239 29698 41248
rect 28816 41200 28868 41206
rect 28816 41142 28868 41148
rect 28264 40928 28316 40934
rect 28264 40870 28316 40876
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 28540 40928 28592 40934
rect 28540 40870 28592 40876
rect 28276 40526 28304 40870
rect 28552 40730 28580 40870
rect 28540 40724 28592 40730
rect 28540 40666 28592 40672
rect 28264 40520 28316 40526
rect 28264 40462 28316 40468
rect 28276 40186 28304 40462
rect 28172 40180 28224 40186
rect 28172 40122 28224 40128
rect 28264 40180 28316 40186
rect 28264 40122 28316 40128
rect 28184 38962 28212 40122
rect 28264 39976 28316 39982
rect 28264 39918 28316 39924
rect 28276 39098 28304 39918
rect 28264 39092 28316 39098
rect 28264 39034 28316 39040
rect 28172 38956 28224 38962
rect 28172 38898 28224 38904
rect 28908 38956 28960 38962
rect 28908 38898 28960 38904
rect 28920 37466 28948 38898
rect 29656 38282 29684 41239
rect 30024 39506 30052 42570
rect 30380 42560 30432 42566
rect 30380 42502 30432 42508
rect 30656 42560 30708 42566
rect 30656 42502 30708 42508
rect 30748 42560 30800 42566
rect 30748 42502 30800 42508
rect 30392 42294 30420 42502
rect 30380 42288 30432 42294
rect 30380 42230 30432 42236
rect 30564 42288 30616 42294
rect 30564 42230 30616 42236
rect 30196 42084 30248 42090
rect 30196 42026 30248 42032
rect 30472 42084 30524 42090
rect 30472 42026 30524 42032
rect 30102 41712 30158 41721
rect 30102 41647 30104 41656
rect 30156 41647 30158 41656
rect 30104 41618 30156 41624
rect 30012 39500 30064 39506
rect 29932 39460 30012 39488
rect 29828 39432 29880 39438
rect 29828 39374 29880 39380
rect 29840 39098 29868 39374
rect 29828 39092 29880 39098
rect 29828 39034 29880 39040
rect 29932 39030 29960 39460
rect 30012 39442 30064 39448
rect 30208 39438 30236 42026
rect 30484 41818 30512 42026
rect 30380 41812 30432 41818
rect 30380 41754 30432 41760
rect 30472 41812 30524 41818
rect 30472 41754 30524 41760
rect 30288 41608 30340 41614
rect 30288 41550 30340 41556
rect 30300 41274 30328 41550
rect 30392 41478 30420 41754
rect 30472 41540 30524 41546
rect 30576 41528 30604 42230
rect 30668 42226 30696 42502
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 30656 42016 30708 42022
rect 30656 41958 30708 41964
rect 30668 41818 30696 41958
rect 30656 41812 30708 41818
rect 30656 41754 30708 41760
rect 30760 41698 30788 42502
rect 30852 41818 30880 43658
rect 31668 43104 31720 43110
rect 31668 43046 31720 43052
rect 31024 42696 31076 42702
rect 31024 42638 31076 42644
rect 30840 41812 30892 41818
rect 30840 41754 30892 41760
rect 30668 41670 30788 41698
rect 30932 41676 30984 41682
rect 30668 41546 30696 41670
rect 30932 41618 30984 41624
rect 30748 41608 30800 41614
rect 30748 41550 30800 41556
rect 30524 41500 30604 41528
rect 30656 41540 30708 41546
rect 30472 41482 30524 41488
rect 30656 41482 30708 41488
rect 30380 41472 30432 41478
rect 30380 41414 30432 41420
rect 30288 41268 30340 41274
rect 30288 41210 30340 41216
rect 30564 41064 30616 41070
rect 30760 41052 30788 41550
rect 30944 41414 30972 41618
rect 30852 41386 30972 41414
rect 30852 41274 30880 41386
rect 31036 41290 31064 42638
rect 31680 42362 31708 43046
rect 31864 42702 31892 43794
rect 31944 43648 31996 43654
rect 31944 43590 31996 43596
rect 31956 42906 31984 43590
rect 31944 42900 31996 42906
rect 31944 42842 31996 42848
rect 31944 42764 31996 42770
rect 31944 42706 31996 42712
rect 31852 42696 31904 42702
rect 31852 42638 31904 42644
rect 31760 42560 31812 42566
rect 31760 42502 31812 42508
rect 31772 42362 31800 42502
rect 31484 42356 31536 42362
rect 31484 42298 31536 42304
rect 31668 42356 31720 42362
rect 31668 42298 31720 42304
rect 31760 42356 31812 42362
rect 31760 42298 31812 42304
rect 31208 42016 31260 42022
rect 31208 41958 31260 41964
rect 31220 41614 31248 41958
rect 31208 41608 31260 41614
rect 31208 41550 31260 41556
rect 30840 41268 30892 41274
rect 30840 41210 30892 41216
rect 30944 41262 31064 41290
rect 30944 41206 30972 41262
rect 30932 41200 30984 41206
rect 30932 41142 30984 41148
rect 31220 41138 31248 41550
rect 31392 41540 31444 41546
rect 31392 41482 31444 41488
rect 31208 41132 31260 41138
rect 31260 41092 31340 41120
rect 31208 41074 31260 41080
rect 30616 41024 30788 41052
rect 30564 41006 30616 41012
rect 30288 40928 30340 40934
rect 30288 40870 30340 40876
rect 30300 39846 30328 40870
rect 30760 40458 30788 41024
rect 30932 41064 30984 41070
rect 31116 41064 31168 41070
rect 30932 41006 30984 41012
rect 31114 41032 31116 41041
rect 31168 41032 31170 41041
rect 30748 40452 30800 40458
rect 30748 40394 30800 40400
rect 30944 40118 30972 41006
rect 31114 40967 31170 40976
rect 31208 40928 31260 40934
rect 31208 40870 31260 40876
rect 30932 40112 30984 40118
rect 30932 40054 30984 40060
rect 30288 39840 30340 39846
rect 30288 39782 30340 39788
rect 30300 39658 30328 39782
rect 30300 39630 30604 39658
rect 30288 39568 30340 39574
rect 30288 39510 30340 39516
rect 30196 39432 30248 39438
rect 30196 39374 30248 39380
rect 30012 39296 30064 39302
rect 30012 39238 30064 39244
rect 30024 39098 30052 39238
rect 30012 39092 30064 39098
rect 30208 39080 30236 39374
rect 30012 39034 30064 39040
rect 30116 39052 30236 39080
rect 29920 39024 29972 39030
rect 29920 38966 29972 38972
rect 30116 38962 30144 39052
rect 30104 38956 30156 38962
rect 30104 38898 30156 38904
rect 29736 38752 29788 38758
rect 29736 38694 29788 38700
rect 29748 38350 29776 38694
rect 29736 38344 29788 38350
rect 29736 38286 29788 38292
rect 30012 38344 30064 38350
rect 30064 38304 30144 38332
rect 30012 38286 30064 38292
rect 29368 38276 29420 38282
rect 29368 38218 29420 38224
rect 29644 38276 29696 38282
rect 29644 38218 29696 38224
rect 29092 38208 29144 38214
rect 29092 38150 29144 38156
rect 29104 38010 29132 38150
rect 29092 38004 29144 38010
rect 29092 37946 29144 37952
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 28908 37460 28960 37466
rect 28908 37402 28960 37408
rect 29104 37126 29132 37742
rect 29092 37120 29144 37126
rect 29092 37062 29144 37068
rect 27988 36848 28040 36854
rect 27988 36790 28040 36796
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 27816 36242 27844 36518
rect 27804 36236 27856 36242
rect 27804 36178 27856 36184
rect 27816 35154 27844 36178
rect 27804 35148 27856 35154
rect 27804 35090 27856 35096
rect 27724 35006 27844 35034
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 26516 34604 26568 34610
rect 26516 34546 26568 34552
rect 27620 34604 27672 34610
rect 27620 34546 27672 34552
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33658 27568 33798
rect 27528 33652 27580 33658
rect 27528 33594 27580 33600
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 26344 32978 26372 33458
rect 27724 33114 27752 33458
rect 27712 33108 27764 33114
rect 27712 33050 27764 33056
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26608 32972 26660 32978
rect 26608 32914 26660 32920
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 32570 26096 32846
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 25964 32360 26016 32366
rect 25964 32302 26016 32308
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25516 29510 25544 31758
rect 25976 31482 26004 32302
rect 26344 31890 26372 32914
rect 26516 32224 26568 32230
rect 26516 32166 26568 32172
rect 26424 31952 26476 31958
rect 26424 31894 26476 31900
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 26252 31278 26280 31758
rect 26332 31680 26384 31686
rect 26332 31622 26384 31628
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 26344 30734 26372 31622
rect 26436 31498 26464 31894
rect 26528 31822 26556 32166
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26436 31470 26556 31498
rect 26528 31278 26556 31470
rect 26620 31362 26648 32914
rect 27344 32768 27396 32774
rect 27344 32710 27396 32716
rect 27356 32570 27384 32710
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27436 32360 27488 32366
rect 27436 32302 27488 32308
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 26712 31482 26740 31758
rect 26700 31476 26752 31482
rect 26700 31418 26752 31424
rect 26620 31346 26832 31362
rect 26620 31340 26844 31346
rect 26620 31334 26792 31340
rect 26792 31282 26844 31288
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 26332 30728 26384 30734
rect 26332 30670 26384 30676
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 25424 28218 25452 28426
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25516 27470 25544 29446
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25792 27130 25820 29582
rect 26160 29034 26188 30126
rect 26148 29028 26200 29034
rect 26148 28970 26200 28976
rect 26436 28762 26464 31214
rect 26804 30938 26832 31282
rect 27068 31272 27120 31278
rect 27068 31214 27120 31220
rect 26792 30932 26844 30938
rect 26792 30874 26844 30880
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26620 28762 26648 30194
rect 26792 30048 26844 30054
rect 26792 29990 26844 29996
rect 26804 29238 26832 29990
rect 27080 29850 27108 31214
rect 27160 30728 27212 30734
rect 27160 30670 27212 30676
rect 27172 29850 27200 30670
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 27356 30326 27384 30534
rect 27344 30320 27396 30326
rect 27344 30262 27396 30268
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 26792 29232 26844 29238
rect 26792 29174 26844 29180
rect 26424 28756 26476 28762
rect 26424 28698 26476 28704
rect 26608 28756 26660 28762
rect 26608 28698 26660 28704
rect 26436 28082 26464 28698
rect 27448 28218 27476 32302
rect 27540 31210 27568 32302
rect 27712 31884 27764 31890
rect 27712 31826 27764 31832
rect 27724 31754 27752 31826
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27528 31204 27580 31210
rect 27528 31146 27580 31152
rect 27540 29782 27568 31146
rect 27724 30326 27752 31690
rect 27816 30802 27844 35006
rect 27896 35012 27948 35018
rect 27896 34954 27948 34960
rect 27908 34746 27936 34954
rect 27896 34740 27948 34746
rect 27896 34682 27948 34688
rect 28000 33998 28028 36790
rect 29000 36576 29052 36582
rect 29000 36518 29052 36524
rect 29012 36378 29040 36518
rect 29000 36372 29052 36378
rect 29000 36314 29052 36320
rect 29104 36106 29132 37062
rect 29276 36916 29328 36922
rect 29276 36858 29328 36864
rect 29288 36786 29316 36858
rect 29380 36786 29408 38218
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 30024 37262 30052 37606
rect 30012 37256 30064 37262
rect 30012 37198 30064 37204
rect 29920 37120 29972 37126
rect 29920 37062 29972 37068
rect 29932 36922 29960 37062
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 29276 36780 29328 36786
rect 29276 36722 29328 36728
rect 29368 36780 29420 36786
rect 29368 36722 29420 36728
rect 29184 36304 29236 36310
rect 29184 36246 29236 36252
rect 29092 36100 29144 36106
rect 29092 36042 29144 36048
rect 29196 36038 29224 36246
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 29380 35986 29408 36722
rect 29840 36650 29868 36858
rect 30116 36786 30144 38304
rect 30300 37126 30328 39510
rect 30380 39500 30432 39506
rect 30380 39442 30432 39448
rect 30392 38554 30420 39442
rect 30472 39296 30524 39302
rect 30472 39238 30524 39244
rect 30484 39098 30512 39238
rect 30576 39098 30604 39630
rect 30472 39092 30524 39098
rect 30472 39034 30524 39040
rect 30564 39092 30616 39098
rect 30564 39034 30616 39040
rect 30564 38752 30616 38758
rect 30564 38694 30616 38700
rect 30380 38548 30432 38554
rect 30380 38490 30432 38496
rect 30392 37874 30420 38490
rect 30576 38350 30604 38694
rect 30944 38350 30972 40054
rect 31220 38962 31248 40870
rect 31312 40730 31340 41092
rect 31404 40934 31432 41482
rect 31392 40928 31444 40934
rect 31392 40870 31444 40876
rect 31300 40724 31352 40730
rect 31300 40666 31352 40672
rect 31496 39370 31524 42298
rect 31772 42242 31800 42298
rect 31588 42214 31800 42242
rect 31852 42220 31904 42226
rect 31588 41614 31616 42214
rect 31852 42162 31904 42168
rect 31668 42152 31720 42158
rect 31668 42094 31720 42100
rect 31680 41682 31708 42094
rect 31760 42016 31812 42022
rect 31760 41958 31812 41964
rect 31668 41676 31720 41682
rect 31668 41618 31720 41624
rect 31576 41608 31628 41614
rect 31576 41550 31628 41556
rect 31588 41290 31616 41550
rect 31588 41274 31708 41290
rect 31588 41268 31720 41274
rect 31588 41262 31668 41268
rect 31668 41210 31720 41216
rect 31576 41200 31628 41206
rect 31574 41168 31576 41177
rect 31628 41168 31630 41177
rect 31574 41103 31630 41112
rect 31576 41064 31628 41070
rect 31576 41006 31628 41012
rect 31588 40594 31616 41006
rect 31772 41002 31800 41958
rect 31864 41818 31892 42162
rect 31852 41812 31904 41818
rect 31852 41754 31904 41760
rect 31864 41478 31892 41754
rect 31956 41682 31984 42706
rect 31944 41676 31996 41682
rect 31944 41618 31996 41624
rect 31852 41472 31904 41478
rect 31852 41414 31904 41420
rect 31944 41472 31996 41478
rect 31944 41414 31996 41420
rect 31956 41154 31984 41414
rect 31864 41138 31984 41154
rect 31852 41132 31984 41138
rect 31904 41126 31984 41132
rect 31852 41074 31904 41080
rect 31944 41064 31996 41070
rect 31944 41006 31996 41012
rect 31760 40996 31812 41002
rect 31760 40938 31812 40944
rect 31956 40730 31984 41006
rect 31944 40724 31996 40730
rect 31944 40666 31996 40672
rect 31576 40588 31628 40594
rect 31576 40530 31628 40536
rect 31484 39364 31536 39370
rect 31484 39306 31536 39312
rect 31208 38956 31260 38962
rect 31208 38898 31260 38904
rect 30564 38344 30616 38350
rect 30564 38286 30616 38292
rect 30840 38344 30892 38350
rect 30840 38286 30892 38292
rect 30932 38344 30984 38350
rect 30932 38286 30984 38292
rect 30380 37868 30432 37874
rect 30380 37810 30432 37816
rect 30576 37754 30604 38286
rect 30852 38010 30880 38286
rect 30840 38004 30892 38010
rect 30840 37946 30892 37952
rect 30576 37726 30788 37754
rect 30564 37664 30616 37670
rect 30564 37606 30616 37612
rect 30576 37330 30604 37606
rect 30564 37324 30616 37330
rect 30564 37266 30616 37272
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 29920 36712 29972 36718
rect 29920 36654 29972 36660
rect 29828 36644 29880 36650
rect 29828 36586 29880 36592
rect 29736 36576 29788 36582
rect 29736 36518 29788 36524
rect 29748 36174 29776 36518
rect 29932 36310 29960 36654
rect 30300 36582 30328 37062
rect 30380 36780 30432 36786
rect 30380 36722 30432 36728
rect 30392 36582 30420 36722
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 30380 36576 30432 36582
rect 30380 36518 30432 36524
rect 29920 36304 29972 36310
rect 29920 36246 29972 36252
rect 30576 36174 30604 37266
rect 30760 36786 30788 37726
rect 30840 37120 30892 37126
rect 30840 37062 30892 37068
rect 30852 36922 30880 37062
rect 30840 36916 30892 36922
rect 30840 36858 30892 36864
rect 30748 36780 30800 36786
rect 30748 36722 30800 36728
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 29828 36168 29880 36174
rect 29828 36110 29880 36116
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 28080 34944 28132 34950
rect 28080 34886 28132 34892
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 27804 30796 27856 30802
rect 27804 30738 27856 30744
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27528 29776 27580 29782
rect 27528 29718 27580 29724
rect 27540 28626 27568 29718
rect 27724 29238 27752 30262
rect 27712 29232 27764 29238
rect 27712 29174 27764 29180
rect 27528 28620 27580 28626
rect 27528 28562 27580 28568
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26976 27532 27028 27538
rect 26976 27474 27028 27480
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26436 27130 26464 27406
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26160 26246 26188 26726
rect 26988 26518 27016 27474
rect 27540 26926 27568 28562
rect 27724 27674 27752 29174
rect 27712 27668 27764 27674
rect 27712 27610 27764 27616
rect 27724 27402 27752 27610
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27528 26920 27580 26926
rect 27528 26862 27580 26868
rect 27448 26586 27476 26862
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 26976 26512 27028 26518
rect 26976 26454 27028 26460
rect 26148 26240 26200 26246
rect 26148 26182 26200 26188
rect 26160 26042 26188 26182
rect 26148 26036 26200 26042
rect 26148 25978 26200 25984
rect 26608 25900 26660 25906
rect 26608 25842 26660 25848
rect 26620 25498 26648 25842
rect 26988 25838 27016 26454
rect 26976 25832 27028 25838
rect 26976 25774 27028 25780
rect 26608 25492 26660 25498
rect 26608 25434 26660 25440
rect 26988 24954 27016 25774
rect 27540 25362 27568 26862
rect 27724 26314 27752 27338
rect 27712 26308 27764 26314
rect 27712 26250 27764 26256
rect 27724 25974 27752 26250
rect 27712 25968 27764 25974
rect 27712 25910 27764 25916
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26988 24682 27016 24890
rect 26976 24676 27028 24682
rect 26976 24618 27028 24624
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25332 22642 25360 24210
rect 26712 24138 26740 24550
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22778 25544 22918
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25320 22636 25372 22642
rect 25320 22578 25372 22584
rect 25332 22234 25360 22578
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25884 22098 25912 23122
rect 26252 23118 26280 23462
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 25872 22092 25924 22098
rect 26252 22094 26280 23054
rect 26528 22778 26556 23734
rect 26988 23730 27016 24618
rect 27172 24342 27200 25094
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27356 23662 27384 23734
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27264 23322 27292 23598
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27724 23118 27752 24006
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27816 22982 27844 24074
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 26516 22772 26568 22778
rect 26516 22714 26568 22720
rect 27816 22642 27844 22918
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 26252 22066 26372 22094
rect 25872 22034 25924 22040
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 25148 21690 25176 21830
rect 26160 21690 26188 21898
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21010 25176 21422
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25516 19174 25544 19858
rect 25976 19446 26004 20810
rect 25964 19440 26016 19446
rect 25964 19382 26016 19388
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25056 18856 25176 18884
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24964 15434 24992 16526
rect 25056 15706 25084 16526
rect 25148 16250 25176 18856
rect 25516 18630 25544 19110
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25608 18766 25636 18906
rect 26252 18902 26280 19246
rect 26240 18896 26292 18902
rect 26240 18838 26292 18844
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25608 18426 25636 18702
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 26160 18290 26188 18566
rect 26344 18358 26372 22066
rect 27540 21486 27568 22510
rect 27712 21956 27764 21962
rect 27712 21898 27764 21904
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27632 21622 27660 21830
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27724 20874 27752 21898
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26804 19378 26832 19790
rect 26976 19780 27028 19786
rect 26976 19722 27028 19728
rect 26988 19378 27016 19722
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 27172 19446 27200 19654
rect 27724 19446 27752 20810
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 26332 18352 26384 18358
rect 26332 18294 26384 18300
rect 26700 18352 26752 18358
rect 26700 18294 26752 18300
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 26344 17746 26372 18022
rect 26332 17740 26384 17746
rect 26332 17682 26384 17688
rect 26712 17610 26740 18294
rect 27724 18290 27752 18702
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27724 17882 27752 18226
rect 27712 17876 27764 17882
rect 27712 17818 27764 17824
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26712 17270 26740 17546
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 27264 17134 27292 17478
rect 27528 17264 27580 17270
rect 27528 17206 27580 17212
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27540 16794 27568 17206
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 27632 16658 27660 16934
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25332 16114 25360 16526
rect 25320 16108 25372 16114
rect 25320 16050 25372 16056
rect 25424 16046 25452 16594
rect 27632 16114 27660 16594
rect 27908 16182 27936 30534
rect 28092 23066 28120 34886
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28184 24206 28212 34546
rect 28552 31958 28580 34614
rect 28724 33992 28776 33998
rect 28724 33934 28776 33940
rect 28632 32768 28684 32774
rect 28632 32710 28684 32716
rect 28644 32570 28672 32710
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28632 32020 28684 32026
rect 28632 31962 28684 31968
rect 28540 31952 28592 31958
rect 28540 31894 28592 31900
rect 28644 31482 28672 31962
rect 28632 31476 28684 31482
rect 28632 31418 28684 31424
rect 28448 30184 28500 30190
rect 28448 30126 28500 30132
rect 28460 29714 28488 30126
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28448 29708 28500 29714
rect 28448 29650 28500 29656
rect 28460 29102 28488 29650
rect 28644 29578 28672 29786
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28448 29096 28500 29102
rect 28448 29038 28500 29044
rect 28460 27334 28488 29038
rect 28644 28966 28672 29514
rect 28632 28960 28684 28966
rect 28632 28902 28684 28908
rect 28644 28558 28672 28902
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 27130 28488 27270
rect 28448 27124 28500 27130
rect 28448 27066 28500 27072
rect 28632 26852 28684 26858
rect 28632 26794 28684 26800
rect 28644 26450 28672 26794
rect 28632 26444 28684 26450
rect 28632 26386 28684 26392
rect 28736 24818 28764 33934
rect 28908 33108 28960 33114
rect 28908 33050 28960 33056
rect 28816 32972 28868 32978
rect 28816 32914 28868 32920
rect 28828 32298 28856 32914
rect 28920 32434 28948 33050
rect 28908 32428 28960 32434
rect 28908 32370 28960 32376
rect 28816 32292 28868 32298
rect 28816 32234 28868 32240
rect 28920 32026 28948 32370
rect 28908 32020 28960 32026
rect 28908 31962 28960 31968
rect 28816 31952 28868 31958
rect 28816 31894 28868 31900
rect 28828 31754 28856 31894
rect 28828 31726 28948 31754
rect 28816 26920 28868 26926
rect 28816 26862 28868 26868
rect 28828 26586 28856 26862
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28264 24064 28316 24070
rect 28264 24006 28316 24012
rect 28276 23118 28304 24006
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28264 23112 28316 23118
rect 28092 23038 28212 23066
rect 28264 23054 28316 23060
rect 28184 22982 28212 23038
rect 28172 22976 28224 22982
rect 28172 22918 28224 22924
rect 28184 22778 28212 22918
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28184 22166 28212 22578
rect 28552 22506 28580 23734
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28828 23186 28856 23462
rect 28816 23180 28868 23186
rect 28816 23122 28868 23128
rect 28920 23066 28948 31726
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 29012 30190 29040 30670
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 29012 29850 29040 30126
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 29012 26586 29040 26930
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 29012 26382 29040 26522
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 29012 25702 29040 26318
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29012 25158 29040 25638
rect 29092 25356 29144 25362
rect 29092 25298 29144 25304
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 29104 24954 29132 25298
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29196 24206 29224 35974
rect 29380 35958 29776 35986
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 29368 34196 29420 34202
rect 29368 34138 29420 34144
rect 29380 33318 29408 34138
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29368 33312 29420 33318
rect 29288 33272 29368 33300
rect 29288 31822 29316 33272
rect 29368 33254 29420 33260
rect 29472 33046 29500 33390
rect 29564 33318 29592 35634
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29460 33040 29512 33046
rect 29460 32982 29512 32988
rect 29564 32842 29592 33254
rect 29644 32972 29696 32978
rect 29644 32914 29696 32920
rect 29552 32836 29604 32842
rect 29552 32778 29604 32784
rect 29656 32570 29684 32914
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29368 32360 29420 32366
rect 29368 32302 29420 32308
rect 29276 31816 29328 31822
rect 29276 31758 29328 31764
rect 29380 31346 29408 32302
rect 29368 31340 29420 31346
rect 29368 31282 29420 31288
rect 29380 29850 29408 31282
rect 29552 30116 29604 30122
rect 29552 30058 29604 30064
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 29564 29646 29592 30058
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29276 27124 29328 27130
rect 29276 27066 29328 27072
rect 29288 26382 29316 27066
rect 29644 26920 29696 26926
rect 29644 26862 29696 26868
rect 29460 26444 29512 26450
rect 29460 26386 29512 26392
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29288 25906 29316 26318
rect 29472 26246 29500 26386
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29460 26240 29512 26246
rect 29460 26182 29512 26188
rect 29276 25900 29328 25906
rect 29276 25842 29328 25848
rect 29288 24954 29316 25842
rect 29472 25770 29500 26182
rect 29460 25764 29512 25770
rect 29460 25706 29512 25712
rect 29276 24948 29328 24954
rect 29276 24890 29328 24896
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29288 24410 29316 24754
rect 29472 24614 29500 25706
rect 29564 25702 29592 26250
rect 29656 26042 29684 26862
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29748 25702 29776 35958
rect 29840 35562 29868 36110
rect 30024 35698 30052 36110
rect 30944 35834 30972 38286
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 31036 36786 31064 36858
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31680 36378 31708 36654
rect 31668 36372 31720 36378
rect 31668 36314 31720 36320
rect 30932 35828 30984 35834
rect 30932 35770 30984 35776
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 29920 35624 29972 35630
rect 29920 35566 29972 35572
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 29828 35556 29880 35562
rect 29828 35498 29880 35504
rect 29932 35086 29960 35566
rect 30104 35556 30156 35562
rect 30104 35498 30156 35504
rect 30116 35086 30144 35498
rect 30300 35290 30328 35566
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 30104 35080 30156 35086
rect 30104 35022 30156 35028
rect 29932 32434 29960 35022
rect 30288 34944 30340 34950
rect 30288 34886 30340 34892
rect 30102 33144 30158 33153
rect 30300 33114 30328 34886
rect 31668 34672 31720 34678
rect 31668 34614 31720 34620
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 30748 33448 30800 33454
rect 30748 33390 30800 33396
rect 30760 33114 30788 33390
rect 30102 33079 30158 33088
rect 30288 33108 30340 33114
rect 30116 33046 30144 33079
rect 30288 33050 30340 33056
rect 30748 33108 30800 33114
rect 30748 33050 30800 33056
rect 30104 33040 30156 33046
rect 30104 32982 30156 32988
rect 31496 32910 31524 34478
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30932 32904 30984 32910
rect 30932 32846 30984 32852
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 30208 32434 30236 32846
rect 30944 32570 30972 32846
rect 31404 32570 31432 32846
rect 31680 32842 31708 34614
rect 31760 33448 31812 33454
rect 31760 33390 31812 33396
rect 31772 32978 31800 33390
rect 31944 33108 31996 33114
rect 31944 33050 31996 33056
rect 31760 32972 31812 32978
rect 31760 32914 31812 32920
rect 31668 32836 31720 32842
rect 31668 32778 31720 32784
rect 30932 32564 30984 32570
rect 30932 32506 30984 32512
rect 31392 32564 31444 32570
rect 31392 32506 31444 32512
rect 31772 32502 31800 32914
rect 31956 32910 31984 33050
rect 31944 32904 31996 32910
rect 31944 32846 31996 32852
rect 31760 32496 31812 32502
rect 31760 32438 31812 32444
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 30196 32428 30248 32434
rect 30196 32370 30248 32376
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29840 31482 29868 31826
rect 29828 31476 29880 31482
rect 29828 31418 29880 31424
rect 29932 31414 29960 32370
rect 30852 32026 30880 32370
rect 30840 32020 30892 32026
rect 30840 31962 30892 31968
rect 29920 31408 29972 31414
rect 29920 31350 29972 31356
rect 29932 30258 29960 31350
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 30116 30938 30144 31214
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30196 30796 30248 30802
rect 30196 30738 30248 30744
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29932 30138 29960 30194
rect 29932 30110 30144 30138
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 29932 29850 29960 29990
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 30024 29714 30052 29990
rect 30116 29782 30144 30110
rect 30208 29850 30236 30738
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 30300 29850 30328 30126
rect 30196 29844 30248 29850
rect 30196 29786 30248 29792
rect 30288 29844 30340 29850
rect 30288 29786 30340 29792
rect 30104 29776 30156 29782
rect 30104 29718 30156 29724
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 30024 29306 30052 29650
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30024 26586 30052 29242
rect 30116 29170 30144 29718
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30484 29238 30512 29582
rect 30472 29232 30524 29238
rect 30472 29174 30524 29180
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30116 27130 30144 29106
rect 31852 28484 31904 28490
rect 31852 28426 31904 28432
rect 31864 27674 31892 28426
rect 31852 27668 31904 27674
rect 31852 27610 31904 27616
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30104 27124 30156 27130
rect 30104 27066 30156 27072
rect 30668 26994 30696 27270
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 31864 26314 31892 27610
rect 30840 26308 30892 26314
rect 30840 26250 30892 26256
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 30852 26042 30880 26250
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29736 25696 29788 25702
rect 29736 25638 29788 25644
rect 29564 25498 29592 25638
rect 31496 25498 31524 25774
rect 31588 25498 31616 25842
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31576 25492 31628 25498
rect 31576 25434 31628 25440
rect 31944 25492 31996 25498
rect 31944 25434 31996 25440
rect 31956 25294 31984 25434
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 29828 25220 29880 25226
rect 29828 25162 29880 25168
rect 29840 24818 29868 25162
rect 31852 25152 31904 25158
rect 31852 25094 31904 25100
rect 29920 24948 29972 24954
rect 29920 24890 29972 24896
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29460 24608 29512 24614
rect 29460 24550 29512 24556
rect 29276 24404 29328 24410
rect 29276 24346 29328 24352
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 28828 23050 28948 23066
rect 29012 23050 29040 23258
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 28816 23044 28948 23050
rect 28868 23038 28948 23044
rect 29000 23044 29052 23050
rect 28816 22986 28868 22992
rect 29000 22986 29052 22992
rect 29104 22982 29132 23054
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28540 22500 28592 22506
rect 28540 22442 28592 22448
rect 28172 22160 28224 22166
rect 28172 22102 28224 22108
rect 28080 21684 28132 21690
rect 28080 21626 28132 21632
rect 28092 21350 28120 21626
rect 28184 21486 28212 22102
rect 28552 21962 28580 22442
rect 28920 21962 28948 22578
rect 29104 22234 29132 22918
rect 29196 22642 29224 24142
rect 29288 22642 29316 24346
rect 29472 24138 29500 24550
rect 29748 24410 29776 24686
rect 29736 24404 29788 24410
rect 29736 24346 29788 24352
rect 29932 24206 29960 24890
rect 31864 24886 31892 25094
rect 31956 24954 31984 25230
rect 31944 24948 31996 24954
rect 31944 24890 31996 24896
rect 31852 24880 31904 24886
rect 31852 24822 31904 24828
rect 31944 24336 31996 24342
rect 31944 24278 31996 24284
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 29460 24132 29512 24138
rect 29460 24074 29512 24080
rect 29368 23656 29420 23662
rect 29368 23598 29420 23604
rect 29380 23050 29408 23598
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 29276 22636 29328 22642
rect 29276 22578 29328 22584
rect 29092 22228 29144 22234
rect 29092 22170 29144 22176
rect 29288 22030 29316 22578
rect 29380 22166 29408 22714
rect 29368 22160 29420 22166
rect 29368 22102 29420 22108
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28908 21956 28960 21962
rect 28908 21898 28960 21904
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28920 21418 28948 21898
rect 29288 21622 29316 21966
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 28092 20806 28120 21286
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 29012 19922 29040 21286
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28736 19514 28764 19790
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28632 18828 28684 18834
rect 28632 18770 28684 18776
rect 28644 18426 28672 18770
rect 28632 18420 28684 18426
rect 28632 18362 28684 18368
rect 28736 18290 28764 19246
rect 28920 19242 28948 19722
rect 29012 19718 29040 19858
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 29012 19378 29040 19654
rect 29196 19378 29224 19994
rect 29288 19446 29316 21558
rect 29472 20058 29500 24074
rect 31956 23594 31984 24278
rect 31944 23588 31996 23594
rect 31944 23530 31996 23536
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29748 22778 29776 23258
rect 30932 23180 30984 23186
rect 30932 23122 30984 23128
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30300 22778 30328 23054
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30392 22778 30420 22986
rect 29736 22772 29788 22778
rect 29736 22714 29788 22720
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30380 22772 30432 22778
rect 30380 22714 30432 22720
rect 30852 22506 30880 22986
rect 30944 22778 30972 23122
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 30840 22500 30892 22506
rect 30840 22442 30892 22448
rect 29644 22432 29696 22438
rect 29644 22374 29696 22380
rect 29656 22098 29684 22374
rect 31956 22234 31984 23530
rect 31944 22228 31996 22234
rect 31944 22170 31996 22176
rect 29644 22092 29696 22098
rect 32048 22094 32076 45766
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 33048 43852 33100 43858
rect 33048 43794 33100 43800
rect 32220 43376 32272 43382
rect 32220 43318 32272 43324
rect 32232 43110 32260 43318
rect 32220 43104 32272 43110
rect 32220 43046 32272 43052
rect 32128 41132 32180 41138
rect 32128 41074 32180 41080
rect 32140 41041 32168 41074
rect 32126 41032 32182 41041
rect 32126 40967 32182 40976
rect 32232 39506 32260 43046
rect 33060 42906 33088 43794
rect 33968 43648 34020 43654
rect 33968 43590 34020 43596
rect 33876 43308 33928 43314
rect 33876 43250 33928 43256
rect 33048 42900 33100 42906
rect 33048 42842 33100 42848
rect 32496 42832 32548 42838
rect 32496 42774 32548 42780
rect 32508 42566 32536 42774
rect 32680 42696 32732 42702
rect 32680 42638 32732 42644
rect 33232 42696 33284 42702
rect 33232 42638 33284 42644
rect 32588 42628 32640 42634
rect 32588 42570 32640 42576
rect 32496 42560 32548 42566
rect 32496 42502 32548 42508
rect 32508 41614 32536 42502
rect 32600 42362 32628 42570
rect 32588 42356 32640 42362
rect 32588 42298 32640 42304
rect 32600 41721 32628 42298
rect 32586 41712 32642 41721
rect 32586 41647 32642 41656
rect 32496 41608 32548 41614
rect 32496 41550 32548 41556
rect 32496 41200 32548 41206
rect 32494 41168 32496 41177
rect 32548 41168 32550 41177
rect 32404 41132 32456 41138
rect 32494 41103 32550 41112
rect 32404 41074 32456 41080
rect 32416 40594 32444 41074
rect 32404 40588 32456 40594
rect 32404 40530 32456 40536
rect 32220 39500 32272 39506
rect 32220 39442 32272 39448
rect 32416 39098 32444 40530
rect 32404 39092 32456 39098
rect 32404 39034 32456 39040
rect 32600 38654 32628 41647
rect 32692 41614 32720 42638
rect 33140 42560 33192 42566
rect 33140 42502 33192 42508
rect 32772 42016 32824 42022
rect 32772 41958 32824 41964
rect 32784 41682 32812 41958
rect 33152 41818 33180 42502
rect 33244 42294 33272 42638
rect 33324 42560 33376 42566
rect 33324 42502 33376 42508
rect 33232 42288 33284 42294
rect 33232 42230 33284 42236
rect 33336 42226 33364 42502
rect 33784 42356 33836 42362
rect 33784 42298 33836 42304
rect 33692 42288 33744 42294
rect 33692 42230 33744 42236
rect 33324 42220 33376 42226
rect 33324 42162 33376 42168
rect 33508 42016 33560 42022
rect 33508 41958 33560 41964
rect 33140 41812 33192 41818
rect 33140 41754 33192 41760
rect 33048 41744 33100 41750
rect 33048 41686 33100 41692
rect 32772 41676 32824 41682
rect 32772 41618 32824 41624
rect 32680 41608 32732 41614
rect 32680 41550 32732 41556
rect 33060 41206 33088 41686
rect 33520 41614 33548 41958
rect 33508 41608 33560 41614
rect 33508 41550 33560 41556
rect 33598 41576 33654 41585
rect 33416 41540 33468 41546
rect 33598 41511 33600 41520
rect 33416 41482 33468 41488
rect 33652 41511 33654 41520
rect 33600 41482 33652 41488
rect 33428 41414 33456 41482
rect 33428 41386 33640 41414
rect 33048 41200 33100 41206
rect 33048 41142 33100 41148
rect 33612 41138 33640 41386
rect 33704 41274 33732 42230
rect 33796 41818 33824 42298
rect 33784 41812 33836 41818
rect 33784 41754 33836 41760
rect 33784 41608 33836 41614
rect 33784 41550 33836 41556
rect 33692 41268 33744 41274
rect 33692 41210 33744 41216
rect 33796 41138 33824 41550
rect 33600 41132 33652 41138
rect 33600 41074 33652 41080
rect 33784 41132 33836 41138
rect 33784 41074 33836 41080
rect 32968 39086 33456 39114
rect 32968 38978 32996 39086
rect 32876 38962 32996 38978
rect 33060 38962 33180 38978
rect 33428 38962 33456 39086
rect 33612 39030 33640 41074
rect 33888 39030 33916 43250
rect 33980 43246 34008 43590
rect 35532 43308 35584 43314
rect 35532 43250 35584 43256
rect 33968 43240 34020 43246
rect 33968 43182 34020 43188
rect 34244 43240 34296 43246
rect 34244 43182 34296 43188
rect 34256 42362 34284 43182
rect 35544 43110 35572 43250
rect 35532 43104 35584 43110
rect 35532 43046 35584 43052
rect 35716 43104 35768 43110
rect 35716 43046 35768 43052
rect 36912 43104 36964 43110
rect 36912 43046 36964 43052
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35728 42770 35756 43046
rect 35256 42764 35308 42770
rect 35256 42706 35308 42712
rect 35716 42764 35768 42770
rect 35716 42706 35768 42712
rect 34888 42560 34940 42566
rect 34888 42502 34940 42508
rect 34900 42362 34928 42502
rect 34244 42356 34296 42362
rect 34244 42298 34296 42304
rect 34888 42356 34940 42362
rect 34888 42298 34940 42304
rect 34152 42288 34204 42294
rect 34152 42230 34204 42236
rect 34704 42288 34756 42294
rect 34704 42230 34756 42236
rect 34796 42288 34848 42294
rect 34796 42230 34848 42236
rect 34164 41614 34192 42230
rect 34716 42090 34744 42230
rect 34704 42084 34756 42090
rect 34704 42026 34756 42032
rect 34716 41750 34744 42026
rect 34704 41744 34756 41750
rect 34704 41686 34756 41692
rect 34808 41682 34836 42230
rect 35268 42226 35296 42706
rect 35256 42220 35308 42226
rect 35256 42162 35308 42168
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34796 41676 34848 41682
rect 34796 41618 34848 41624
rect 34060 41608 34112 41614
rect 34060 41550 34112 41556
rect 34152 41608 34204 41614
rect 34704 41608 34756 41614
rect 34152 41550 34204 41556
rect 34334 41576 34390 41585
rect 34072 41460 34100 41550
rect 34704 41550 34756 41556
rect 34334 41511 34336 41520
rect 34388 41511 34390 41520
rect 34336 41482 34388 41488
rect 34072 41432 34284 41460
rect 34256 41274 34284 41432
rect 34244 41268 34296 41274
rect 34244 41210 34296 41216
rect 34348 41138 34376 41482
rect 34716 41206 34744 41550
rect 34808 41274 34836 41618
rect 35532 41540 35584 41546
rect 35532 41482 35584 41488
rect 35070 41304 35126 41313
rect 34796 41268 34848 41274
rect 35544 41274 35572 41482
rect 35070 41239 35072 41248
rect 34796 41210 34848 41216
rect 35124 41239 35126 41248
rect 35532 41268 35584 41274
rect 35072 41210 35124 41216
rect 35532 41210 35584 41216
rect 34704 41200 34756 41206
rect 34704 41142 34756 41148
rect 34336 41132 34388 41138
rect 34336 41074 34388 41080
rect 34520 41132 34572 41138
rect 34520 41074 34572 41080
rect 34532 41018 34560 41074
rect 34440 40990 34560 41018
rect 34440 40934 34468 40990
rect 34428 40928 34480 40934
rect 34428 40870 34480 40876
rect 35808 40928 35860 40934
rect 35808 40870 35860 40876
rect 35900 40928 35952 40934
rect 35900 40870 35952 40876
rect 34060 40112 34112 40118
rect 34060 40054 34112 40060
rect 33600 39024 33652 39030
rect 33600 38966 33652 38972
rect 33876 39024 33928 39030
rect 33876 38966 33928 38972
rect 32864 38956 32996 38962
rect 32916 38950 32996 38956
rect 33048 38956 33180 38962
rect 32864 38898 32916 38904
rect 33100 38950 33180 38956
rect 33048 38898 33100 38904
rect 33152 38826 33180 38950
rect 33416 38956 33468 38962
rect 33416 38898 33468 38904
rect 33140 38820 33192 38826
rect 33140 38762 33192 38768
rect 33324 38820 33376 38826
rect 33324 38762 33376 38768
rect 32600 38626 32720 38654
rect 32404 38344 32456 38350
rect 32404 38286 32456 38292
rect 32416 37874 32444 38286
rect 32404 37868 32456 37874
rect 32404 37810 32456 37816
rect 32416 37262 32444 37810
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 32416 36718 32444 37198
rect 32404 36712 32456 36718
rect 32404 36654 32456 36660
rect 32416 35834 32444 36654
rect 32692 36174 32720 38626
rect 33152 38554 33180 38762
rect 33140 38548 33192 38554
rect 33140 38490 33192 38496
rect 33336 38418 33364 38762
rect 33324 38412 33376 38418
rect 33324 38354 33376 38360
rect 33428 38350 33456 38898
rect 33508 38752 33560 38758
rect 33508 38694 33560 38700
rect 33520 38350 33548 38694
rect 33416 38344 33468 38350
rect 33416 38286 33468 38292
rect 33508 38344 33560 38350
rect 33508 38286 33560 38292
rect 33692 38344 33744 38350
rect 33692 38286 33744 38292
rect 32772 38208 32824 38214
rect 32772 38150 32824 38156
rect 33232 38208 33284 38214
rect 33232 38150 33284 38156
rect 33508 38208 33560 38214
rect 33508 38150 33560 38156
rect 32784 37874 32812 38150
rect 32772 37868 32824 37874
rect 32772 37810 32824 37816
rect 32784 37262 32812 37810
rect 33244 37670 33272 38150
rect 33232 37664 33284 37670
rect 33232 37606 33284 37612
rect 33244 37466 33272 37606
rect 33232 37460 33284 37466
rect 33232 37402 33284 37408
rect 32772 37256 32824 37262
rect 32772 37198 32824 37204
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32784 36786 32812 37198
rect 32772 36780 32824 36786
rect 32772 36722 32824 36728
rect 32864 36644 32916 36650
rect 32864 36586 32916 36592
rect 32876 36378 32904 36586
rect 33048 36576 33100 36582
rect 33048 36518 33100 36524
rect 32864 36372 32916 36378
rect 32864 36314 32916 36320
rect 33060 36174 33088 36518
rect 32680 36168 32732 36174
rect 32680 36110 32732 36116
rect 32772 36168 32824 36174
rect 32772 36110 32824 36116
rect 33048 36168 33100 36174
rect 33048 36110 33100 36116
rect 32404 35828 32456 35834
rect 32404 35770 32456 35776
rect 32588 34672 32640 34678
rect 32588 34614 32640 34620
rect 32600 34406 32628 34614
rect 32588 34400 32640 34406
rect 32588 34342 32640 34348
rect 32128 33312 32180 33318
rect 32128 33254 32180 33260
rect 32140 32978 32168 33254
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 32496 32972 32548 32978
rect 32496 32914 32548 32920
rect 32220 32768 32272 32774
rect 32220 32710 32272 32716
rect 32232 32502 32260 32710
rect 32220 32496 32272 32502
rect 32220 32438 32272 32444
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32416 32026 32444 32370
rect 32404 32020 32456 32026
rect 32404 31962 32456 31968
rect 32508 31958 32536 32914
rect 32600 32434 32628 34342
rect 32692 33114 32720 36110
rect 32784 35834 32812 36110
rect 32864 36100 32916 36106
rect 32864 36042 32916 36048
rect 32876 35834 32904 36042
rect 32772 35828 32824 35834
rect 32772 35770 32824 35776
rect 32864 35828 32916 35834
rect 32864 35770 32916 35776
rect 33152 35086 33180 37198
rect 33416 36644 33468 36650
rect 33416 36586 33468 36592
rect 33428 35698 33456 36586
rect 33416 35692 33468 35698
rect 33416 35634 33468 35640
rect 33520 35562 33548 38150
rect 33704 38010 33732 38286
rect 33692 38004 33744 38010
rect 33692 37946 33744 37952
rect 33784 36780 33836 36786
rect 33784 36722 33836 36728
rect 33600 35624 33652 35630
rect 33600 35566 33652 35572
rect 33508 35556 33560 35562
rect 33508 35498 33560 35504
rect 33520 35086 33548 35498
rect 33612 35290 33640 35566
rect 33600 35284 33652 35290
rect 33600 35226 33652 35232
rect 33140 35080 33192 35086
rect 33140 35022 33192 35028
rect 33324 35080 33376 35086
rect 33324 35022 33376 35028
rect 33508 35080 33560 35086
rect 33508 35022 33560 35028
rect 33152 34746 33180 35022
rect 33336 34746 33364 35022
rect 33140 34740 33192 34746
rect 33140 34682 33192 34688
rect 33324 34740 33376 34746
rect 33324 34682 33376 34688
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 33048 34196 33100 34202
rect 33100 34156 33180 34184
rect 33048 34138 33100 34144
rect 33048 34060 33100 34066
rect 32968 34020 33048 34048
rect 32864 33924 32916 33930
rect 32864 33866 32916 33872
rect 32680 33108 32732 33114
rect 32680 33050 32732 33056
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32496 31952 32548 31958
rect 32496 31894 32548 31900
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32324 31482 32352 31758
rect 32508 31482 32536 31758
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32496 31476 32548 31482
rect 32496 31418 32548 31424
rect 32600 30326 32628 32370
rect 32692 32230 32720 33050
rect 32680 32224 32732 32230
rect 32680 32166 32732 32172
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32220 30048 32272 30054
rect 32220 29990 32272 29996
rect 32232 29782 32260 29990
rect 32312 29844 32364 29850
rect 32312 29786 32364 29792
rect 32220 29776 32272 29782
rect 32220 29718 32272 29724
rect 32220 29504 32272 29510
rect 32220 29446 32272 29452
rect 32232 29306 32260 29446
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32324 29034 32352 29786
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32312 29028 32364 29034
rect 32312 28970 32364 28976
rect 32692 28558 32720 29106
rect 32680 28552 32732 28558
rect 32680 28494 32732 28500
rect 32692 28422 32720 28494
rect 32680 28416 32732 28422
rect 32680 28358 32732 28364
rect 32220 26444 32272 26450
rect 32220 26386 32272 26392
rect 32128 26240 32180 26246
rect 32128 26182 32180 26188
rect 32140 25974 32168 26182
rect 32128 25968 32180 25974
rect 32128 25910 32180 25916
rect 32232 25906 32260 26386
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 32128 25764 32180 25770
rect 32128 25706 32180 25712
rect 32140 25362 32168 25706
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 32232 25294 32260 25842
rect 32404 25696 32456 25702
rect 32404 25638 32456 25644
rect 32220 25288 32272 25294
rect 32220 25230 32272 25236
rect 32416 25158 32444 25638
rect 32404 25152 32456 25158
rect 32404 25094 32456 25100
rect 32220 24880 32272 24886
rect 32508 24834 32536 25842
rect 32692 25498 32720 25842
rect 32680 25492 32732 25498
rect 32680 25434 32732 25440
rect 32272 24828 32536 24834
rect 32220 24822 32536 24828
rect 32128 24812 32180 24818
rect 32232 24806 32536 24822
rect 32128 24754 32180 24760
rect 32140 24410 32168 24754
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32140 23322 32168 23666
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 29644 22034 29696 22040
rect 31864 22066 32076 22094
rect 29656 21554 29684 22034
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29748 21690 29776 21830
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 29656 19514 29684 19858
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29748 19514 29776 19654
rect 31036 19514 31064 19790
rect 31312 19786 31340 20402
rect 31404 19990 31432 20402
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 31392 19984 31444 19990
rect 31392 19926 31444 19932
rect 31666 19952 31722 19961
rect 31404 19854 31432 19926
rect 31666 19887 31668 19896
rect 31720 19887 31722 19896
rect 31668 19858 31720 19864
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31300 19780 31352 19786
rect 31300 19722 31352 19728
rect 31404 19514 31432 19790
rect 31772 19718 31800 20266
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 29276 19440 29328 19446
rect 29276 19382 29328 19388
rect 31864 19394 31892 22066
rect 32036 21004 32088 21010
rect 32036 20946 32088 20952
rect 32048 20602 32076 20946
rect 32036 20596 32088 20602
rect 32036 20538 32088 20544
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 31956 20058 31984 20402
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 31956 19854 31984 19994
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31956 19514 31984 19790
rect 31944 19508 31996 19514
rect 31944 19450 31996 19456
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 28908 19236 28960 19242
rect 28908 19178 28960 19184
rect 28816 18896 28868 18902
rect 28920 18884 28948 19178
rect 28868 18856 28948 18884
rect 28816 18838 28868 18844
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29012 18222 29040 19314
rect 29288 19310 29316 19382
rect 31484 19372 31536 19378
rect 31864 19366 31984 19394
rect 31484 19314 31536 19320
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30760 18766 30788 19110
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 31496 18222 31524 19314
rect 31760 19168 31812 19174
rect 31760 19110 31812 19116
rect 31772 18834 31800 19110
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31852 18692 31904 18698
rect 31852 18634 31904 18640
rect 31864 18358 31892 18634
rect 31852 18352 31904 18358
rect 31852 18294 31904 18300
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 31484 18216 31536 18222
rect 31484 18158 31536 18164
rect 30944 17882 30972 18158
rect 30932 17876 30984 17882
rect 30932 17818 30984 17824
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 28092 16794 28120 17478
rect 28920 17338 28948 17614
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 30932 17264 30984 17270
rect 30932 17206 30984 17212
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 28920 16590 28948 17070
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16250 28212 16458
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 27896 16176 27948 16182
rect 27896 16118 27948 16124
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 14618 25176 15302
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 25044 14068 25096 14074
rect 25424 14056 25452 15982
rect 25608 15026 25636 15982
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25884 14958 25912 15506
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25884 14482 25912 14894
rect 25872 14476 25924 14482
rect 25872 14418 25924 14424
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25096 14028 25452 14056
rect 25044 14010 25096 14016
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24964 13530 24992 13738
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24872 11354 24900 13330
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24964 12918 24992 13262
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 25056 12782 25084 14010
rect 25608 13938 25636 14214
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25608 13462 25636 13874
rect 25596 13456 25648 13462
rect 25596 13398 25648 13404
rect 25884 13326 25912 14418
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25792 12986 25820 13194
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25228 12912 25280 12918
rect 25228 12854 25280 12860
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25240 11898 25268 12854
rect 25884 12782 25912 13262
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25148 11354 25176 11698
rect 25424 11694 25452 12718
rect 25976 11762 26004 14962
rect 26068 13462 26096 15982
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26344 14958 26372 15302
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26160 14618 26188 14758
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 25148 10130 25176 11290
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25332 10810 25360 11086
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25424 10538 25452 11630
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25424 10198 25452 10474
rect 25412 10192 25464 10198
rect 25412 10134 25464 10140
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25056 8634 25084 8910
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25240 8634 25268 8774
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25332 8430 25360 8978
rect 25608 8634 25636 9862
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25700 9178 25728 9318
rect 25792 9178 25820 10066
rect 25976 9450 26004 11698
rect 26160 11694 26188 14010
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26252 12986 26280 13126
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26068 11150 26096 11630
rect 26160 11286 26188 11630
rect 26148 11280 26200 11286
rect 26148 11222 26200 11228
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26068 10810 26096 11086
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 26160 10130 26188 11222
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 25964 9444 26016 9450
rect 25964 9386 26016 9392
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 26160 9042 26188 10066
rect 26252 9518 26280 10542
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25332 7546 25360 8366
rect 25608 8090 25636 8570
rect 25792 8430 25820 8842
rect 26344 8634 26372 14894
rect 26528 14278 26556 15642
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26804 14482 26832 15506
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26896 15026 26924 15302
rect 26884 15020 26936 15026
rect 26884 14962 26936 14968
rect 26792 14476 26844 14482
rect 26620 14436 26792 14464
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26528 13190 26556 14214
rect 26620 14074 26648 14436
rect 26792 14418 26844 14424
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 14074 26740 14214
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26620 13530 26648 14010
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 26804 13530 26832 13738
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26608 13320 26660 13326
rect 26792 13320 26844 13326
rect 26660 13280 26792 13308
rect 26608 13262 26660 13268
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26516 10532 26568 10538
rect 26516 10474 26568 10480
rect 26528 10130 26556 10474
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26712 9674 26740 13280
rect 26792 13262 26844 13268
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 26804 10266 26832 10610
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 26804 9722 26832 10202
rect 26436 9646 26740 9674
rect 26792 9716 26844 9722
rect 26792 9658 26844 9664
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23584 6322 23612 6802
rect 24412 6798 24440 7278
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24320 6390 24348 6734
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23768 5914 23796 6054
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 23112 5092 23164 5098
rect 23112 5034 23164 5040
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 23124 4622 23152 5034
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4826 23244 4966
rect 23584 4826 23612 5510
rect 23860 5166 23888 5850
rect 23952 5710 23980 6054
rect 24320 5846 24348 6326
rect 24412 6322 24440 6734
rect 24872 6730 24900 7346
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 25056 6662 25084 6938
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24780 6322 24808 6598
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 24136 5098 24164 5646
rect 24320 5574 24348 5782
rect 24412 5710 24440 6258
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24320 5234 24348 5510
rect 24872 5234 24900 6122
rect 25056 6118 25084 6598
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25240 5914 25268 6054
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23768 4690 23796 4966
rect 23860 4826 23888 4966
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19524 4004 19576 4010
rect 19444 3964 19524 3992
rect 19524 3946 19576 3952
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3602 18736 3878
rect 19628 3738 19656 4082
rect 20548 4078 20576 4558
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 23768 3534 23796 4626
rect 24504 3738 24532 4966
rect 24872 4622 24900 5170
rect 25228 5092 25280 5098
rect 25332 5080 25360 6938
rect 25792 6866 25820 8366
rect 26436 8362 26464 9646
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26712 8090 26740 8434
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26896 7546 26924 14962
rect 26988 14618 27016 15438
rect 27068 14952 27120 14958
rect 27068 14894 27120 14900
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 27080 14278 27108 14894
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26988 11676 27016 13262
rect 27080 11898 27108 14214
rect 28920 14074 28948 16526
rect 29196 16182 29224 16526
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29380 16114 29408 16390
rect 30944 16182 30972 17206
rect 31116 16992 31168 16998
rect 31116 16934 31168 16940
rect 30932 16176 30984 16182
rect 30932 16118 30984 16124
rect 31128 16114 31156 16934
rect 31956 16726 31984 19366
rect 32140 19310 32168 22510
rect 32324 21146 32352 24142
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 32416 23322 32444 23666
rect 32404 23316 32456 23322
rect 32404 23258 32456 23264
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32416 20466 32444 20878
rect 32508 20602 32536 24806
rect 32680 24676 32732 24682
rect 32680 24618 32732 24624
rect 32692 24410 32720 24618
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 32876 24342 32904 33866
rect 32968 33046 32996 34020
rect 33048 34002 33100 34008
rect 33152 33998 33180 34156
rect 33244 34066 33272 34546
rect 33324 34400 33376 34406
rect 33324 34342 33376 34348
rect 33336 34202 33364 34342
rect 33324 34196 33376 34202
rect 33324 34138 33376 34144
rect 33232 34060 33284 34066
rect 33232 34002 33284 34008
rect 33140 33992 33192 33998
rect 33140 33934 33192 33940
rect 33140 33856 33192 33862
rect 33140 33798 33192 33804
rect 32956 33040 33008 33046
rect 32956 32982 33008 32988
rect 33048 33040 33100 33046
rect 33048 32982 33100 32988
rect 33060 32434 33088 32982
rect 33048 32428 33100 32434
rect 33048 32370 33100 32376
rect 33152 32366 33180 33798
rect 33244 32910 33272 34002
rect 33416 33992 33468 33998
rect 33336 33940 33416 33946
rect 33336 33934 33468 33940
rect 33336 33918 33456 33934
rect 33336 32978 33364 33918
rect 33416 33856 33468 33862
rect 33416 33798 33468 33804
rect 33324 32972 33376 32978
rect 33324 32914 33376 32920
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 33140 32360 33192 32366
rect 33140 32302 33192 32308
rect 33244 32026 33272 32846
rect 33324 32768 33376 32774
rect 33324 32710 33376 32716
rect 33336 32314 33364 32710
rect 33428 32434 33456 33798
rect 33520 32910 33548 35022
rect 33598 34640 33654 34649
rect 33598 34575 33600 34584
rect 33652 34575 33654 34584
rect 33600 34546 33652 34552
rect 33692 34196 33744 34202
rect 33692 34138 33744 34144
rect 33600 33992 33652 33998
rect 33600 33934 33652 33940
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33612 32502 33640 33934
rect 33704 33046 33732 34138
rect 33796 34082 33824 36722
rect 33888 34202 33916 38966
rect 34072 38962 34100 40054
rect 34336 40044 34388 40050
rect 34336 39986 34388 39992
rect 34348 39302 34376 39986
rect 34440 39982 34468 40870
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35256 40520 35308 40526
rect 35256 40462 35308 40468
rect 35268 40186 35296 40462
rect 35820 40458 35848 40870
rect 35532 40452 35584 40458
rect 35532 40394 35584 40400
rect 35808 40452 35860 40458
rect 35808 40394 35860 40400
rect 35544 40186 35572 40394
rect 35256 40180 35308 40186
rect 35256 40122 35308 40128
rect 35532 40180 35584 40186
rect 35532 40122 35584 40128
rect 34428 39976 34480 39982
rect 34428 39918 34480 39924
rect 35440 39976 35492 39982
rect 35440 39918 35492 39924
rect 34152 39296 34204 39302
rect 34152 39238 34204 39244
rect 34336 39296 34388 39302
rect 34336 39238 34388 39244
rect 34060 38956 34112 38962
rect 34060 38898 34112 38904
rect 34072 38842 34100 38898
rect 34164 38894 34192 39238
rect 34348 38962 34376 39238
rect 34336 38956 34388 38962
rect 34336 38898 34388 38904
rect 33980 38814 34100 38842
rect 34152 38888 34204 38894
rect 34152 38830 34204 38836
rect 33980 38554 34008 38814
rect 34060 38752 34112 38758
rect 34060 38694 34112 38700
rect 33968 38548 34020 38554
rect 33968 38490 34020 38496
rect 34072 38350 34100 38694
rect 34440 38350 34468 39918
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35452 39098 35480 39918
rect 35624 39432 35676 39438
rect 35624 39374 35676 39380
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 35636 38962 35664 39374
rect 35820 39370 35848 40394
rect 35912 40390 35940 40870
rect 35992 40520 36044 40526
rect 35992 40462 36044 40468
rect 35900 40384 35952 40390
rect 35900 40326 35952 40332
rect 35912 40050 35940 40326
rect 35900 40044 35952 40050
rect 35900 39986 35952 39992
rect 36004 39438 36032 40462
rect 36924 40458 36952 43046
rect 38016 40520 38068 40526
rect 38016 40462 38068 40468
rect 36912 40452 36964 40458
rect 36912 40394 36964 40400
rect 37188 40384 37240 40390
rect 37188 40326 37240 40332
rect 35992 39432 36044 39438
rect 35992 39374 36044 39380
rect 35808 39364 35860 39370
rect 35808 39306 35860 39312
rect 35900 39364 35952 39370
rect 35900 39306 35952 39312
rect 35256 38956 35308 38962
rect 35256 38898 35308 38904
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 35716 38956 35768 38962
rect 35716 38898 35768 38904
rect 34704 38888 34756 38894
rect 34704 38830 34756 38836
rect 34716 38554 34744 38830
rect 34796 38752 34848 38758
rect 34796 38694 34848 38700
rect 35268 38706 35296 38898
rect 35532 38888 35584 38894
rect 35532 38830 35584 38836
rect 34704 38548 34756 38554
rect 34704 38490 34756 38496
rect 34808 38350 34836 38694
rect 35268 38678 35388 38706
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35360 38554 35388 38678
rect 35348 38548 35400 38554
rect 35348 38490 35400 38496
rect 34060 38344 34112 38350
rect 34060 38286 34112 38292
rect 34428 38344 34480 38350
rect 34428 38286 34480 38292
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 35348 38344 35400 38350
rect 35348 38286 35400 38292
rect 33968 36780 34020 36786
rect 33968 36722 34020 36728
rect 33980 35834 34008 36722
rect 34072 35834 34100 38286
rect 34808 38214 34836 38286
rect 35360 38214 35388 38286
rect 35544 38282 35572 38830
rect 35728 38554 35756 38898
rect 35716 38548 35768 38554
rect 35716 38490 35768 38496
rect 35532 38276 35584 38282
rect 35532 38218 35584 38224
rect 34796 38208 34848 38214
rect 34796 38150 34848 38156
rect 35348 38208 35400 38214
rect 35348 38150 35400 38156
rect 34612 36848 34664 36854
rect 34612 36790 34664 36796
rect 34336 36780 34388 36786
rect 34336 36722 34388 36728
rect 34348 36281 34376 36722
rect 34520 36576 34572 36582
rect 34520 36518 34572 36524
rect 34532 36378 34560 36518
rect 34520 36372 34572 36378
rect 34520 36314 34572 36320
rect 34334 36272 34390 36281
rect 34334 36207 34390 36216
rect 33968 35828 34020 35834
rect 33968 35770 34020 35776
rect 34060 35828 34112 35834
rect 34060 35770 34112 35776
rect 34152 35692 34204 35698
rect 34152 35634 34204 35640
rect 34164 35290 34192 35634
rect 34152 35284 34204 35290
rect 34152 35226 34204 35232
rect 34060 34604 34112 34610
rect 34060 34546 34112 34552
rect 34072 34202 34100 34546
rect 33876 34196 33928 34202
rect 33876 34138 33928 34144
rect 34060 34196 34112 34202
rect 34060 34138 34112 34144
rect 33796 34054 33916 34082
rect 33692 33040 33744 33046
rect 33692 32982 33744 32988
rect 33784 32904 33836 32910
rect 33784 32846 33836 32852
rect 33796 32570 33824 32846
rect 33888 32842 33916 34054
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 33980 33658 34008 33934
rect 33968 33652 34020 33658
rect 33968 33594 34020 33600
rect 34060 33380 34112 33386
rect 34060 33322 34112 33328
rect 34072 32842 34100 33322
rect 34348 32910 34376 36207
rect 34624 35834 34652 36790
rect 34704 36032 34756 36038
rect 34808 36020 34836 38150
rect 35532 37800 35584 37806
rect 35532 37742 35584 37748
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35544 37330 35572 37742
rect 35532 37324 35584 37330
rect 35532 37266 35584 37272
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35544 36378 35572 37266
rect 35716 36712 35768 36718
rect 35820 36700 35848 39306
rect 35912 39098 35940 39306
rect 35900 39092 35952 39098
rect 35900 39034 35952 39040
rect 36004 38554 36032 39374
rect 37200 39370 37228 40326
rect 38028 39982 38056 40462
rect 40500 40112 40552 40118
rect 40500 40054 40552 40060
rect 38016 39976 38068 39982
rect 38016 39918 38068 39924
rect 39120 39976 39172 39982
rect 39120 39918 39172 39924
rect 38028 39438 38056 39918
rect 38016 39432 38068 39438
rect 38016 39374 38068 39380
rect 38292 39432 38344 39438
rect 38292 39374 38344 39380
rect 37188 39364 37240 39370
rect 37188 39306 37240 39312
rect 36268 39296 36320 39302
rect 36268 39238 36320 39244
rect 36280 38962 36308 39238
rect 36268 38956 36320 38962
rect 36268 38898 36320 38904
rect 37004 38956 37056 38962
rect 37004 38898 37056 38904
rect 37016 38554 37044 38898
rect 35992 38548 36044 38554
rect 35992 38490 36044 38496
rect 37004 38548 37056 38554
rect 37004 38490 37056 38496
rect 35900 37324 35952 37330
rect 35900 37266 35952 37272
rect 35912 36922 35940 37266
rect 35900 36916 35952 36922
rect 35900 36858 35952 36864
rect 36004 36786 36032 38490
rect 37016 38350 37044 38490
rect 36544 38344 36596 38350
rect 36544 38286 36596 38292
rect 37004 38344 37056 38350
rect 37004 38286 37056 38292
rect 36360 38276 36412 38282
rect 36360 38218 36412 38224
rect 36372 37466 36400 38218
rect 36452 38208 36504 38214
rect 36452 38150 36504 38156
rect 36360 37460 36412 37466
rect 36360 37402 36412 37408
rect 36464 37330 36492 38150
rect 36556 37670 36584 38286
rect 36544 37664 36596 37670
rect 36544 37606 36596 37612
rect 36452 37324 36504 37330
rect 36452 37266 36504 37272
rect 36174 37224 36230 37233
rect 36174 37159 36230 37168
rect 36188 36786 36216 37159
rect 36556 36854 36584 37606
rect 36820 37460 36872 37466
rect 36820 37402 36872 37408
rect 36544 36848 36596 36854
rect 36544 36790 36596 36796
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 35768 36672 35848 36700
rect 35716 36654 35768 36660
rect 36176 36576 36228 36582
rect 36176 36518 36228 36524
rect 35532 36372 35584 36378
rect 35532 36314 35584 36320
rect 35716 36100 35768 36106
rect 35716 36042 35768 36048
rect 34756 35992 34836 36020
rect 34704 35974 34756 35980
rect 34612 35828 34664 35834
rect 34612 35770 34664 35776
rect 34716 35698 34744 35974
rect 35728 35834 35756 36042
rect 35716 35828 35768 35834
rect 35716 35770 35768 35776
rect 34704 35692 34756 35698
rect 34704 35634 34756 35640
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35728 35290 35756 35770
rect 35716 35284 35768 35290
rect 35716 35226 35768 35232
rect 36188 34950 36216 36518
rect 36176 34944 36228 34950
rect 36176 34886 36228 34892
rect 36268 34944 36320 34950
rect 36268 34886 36320 34892
rect 36188 34592 36216 34886
rect 36280 34746 36308 34886
rect 36268 34740 36320 34746
rect 36268 34682 36320 34688
rect 36832 34610 36860 37402
rect 37004 37324 37056 37330
rect 37004 37266 37056 37272
rect 36544 34604 36596 34610
rect 36188 34564 36544 34592
rect 36544 34546 36596 34552
rect 36820 34604 36872 34610
rect 36820 34546 36872 34552
rect 34520 34536 34572 34542
rect 34520 34478 34572 34484
rect 34336 32904 34388 32910
rect 34336 32846 34388 32852
rect 33876 32836 33928 32842
rect 33876 32778 33928 32784
rect 34060 32836 34112 32842
rect 34060 32778 34112 32784
rect 33784 32564 33836 32570
rect 33784 32506 33836 32512
rect 33600 32496 33652 32502
rect 33600 32438 33652 32444
rect 33416 32428 33468 32434
rect 33416 32370 33468 32376
rect 33336 32286 33456 32314
rect 33232 32020 33284 32026
rect 33232 31962 33284 31968
rect 33048 31204 33100 31210
rect 33048 31146 33100 31152
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32968 30122 32996 30670
rect 32956 30116 33008 30122
rect 32956 30058 33008 30064
rect 32968 29850 32996 30058
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 33060 28626 33088 31146
rect 33324 30796 33376 30802
rect 33324 30738 33376 30744
rect 33336 30394 33364 30738
rect 33324 30388 33376 30394
rect 33324 30330 33376 30336
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33140 30048 33192 30054
rect 33140 29990 33192 29996
rect 33152 29306 33180 29990
rect 33336 29850 33364 30194
rect 33324 29844 33376 29850
rect 33324 29786 33376 29792
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 33244 29170 33272 29446
rect 33336 29170 33364 29514
rect 33232 29164 33284 29170
rect 33232 29106 33284 29112
rect 33324 29164 33376 29170
rect 33324 29106 33376 29112
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 33152 28558 33180 28902
rect 33428 28694 33456 32286
rect 33784 32224 33836 32230
rect 33784 32166 33836 32172
rect 33508 31340 33560 31346
rect 33508 31282 33560 31288
rect 33600 31340 33652 31346
rect 33600 31282 33652 31288
rect 33520 30938 33548 31282
rect 33508 30932 33560 30938
rect 33508 30874 33560 30880
rect 33508 30320 33560 30326
rect 33508 30262 33560 30268
rect 33520 29850 33548 30262
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33612 29730 33640 31282
rect 33520 29702 33640 29730
rect 33520 29170 33548 29702
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33612 29306 33640 29582
rect 33600 29300 33652 29306
rect 33600 29242 33652 29248
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33416 28688 33468 28694
rect 33416 28630 33468 28636
rect 33140 28552 33192 28558
rect 33140 28494 33192 28500
rect 33416 26512 33468 26518
rect 33416 26454 33468 26460
rect 33140 26444 33192 26450
rect 33140 26386 33192 26392
rect 33152 26042 33180 26386
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33140 26036 33192 26042
rect 33140 25978 33192 25984
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 33060 25106 33088 25774
rect 33336 25294 33364 26318
rect 33428 25498 33456 26454
rect 33416 25492 33468 25498
rect 33416 25434 33468 25440
rect 33416 25356 33468 25362
rect 33416 25298 33468 25304
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33140 25152 33192 25158
rect 33060 25100 33140 25106
rect 33060 25094 33192 25100
rect 33060 25078 33180 25094
rect 32864 24336 32916 24342
rect 32864 24278 32916 24284
rect 33060 24206 33088 25078
rect 33336 24954 33364 25230
rect 33324 24948 33376 24954
rect 33324 24890 33376 24896
rect 33428 24818 33456 25298
rect 33416 24812 33468 24818
rect 33416 24754 33468 24760
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33048 24200 33100 24206
rect 33048 24142 33100 24148
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32772 24064 32824 24070
rect 32772 24006 32824 24012
rect 32692 23798 32720 24006
rect 32784 23798 32812 24006
rect 32680 23792 32732 23798
rect 32680 23734 32732 23740
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 33060 23730 33088 24142
rect 33244 23798 33272 24686
rect 33520 24274 33548 29106
rect 33796 28558 33824 32166
rect 33888 31482 33916 32778
rect 34348 31754 34376 32846
rect 34532 32842 34560 34478
rect 37016 34474 37044 37266
rect 37200 36106 37228 39306
rect 38028 38758 38056 39374
rect 38304 38826 38332 39374
rect 38752 39364 38804 39370
rect 38752 39306 38804 39312
rect 38660 38956 38712 38962
rect 38660 38898 38712 38904
rect 38292 38820 38344 38826
rect 38292 38762 38344 38768
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 38016 38752 38068 38758
rect 38016 38694 38068 38700
rect 37292 38350 37320 38694
rect 38304 38418 38332 38762
rect 38672 38593 38700 38898
rect 38764 38758 38792 39306
rect 38752 38752 38804 38758
rect 38752 38694 38804 38700
rect 38658 38584 38714 38593
rect 38658 38519 38714 38528
rect 38292 38412 38344 38418
rect 38292 38354 38344 38360
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 37292 37806 37320 38286
rect 38292 37868 38344 37874
rect 38292 37810 38344 37816
rect 37280 37800 37332 37806
rect 37280 37742 37332 37748
rect 37372 37800 37424 37806
rect 37372 37742 37424 37748
rect 37280 37120 37332 37126
rect 37384 37074 37412 37742
rect 37648 37664 37700 37670
rect 37648 37606 37700 37612
rect 37332 37068 37412 37074
rect 37280 37062 37412 37068
rect 37292 37046 37412 37062
rect 37292 36582 37320 37046
rect 37660 36854 37688 37606
rect 38304 37466 38332 37810
rect 38568 37800 38620 37806
rect 38568 37742 38620 37748
rect 38292 37460 38344 37466
rect 38292 37402 38344 37408
rect 38016 37256 38068 37262
rect 38016 37198 38068 37204
rect 38028 36922 38056 37198
rect 38304 37194 38332 37402
rect 38292 37188 38344 37194
rect 38292 37130 38344 37136
rect 38384 37188 38436 37194
rect 38384 37130 38436 37136
rect 38016 36916 38068 36922
rect 38016 36858 38068 36864
rect 37648 36848 37700 36854
rect 37648 36790 37700 36796
rect 37280 36576 37332 36582
rect 37280 36518 37332 36524
rect 37740 36576 37792 36582
rect 37740 36518 37792 36524
rect 38292 36576 38344 36582
rect 38292 36518 38344 36524
rect 37188 36100 37240 36106
rect 37188 36042 37240 36048
rect 37200 35766 37228 36042
rect 37188 35760 37240 35766
rect 37188 35702 37240 35708
rect 37188 35080 37240 35086
rect 37188 35022 37240 35028
rect 37096 34536 37148 34542
rect 37096 34478 37148 34484
rect 37004 34468 37056 34474
rect 37004 34410 37056 34416
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 37016 34202 37044 34410
rect 37004 34196 37056 34202
rect 37004 34138 37056 34144
rect 37016 34082 37044 34138
rect 36924 34054 37044 34082
rect 35900 33856 35952 33862
rect 35900 33798 35952 33804
rect 36636 33856 36688 33862
rect 36636 33798 36688 33804
rect 35532 33652 35584 33658
rect 35532 33594 35584 33600
rect 34796 33448 34848 33454
rect 34796 33390 34848 33396
rect 34808 33114 34836 33390
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 35544 33046 35572 33594
rect 35912 33522 35940 33798
rect 35900 33516 35952 33522
rect 35900 33458 35952 33464
rect 35992 33448 36044 33454
rect 35992 33390 36044 33396
rect 36004 33114 36032 33390
rect 36544 33312 36596 33318
rect 36544 33254 36596 33260
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 35532 33040 35584 33046
rect 35532 32982 35584 32988
rect 34520 32836 34572 32842
rect 34520 32778 34572 32784
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 34072 31726 34376 31754
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33980 31482 34008 31622
rect 33876 31476 33928 31482
rect 33876 31418 33928 31424
rect 33968 31476 34020 31482
rect 33968 31418 34020 31424
rect 34072 31346 34100 31726
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 33876 31136 33928 31142
rect 33876 31078 33928 31084
rect 33888 30938 33916 31078
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 34072 29102 34100 31282
rect 34808 30734 34836 31758
rect 35544 31346 35572 32982
rect 35636 32978 35756 32994
rect 35636 32972 35768 32978
rect 35636 32966 35716 32972
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 35440 31204 35492 31210
rect 35440 31146 35492 31152
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30734 35480 31146
rect 35636 31142 35664 32966
rect 35716 32914 35768 32920
rect 35900 31952 35952 31958
rect 35900 31894 35952 31900
rect 35624 31136 35676 31142
rect 35624 31078 35676 31084
rect 35636 30734 35664 31078
rect 35912 30802 35940 31894
rect 36556 31890 36584 33254
rect 36648 32842 36676 33798
rect 36820 33516 36872 33522
rect 36820 33458 36872 33464
rect 36636 32836 36688 32842
rect 36636 32778 36688 32784
rect 36832 32230 36860 33458
rect 36924 33114 36952 34054
rect 37004 33992 37056 33998
rect 37004 33934 37056 33940
rect 37016 33318 37044 33934
rect 37004 33312 37056 33318
rect 37004 33254 37056 33260
rect 37108 33114 37136 34478
rect 37200 33590 37228 35022
rect 37292 34066 37320 36518
rect 37752 36038 37780 36518
rect 37740 36032 37792 36038
rect 37740 35974 37792 35980
rect 37752 35630 37780 35974
rect 37924 35828 37976 35834
rect 37924 35770 37976 35776
rect 37740 35624 37792 35630
rect 37740 35566 37792 35572
rect 37372 34672 37424 34678
rect 37372 34614 37424 34620
rect 37280 34060 37332 34066
rect 37280 34002 37332 34008
rect 37280 33856 37332 33862
rect 37280 33798 37332 33804
rect 37188 33584 37240 33590
rect 37188 33526 37240 33532
rect 36912 33108 36964 33114
rect 36912 33050 36964 33056
rect 37096 33108 37148 33114
rect 37096 33050 37148 33056
rect 37292 32910 37320 33798
rect 37384 32910 37412 34614
rect 37936 34610 37964 35770
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 37648 34060 37700 34066
rect 37648 34002 37700 34008
rect 37660 33590 37688 34002
rect 38028 33930 38056 34886
rect 38304 34610 38332 36518
rect 38396 35834 38424 37130
rect 38580 36938 38608 37742
rect 38764 37670 38792 38694
rect 39132 38554 39160 39918
rect 39304 39500 39356 39506
rect 39304 39442 39356 39448
rect 39316 38593 39344 39442
rect 39856 39432 39908 39438
rect 39856 39374 39908 39380
rect 39488 39296 39540 39302
rect 39488 39238 39540 39244
rect 39396 39024 39448 39030
rect 39396 38966 39448 38972
rect 39302 38584 39358 38593
rect 39120 38548 39172 38554
rect 39302 38519 39358 38528
rect 39120 38490 39172 38496
rect 39212 38412 39264 38418
rect 39212 38354 39264 38360
rect 38936 38208 38988 38214
rect 38936 38150 38988 38156
rect 38948 37874 38976 38150
rect 38936 37868 38988 37874
rect 38936 37810 38988 37816
rect 39120 37868 39172 37874
rect 39120 37810 39172 37816
rect 38752 37664 38804 37670
rect 38752 37606 38804 37612
rect 39132 37466 39160 37810
rect 39120 37460 39172 37466
rect 39120 37402 39172 37408
rect 39224 37194 39252 38354
rect 39316 38350 39344 38519
rect 39304 38344 39356 38350
rect 39304 38286 39356 38292
rect 39316 37874 39344 38286
rect 39304 37868 39356 37874
rect 39304 37810 39356 37816
rect 39316 37466 39344 37810
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 39408 37210 39436 38966
rect 39500 38654 39528 39238
rect 39868 38962 39896 39374
rect 40132 39364 40184 39370
rect 40132 39306 40184 39312
rect 40040 39296 40092 39302
rect 40040 39238 40092 39244
rect 39856 38956 39908 38962
rect 39856 38898 39908 38904
rect 39764 38888 39816 38894
rect 39764 38830 39816 38836
rect 39500 38626 39620 38654
rect 39592 38282 39620 38626
rect 39776 38486 39804 38830
rect 39764 38480 39816 38486
rect 39764 38422 39816 38428
rect 39580 38276 39632 38282
rect 39580 38218 39632 38224
rect 39592 37942 39620 38218
rect 39580 37936 39632 37942
rect 39580 37878 39632 37884
rect 39672 37664 39724 37670
rect 39672 37606 39724 37612
rect 39408 37194 39620 37210
rect 39212 37188 39264 37194
rect 39408 37188 39632 37194
rect 39408 37182 39580 37188
rect 39212 37130 39264 37136
rect 39580 37130 39632 37136
rect 38660 37120 38712 37126
rect 38660 37062 38712 37068
rect 38488 36922 38608 36938
rect 38476 36916 38608 36922
rect 38528 36910 38608 36916
rect 38672 36938 38700 37062
rect 38672 36910 38792 36938
rect 38476 36858 38528 36864
rect 38764 36242 38792 36910
rect 39224 36854 39252 37130
rect 39488 37120 39540 37126
rect 39488 37062 39540 37068
rect 39500 36854 39528 37062
rect 39684 36854 39712 37606
rect 39212 36848 39264 36854
rect 39212 36790 39264 36796
rect 39488 36848 39540 36854
rect 39488 36790 39540 36796
rect 39672 36848 39724 36854
rect 39672 36790 39724 36796
rect 39224 36378 39252 36790
rect 39212 36372 39264 36378
rect 39212 36314 39264 36320
rect 38752 36236 38804 36242
rect 38752 36178 38804 36184
rect 39224 36106 39252 36314
rect 39212 36100 39264 36106
rect 39212 36042 39264 36048
rect 38384 35828 38436 35834
rect 38384 35770 38436 35776
rect 38476 35624 38528 35630
rect 38476 35566 38528 35572
rect 38488 34610 38516 35566
rect 39224 35442 39252 36042
rect 39224 35414 39344 35442
rect 38660 35080 38712 35086
rect 38660 35022 38712 35028
rect 38672 34746 38700 35022
rect 39316 35018 39344 35414
rect 39304 35012 39356 35018
rect 39304 34954 39356 34960
rect 38752 34944 38804 34950
rect 38752 34886 38804 34892
rect 38660 34740 38712 34746
rect 38660 34682 38712 34688
rect 38764 34610 38792 34886
rect 38844 34672 38896 34678
rect 38844 34614 38896 34620
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 38476 34604 38528 34610
rect 38476 34546 38528 34552
rect 38752 34604 38804 34610
rect 38752 34546 38804 34552
rect 38108 34400 38160 34406
rect 38108 34342 38160 34348
rect 38016 33924 38068 33930
rect 38016 33866 38068 33872
rect 37648 33584 37700 33590
rect 37648 33526 37700 33532
rect 37280 32904 37332 32910
rect 37280 32846 37332 32852
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 36636 32224 36688 32230
rect 36636 32166 36688 32172
rect 36820 32224 36872 32230
rect 36820 32166 36872 32172
rect 36648 31890 36676 32166
rect 36544 31884 36596 31890
rect 36544 31826 36596 31832
rect 36636 31884 36688 31890
rect 36636 31826 36688 31832
rect 36832 31754 36860 32166
rect 37660 31754 37688 33526
rect 38120 33454 38148 34342
rect 38304 33862 38332 34546
rect 38384 34468 38436 34474
rect 38384 34410 38436 34416
rect 38396 34066 38424 34410
rect 38384 34060 38436 34066
rect 38384 34002 38436 34008
rect 38292 33856 38344 33862
rect 38292 33798 38344 33804
rect 38304 33454 38332 33798
rect 38108 33448 38160 33454
rect 38108 33390 38160 33396
rect 38292 33448 38344 33454
rect 38292 33390 38344 33396
rect 38016 32768 38068 32774
rect 38016 32710 38068 32716
rect 38028 31754 38056 32710
rect 38764 31890 38792 34546
rect 38856 33862 38884 34614
rect 39120 34536 39172 34542
rect 39120 34478 39172 34484
rect 39028 33992 39080 33998
rect 39028 33934 39080 33940
rect 38844 33856 38896 33862
rect 38844 33798 38896 33804
rect 38856 33522 38884 33798
rect 39040 33590 39068 33934
rect 39028 33584 39080 33590
rect 39028 33526 39080 33532
rect 39132 33538 39160 34478
rect 38844 33516 38896 33522
rect 38844 33458 38896 33464
rect 39040 33402 39068 33526
rect 39132 33510 39252 33538
rect 39500 33522 39528 36790
rect 39776 36718 39804 38422
rect 39868 37126 39896 38898
rect 40052 38418 40080 39238
rect 40040 38412 40092 38418
rect 40040 38354 40092 38360
rect 40144 38026 40172 39306
rect 40224 38888 40276 38894
rect 40224 38830 40276 38836
rect 40236 38554 40264 38830
rect 40224 38548 40276 38554
rect 40224 38490 40276 38496
rect 40512 38350 40540 40054
rect 40684 40044 40736 40050
rect 40684 39986 40736 39992
rect 40696 39370 40724 39986
rect 41788 39432 41840 39438
rect 41788 39374 41840 39380
rect 40684 39364 40736 39370
rect 40684 39306 40736 39312
rect 40696 39030 40724 39306
rect 41696 39296 41748 39302
rect 41696 39238 41748 39244
rect 40684 39024 40736 39030
rect 40684 38966 40736 38972
rect 40696 38418 40724 38966
rect 40684 38412 40736 38418
rect 40684 38354 40736 38360
rect 40316 38344 40368 38350
rect 40316 38286 40368 38292
rect 40500 38344 40552 38350
rect 40500 38286 40552 38292
rect 40224 38276 40276 38282
rect 40224 38218 40276 38224
rect 40052 38010 40172 38026
rect 40040 38004 40172 38010
rect 40092 37998 40172 38004
rect 40040 37946 40092 37952
rect 40132 37868 40184 37874
rect 40236 37856 40264 38218
rect 40184 37828 40264 37856
rect 40132 37810 40184 37816
rect 40328 37806 40356 38286
rect 41328 38208 41380 38214
rect 41328 38150 41380 38156
rect 40316 37800 40368 37806
rect 40316 37742 40368 37748
rect 39948 37188 40000 37194
rect 39948 37130 40000 37136
rect 39856 37120 39908 37126
rect 39856 37062 39908 37068
rect 39868 36922 39896 37062
rect 39856 36916 39908 36922
rect 39856 36858 39908 36864
rect 39764 36712 39816 36718
rect 39764 36654 39816 36660
rect 39776 34746 39804 36654
rect 39868 36242 39896 36858
rect 39856 36236 39908 36242
rect 39856 36178 39908 36184
rect 39764 34740 39816 34746
rect 39764 34682 39816 34688
rect 39580 34536 39632 34542
rect 39580 34478 39632 34484
rect 39592 33862 39620 34478
rect 39960 33930 39988 37130
rect 41340 36786 41368 38150
rect 41708 37874 41736 39238
rect 41800 38758 41828 39374
rect 41788 38752 41840 38758
rect 41788 38694 41840 38700
rect 41800 37874 41828 38694
rect 41880 38004 41932 38010
rect 41880 37946 41932 37952
rect 41696 37868 41748 37874
rect 41696 37810 41748 37816
rect 41788 37868 41840 37874
rect 41788 37810 41840 37816
rect 41512 37664 41564 37670
rect 41512 37606 41564 37612
rect 41328 36780 41380 36786
rect 41328 36722 41380 36728
rect 41420 36780 41472 36786
rect 41420 36722 41472 36728
rect 40316 36576 40368 36582
rect 40316 36518 40368 36524
rect 41328 36576 41380 36582
rect 41328 36518 41380 36524
rect 40328 36378 40356 36518
rect 40316 36372 40368 36378
rect 40316 36314 40368 36320
rect 40224 36236 40276 36242
rect 40224 36178 40276 36184
rect 40236 35154 40264 36178
rect 41340 35986 41368 36518
rect 41432 35986 41460 36722
rect 41524 36582 41552 37606
rect 41892 36786 41920 37946
rect 41604 36780 41656 36786
rect 41604 36722 41656 36728
rect 41880 36780 41932 36786
rect 41880 36722 41932 36728
rect 41512 36576 41564 36582
rect 41512 36518 41564 36524
rect 41340 35958 41460 35986
rect 41432 35714 41460 35958
rect 41524 35894 41552 36518
rect 41616 36038 41644 36722
rect 41696 36576 41748 36582
rect 41696 36518 41748 36524
rect 41708 36378 41736 36518
rect 41696 36372 41748 36378
rect 41696 36314 41748 36320
rect 41604 36032 41656 36038
rect 41604 35974 41656 35980
rect 41984 35894 42012 45834
rect 45284 44396 45336 44402
rect 45284 44338 45336 44344
rect 44364 44328 44416 44334
rect 45296 44305 45324 44338
rect 44364 44270 44416 44276
rect 45282 44296 45338 44305
rect 42064 39500 42116 39506
rect 42064 39442 42116 39448
rect 42076 38350 42104 39442
rect 42064 38344 42116 38350
rect 42064 38286 42116 38292
rect 42076 37738 42104 38286
rect 43260 37868 43312 37874
rect 43260 37810 43312 37816
rect 42064 37732 42116 37738
rect 42064 37674 42116 37680
rect 42800 37732 42852 37738
rect 42800 37674 42852 37680
rect 42076 36786 42104 37674
rect 42432 37256 42484 37262
rect 42432 37198 42484 37204
rect 42444 36786 42472 37198
rect 42812 36854 42840 37674
rect 43076 37664 43128 37670
rect 43076 37606 43128 37612
rect 43088 37330 43116 37606
rect 43076 37324 43128 37330
rect 43076 37266 43128 37272
rect 42800 36848 42852 36854
rect 42800 36790 42852 36796
rect 42064 36780 42116 36786
rect 42064 36722 42116 36728
rect 42432 36780 42484 36786
rect 42432 36722 42484 36728
rect 42708 36712 42760 36718
rect 42708 36654 42760 36660
rect 42720 36378 42748 36654
rect 42708 36372 42760 36378
rect 42708 36314 42760 36320
rect 42064 36032 42116 36038
rect 42064 35974 42116 35980
rect 41524 35866 41736 35894
rect 41432 35686 41644 35714
rect 41512 35624 41564 35630
rect 41512 35566 41564 35572
rect 40960 35488 41012 35494
rect 40960 35430 41012 35436
rect 40972 35154 41000 35430
rect 40224 35148 40276 35154
rect 40224 35090 40276 35096
rect 40960 35148 41012 35154
rect 40960 35090 41012 35096
rect 40040 35080 40092 35086
rect 40040 35022 40092 35028
rect 40052 34202 40080 35022
rect 41524 34746 41552 35566
rect 41512 34740 41564 34746
rect 41512 34682 41564 34688
rect 40592 34672 40644 34678
rect 40592 34614 40644 34620
rect 40408 34400 40460 34406
rect 40408 34342 40460 34348
rect 40040 34196 40092 34202
rect 40040 34138 40092 34144
rect 40420 33998 40448 34342
rect 40408 33992 40460 33998
rect 40408 33934 40460 33940
rect 39948 33924 40000 33930
rect 39948 33866 40000 33872
rect 39580 33856 39632 33862
rect 39580 33798 39632 33804
rect 39040 33374 39160 33402
rect 39028 33312 39080 33318
rect 39028 33254 39080 33260
rect 39040 32978 39068 33254
rect 39028 32972 39080 32978
rect 39028 32914 39080 32920
rect 38660 31884 38712 31890
rect 38660 31826 38712 31832
rect 38752 31884 38804 31890
rect 38752 31826 38804 31832
rect 38672 31754 38700 31826
rect 36832 31726 36952 31754
rect 37660 31726 37780 31754
rect 38028 31726 38148 31754
rect 38672 31726 38792 31754
rect 36452 31680 36504 31686
rect 36452 31622 36504 31628
rect 36360 31340 36412 31346
rect 36360 31282 36412 31288
rect 35900 30796 35952 30802
rect 35900 30738 35952 30744
rect 34796 30728 34848 30734
rect 34796 30670 34848 30676
rect 35440 30728 35492 30734
rect 35440 30670 35492 30676
rect 35624 30728 35676 30734
rect 35624 30670 35676 30676
rect 34152 30116 34204 30122
rect 34152 30058 34204 30064
rect 34164 29510 34192 30058
rect 34336 30048 34388 30054
rect 34336 29990 34388 29996
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34164 29238 34192 29446
rect 34152 29232 34204 29238
rect 34152 29174 34204 29180
rect 34060 29096 34112 29102
rect 34060 29038 34112 29044
rect 33876 28688 33928 28694
rect 33876 28630 33928 28636
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33888 28490 33916 28630
rect 33876 28484 33928 28490
rect 33876 28426 33928 28432
rect 33600 26240 33652 26246
rect 33600 26182 33652 26188
rect 33968 26240 34020 26246
rect 33968 26182 34020 26188
rect 33612 25430 33640 26182
rect 33980 25906 34008 26182
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 33600 25424 33652 25430
rect 33600 25366 33652 25372
rect 33612 24750 33640 25366
rect 34072 25294 34100 29038
rect 34164 28558 34192 29174
rect 34348 28558 34376 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35636 29714 35664 30670
rect 36372 30666 36400 31282
rect 36464 30802 36492 31622
rect 36452 30796 36504 30802
rect 36452 30738 36504 30744
rect 36360 30660 36412 30666
rect 36360 30602 36412 30608
rect 35624 29708 35676 29714
rect 35624 29650 35676 29656
rect 36372 29578 36400 30602
rect 35624 29572 35676 29578
rect 35624 29514 35676 29520
rect 36360 29572 36412 29578
rect 36360 29514 36412 29520
rect 35636 29306 35664 29514
rect 35624 29300 35676 29306
rect 35624 29242 35676 29248
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 34808 28762 34836 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 35624 28688 35676 28694
rect 35624 28630 35676 28636
rect 34520 28620 34572 28626
rect 34520 28562 34572 28568
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 34336 28552 34388 28558
rect 34336 28494 34388 28500
rect 34532 27674 34560 28562
rect 34612 28484 34664 28490
rect 34612 28426 34664 28432
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34624 27538 34652 28426
rect 34704 28076 34756 28082
rect 34704 28018 34756 28024
rect 35256 28076 35308 28082
rect 35256 28018 35308 28024
rect 35440 28076 35492 28082
rect 35440 28018 35492 28024
rect 34612 27532 34664 27538
rect 34612 27474 34664 27480
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 34348 27130 34376 27406
rect 34716 27334 34744 28018
rect 34796 27872 34848 27878
rect 34796 27814 34848 27820
rect 35268 27826 35296 28018
rect 35452 27826 35480 28018
rect 34808 27606 34836 27814
rect 35268 27798 35480 27826
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27600 34848 27606
rect 35360 27554 35388 27798
rect 34796 27542 34848 27548
rect 35176 27526 35388 27554
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34336 27124 34388 27130
rect 34336 27066 34388 27072
rect 34428 26920 34480 26926
rect 34428 26862 34480 26868
rect 34440 26364 34468 26862
rect 34716 26586 34744 27270
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34612 26376 34664 26382
rect 34440 26336 34612 26364
rect 34612 26318 34664 26324
rect 34808 26246 34836 26930
rect 35176 26858 35204 27526
rect 35256 27464 35308 27470
rect 35256 27406 35308 27412
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 35268 27130 35296 27406
rect 35256 27124 35308 27130
rect 35256 27066 35308 27072
rect 35164 26852 35216 26858
rect 35164 26794 35216 26800
rect 35268 26738 35296 27066
rect 35452 26926 35480 27406
rect 35636 27062 35664 28630
rect 36084 28620 36136 28626
rect 36084 28562 36136 28568
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35912 27878 35940 28494
rect 35992 28416 36044 28422
rect 35992 28358 36044 28364
rect 35900 27872 35952 27878
rect 35900 27814 35952 27820
rect 35912 27470 35940 27814
rect 35900 27464 35952 27470
rect 35900 27406 35952 27412
rect 35624 27056 35676 27062
rect 35624 26998 35676 27004
rect 35440 26920 35492 26926
rect 35440 26862 35492 26868
rect 35268 26710 35388 26738
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26586 35388 26710
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 35348 26308 35400 26314
rect 35452 26296 35480 26862
rect 35400 26268 35480 26296
rect 35348 26250 35400 26256
rect 34152 26240 34204 26246
rect 34152 26182 34204 26188
rect 34796 26240 34848 26246
rect 34796 26182 34848 26188
rect 34164 25906 34192 26182
rect 34152 25900 34204 25906
rect 34152 25842 34204 25848
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 33876 25220 33928 25226
rect 33876 25162 33928 25168
rect 33968 25220 34020 25226
rect 33968 25162 34020 25168
rect 33888 24954 33916 25162
rect 33980 24954 34008 25162
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 33968 24948 34020 24954
rect 33968 24890 34020 24896
rect 34072 24886 34100 25230
rect 34808 25158 34836 26182
rect 35360 25838 35388 26250
rect 35348 25832 35400 25838
rect 35348 25774 35400 25780
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34980 25152 35032 25158
rect 34980 25094 35032 25100
rect 34060 24880 34112 24886
rect 34060 24822 34112 24828
rect 34992 24818 35020 25094
rect 35440 24880 35492 24886
rect 35440 24822 35492 24828
rect 34980 24812 35032 24818
rect 34980 24754 35032 24760
rect 33600 24744 33652 24750
rect 33600 24686 33652 24692
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33508 24268 33560 24274
rect 33508 24210 33560 24216
rect 33692 24064 33744 24070
rect 33692 24006 33744 24012
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 33232 23792 33284 23798
rect 33232 23734 33284 23740
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 32772 23656 32824 23662
rect 32772 23598 32824 23604
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 32588 23112 32640 23118
rect 32588 23054 32640 23060
rect 32600 22778 32628 23054
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32784 22574 32812 23598
rect 33428 23322 33456 23598
rect 33416 23316 33468 23322
rect 33416 23258 33468 23264
rect 33704 23186 33732 24006
rect 35360 23866 35388 24006
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 33048 23112 33100 23118
rect 33048 23054 33100 23060
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 33060 22710 33088 23054
rect 33048 22704 33100 22710
rect 33048 22646 33100 22652
rect 32772 22568 32824 22574
rect 32772 22510 32824 22516
rect 34060 22432 34112 22438
rect 34060 22374 34112 22380
rect 34072 21962 34100 22374
rect 34152 22228 34204 22234
rect 34152 22170 34204 22176
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32220 20460 32272 20466
rect 32220 20402 32272 20408
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32232 20058 32260 20402
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32220 20052 32272 20058
rect 32220 19994 32272 20000
rect 32324 19961 32352 20334
rect 32416 20058 32444 20402
rect 32404 20052 32456 20058
rect 32404 19994 32456 20000
rect 32508 19990 32536 20402
rect 32772 20392 32824 20398
rect 32772 20334 32824 20340
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 32496 19984 32548 19990
rect 32310 19952 32366 19961
rect 32496 19926 32548 19932
rect 32310 19887 32366 19896
rect 32324 19854 32352 19887
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 32048 18290 32076 18634
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 32140 17898 32168 19246
rect 32220 18896 32272 18902
rect 32404 18896 32456 18902
rect 32272 18856 32404 18884
rect 32220 18838 32272 18844
rect 32404 18838 32456 18844
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32324 18426 32352 18702
rect 32508 18698 32536 19926
rect 32600 19854 32628 20198
rect 32588 19848 32640 19854
rect 32588 19790 32640 19796
rect 32784 18766 32812 20334
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 19310 33088 19654
rect 33874 19408 33930 19417
rect 33416 19372 33468 19378
rect 33874 19343 33876 19352
rect 33416 19314 33468 19320
rect 33928 19343 33930 19352
rect 33876 19314 33928 19320
rect 33048 19304 33100 19310
rect 33048 19246 33100 19252
rect 33060 18970 33088 19246
rect 33428 18970 33456 19314
rect 33048 18964 33100 18970
rect 33048 18906 33100 18912
rect 33416 18964 33468 18970
rect 33416 18906 33468 18912
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 32140 17882 32260 17898
rect 32140 17876 32272 17882
rect 32140 17870 32220 17876
rect 32220 17818 32272 17824
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 32140 17270 32168 17546
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 31944 16720 31996 16726
rect 31944 16662 31996 16668
rect 32232 16114 32260 17818
rect 32416 17746 32444 18566
rect 32600 18358 32628 18566
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 33612 18222 33640 18566
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33612 17882 33640 18158
rect 33600 17876 33652 17882
rect 33600 17818 33652 17824
rect 33704 17746 33732 18566
rect 34072 18222 34100 18634
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 32404 17740 32456 17746
rect 32404 17682 32456 17688
rect 33692 17740 33744 17746
rect 33692 17682 33744 17688
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32876 16182 32904 17546
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 32956 16448 33008 16454
rect 32956 16390 33008 16396
rect 32968 16250 32996 16390
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 32864 16176 32916 16182
rect 32864 16118 32916 16124
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31668 16108 31720 16114
rect 31668 16050 31720 16056
rect 32220 16108 32272 16114
rect 32220 16050 32272 16056
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29012 15706 29040 15846
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 29012 15026 29040 15642
rect 29380 15502 29408 15846
rect 30576 15706 30604 16050
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 29644 15564 29696 15570
rect 29644 15506 29696 15512
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29380 14618 29408 15438
rect 29656 15026 29684 15506
rect 30024 15026 30052 15642
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30300 15026 30328 15438
rect 30484 15026 30512 15438
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30576 15026 30604 15302
rect 30760 15162 30788 15846
rect 31220 15502 31248 16050
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 31496 15502 31524 15982
rect 31680 15638 31708 16050
rect 33060 16046 33088 16526
rect 34164 16182 34192 22170
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 19378 34468 19654
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34348 18426 34376 18702
rect 34336 18420 34388 18426
rect 34336 18362 34388 18368
rect 34532 17746 34560 23054
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34624 22710 34652 22918
rect 34612 22704 34664 22710
rect 34612 22646 34664 22652
rect 34704 19916 34756 19922
rect 34704 19858 34756 19864
rect 34716 19514 34744 19858
rect 34704 19508 34756 19514
rect 34624 19468 34704 19496
rect 34624 18766 34652 19468
rect 34704 19450 34756 19456
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34532 16658 34560 17682
rect 34520 16652 34572 16658
rect 34520 16594 34572 16600
rect 34152 16176 34204 16182
rect 34152 16118 34204 16124
rect 33048 16040 33100 16046
rect 33048 15982 33100 15988
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31852 15904 31904 15910
rect 31852 15846 31904 15852
rect 34060 15904 34112 15910
rect 34060 15846 34112 15852
rect 31668 15632 31720 15638
rect 31668 15574 31720 15580
rect 31772 15502 31800 15846
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 30748 15156 30800 15162
rect 30748 15098 30800 15104
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 29368 14612 29420 14618
rect 29368 14554 29420 14560
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 27264 13462 27292 14010
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 27252 13456 27304 13462
rect 27252 13398 27304 13404
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 27068 11688 27120 11694
rect 26988 11648 27068 11676
rect 27068 11630 27120 11636
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 25884 6866 25912 7278
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 25504 5704 25556 5710
rect 25556 5664 25728 5692
rect 25504 5646 25556 5652
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 25280 5052 25360 5080
rect 25228 5034 25280 5040
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 25424 4486 25452 5170
rect 25516 5166 25544 5510
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17512 3148 17632 3176
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17512 2990 17540 3148
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17592 2984 17644 2990
rect 17972 2972 18000 3334
rect 18156 3194 18184 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 25608 3194 25636 4082
rect 25700 3602 25728 5664
rect 25884 5098 25912 6802
rect 25976 6798 26004 7346
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 25976 5098 26004 6734
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26160 5914 26188 6054
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 26160 5574 26188 5850
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26160 5234 26188 5510
rect 26988 5370 27016 11494
rect 27080 10674 27108 11630
rect 27172 11234 27200 12786
rect 27264 11558 27292 12922
rect 27632 12646 27660 13126
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27724 12442 27752 13330
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27540 11354 27568 11766
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27172 11218 27292 11234
rect 27172 11212 27304 11218
rect 27172 11206 27252 11212
rect 27252 11154 27304 11160
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27080 9722 27108 10610
rect 27172 10198 27200 10610
rect 27160 10192 27212 10198
rect 27160 10134 27212 10140
rect 27264 10130 27292 11154
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27540 10470 27568 10610
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 28000 10266 28028 11698
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10674 28304 11018
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 27068 9716 27120 9722
rect 27068 9658 27120 9664
rect 27264 9518 27292 10066
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 27264 8430 27292 9454
rect 27356 9178 27384 9658
rect 27448 9382 27476 9998
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27356 9042 27384 9114
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27264 7002 27292 8366
rect 27356 8022 27384 8434
rect 27448 8362 27476 9318
rect 27540 9178 27568 9318
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27540 7954 27568 8910
rect 28000 8480 28028 10202
rect 28092 9178 28120 10542
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 28184 8906 28212 10406
rect 28368 9654 28396 12174
rect 28460 11218 28488 13126
rect 28920 12986 28948 13126
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 29012 12714 29040 13126
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 29104 12238 29132 13806
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29288 12986 29316 13262
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29472 12434 29500 14758
rect 30300 14618 30328 14758
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30012 14476 30064 14482
rect 30012 14418 30064 14424
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29656 12442 29684 12786
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 29380 12406 29500 12434
rect 29644 12436 29696 12442
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28828 11626 28856 12038
rect 29012 11762 29040 12174
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 28816 11620 28868 11626
rect 28816 11562 28868 11568
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 28552 11354 28580 11494
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28368 8974 28396 9590
rect 28460 9178 28488 11154
rect 28828 10674 28856 11562
rect 29012 11354 29040 11698
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28920 10690 28948 11086
rect 28920 10674 29132 10690
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28920 10668 29144 10674
rect 28920 10662 29092 10668
rect 28920 9722 28948 10662
rect 29092 10610 29144 10616
rect 29184 10600 29236 10606
rect 29184 10542 29236 10548
rect 29000 10532 29052 10538
rect 29000 10474 29052 10480
rect 29012 10266 29040 10474
rect 29196 10266 29224 10542
rect 29276 10464 29328 10470
rect 29276 10406 29328 10412
rect 29288 10266 29316 10406
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 29184 10260 29236 10266
rect 29184 10202 29236 10208
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29196 9994 29224 10202
rect 29184 9988 29236 9994
rect 29184 9930 29236 9936
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28448 9172 28500 9178
rect 28448 9114 28500 9120
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28184 8634 28212 8842
rect 28368 8634 28396 8910
rect 28460 8634 28488 9114
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28000 8452 28120 8480
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27344 7812 27396 7818
rect 27344 7754 27396 7760
rect 27356 7546 27384 7754
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27540 7342 27568 7890
rect 27908 7886 27936 8366
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27908 7546 27936 7822
rect 28092 7750 28120 8452
rect 28552 7886 28580 8910
rect 28920 8906 28948 9658
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 29184 8900 29236 8906
rect 29184 8842 29236 8848
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29012 8498 29040 8774
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29104 7954 29132 8570
rect 29196 8498 29224 8842
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28080 7744 28132 7750
rect 28080 7686 28132 7692
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27540 6798 27568 7278
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27080 5710 27108 6734
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 27160 5568 27212 5574
rect 27160 5510 27212 5516
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 26988 5234 27016 5306
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 25872 5092 25924 5098
rect 25872 5034 25924 5040
rect 25964 5092 26016 5098
rect 25964 5034 26016 5040
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25792 3738 25820 3878
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25976 3534 26004 5034
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26068 3194 26096 4082
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26528 3058 26556 3538
rect 27080 3194 27108 4082
rect 27172 3942 27200 5510
rect 27356 5098 27384 5578
rect 29012 5098 29040 5646
rect 27344 5092 27396 5098
rect 27344 5034 27396 5040
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28552 4078 28580 4558
rect 29012 4282 29040 5034
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28816 4072 28868 4078
rect 28816 4014 28868 4020
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27356 3194 27384 3878
rect 28552 3738 28580 4014
rect 28828 3738 28856 4014
rect 28540 3732 28592 3738
rect 28540 3674 28592 3680
rect 28816 3732 28868 3738
rect 28816 3674 28868 3680
rect 29012 3534 29040 4218
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 29012 3126 29040 3470
rect 29380 3194 29408 12406
rect 29644 12378 29696 12384
rect 29460 12232 29512 12238
rect 29460 12174 29512 12180
rect 29472 9994 29500 12174
rect 29840 11898 29868 12718
rect 29932 12170 29960 13126
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29828 11892 29880 11898
rect 29748 11852 29828 11880
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29656 10674 29684 10746
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29460 9988 29512 9994
rect 29460 9930 29512 9936
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 29656 9518 29684 9862
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29552 9444 29604 9450
rect 29552 9386 29604 9392
rect 29564 9217 29592 9386
rect 29550 9208 29606 9217
rect 29550 9143 29606 9152
rect 29656 8974 29684 9454
rect 29748 8974 29776 11852
rect 29828 11834 29880 11840
rect 30024 11778 30052 14418
rect 30380 14408 30432 14414
rect 30378 14376 30380 14385
rect 30484 14396 30512 14962
rect 31220 14958 31248 15438
rect 31496 15026 31524 15438
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 31208 14952 31260 14958
rect 31208 14894 31260 14900
rect 30432 14376 30512 14396
rect 30434 14368 30512 14376
rect 30378 14311 30434 14320
rect 31404 14006 31432 14962
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 30840 14000 30892 14006
rect 30840 13942 30892 13948
rect 31392 14000 31444 14006
rect 31392 13942 31444 13948
rect 30472 12776 30524 12782
rect 30472 12718 30524 12724
rect 30484 12434 30512 12718
rect 30748 12640 30800 12646
rect 30748 12582 30800 12588
rect 30760 12442 30788 12582
rect 30748 12436 30800 12442
rect 30484 12406 30696 12434
rect 30668 12238 30696 12406
rect 30748 12378 30800 12384
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 29932 11750 30052 11778
rect 29932 11150 29960 11750
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29840 10470 29868 10746
rect 29932 10674 29960 11086
rect 30024 10674 30052 11630
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 11354 30144 11494
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 30116 10674 30144 11290
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 30012 10668 30064 10674
rect 30012 10610 30064 10616
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 29840 8974 29868 10406
rect 29932 9761 29960 10610
rect 30024 10062 30052 10610
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 29918 9752 29974 9761
rect 29918 9687 29974 9696
rect 29932 9466 29960 9687
rect 30024 9586 30052 9998
rect 30300 9674 30328 12038
rect 30392 11830 30420 12174
rect 30576 11898 30604 12174
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30576 11354 30604 11698
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30668 10010 30696 12174
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30760 11257 30788 12106
rect 30746 11248 30802 11257
rect 30746 11183 30802 11192
rect 30760 11150 30788 11183
rect 30748 11144 30800 11150
rect 30748 11086 30800 11092
rect 30852 11098 30880 13942
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30944 13326 30972 13670
rect 31036 13462 31064 13874
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31024 13456 31076 13462
rect 31024 13398 31076 13404
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30852 11070 30972 11098
rect 30748 11008 30800 11014
rect 30748 10950 30800 10956
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30760 10198 30788 10950
rect 30852 10470 30880 10950
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30748 10192 30800 10198
rect 30748 10134 30800 10140
rect 30668 9982 30788 10010
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30300 9646 30512 9674
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 29932 9438 30052 9466
rect 29920 9376 29972 9382
rect 29920 9318 29972 9324
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29828 8968 29880 8974
rect 29932 8952 29960 9318
rect 29828 8910 29880 8916
rect 29920 8946 29972 8952
rect 29656 8838 29684 8910
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29656 8634 29684 8774
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29748 8090 29776 8910
rect 29840 8634 29868 8910
rect 29920 8888 29972 8894
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 30024 8498 30052 9438
rect 30104 9104 30156 9110
rect 30102 9072 30104 9081
rect 30156 9072 30158 9081
rect 30102 9007 30158 9016
rect 30208 8906 30236 9590
rect 30300 9586 30328 9646
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30286 9208 30342 9217
rect 30286 9143 30288 9152
rect 30340 9143 30342 9152
rect 30288 9114 30340 9120
rect 30484 9042 30512 9646
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30576 9382 30604 9454
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30196 8900 30248 8906
rect 30196 8842 30248 8848
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30300 8498 30328 8774
rect 30668 8498 30696 9522
rect 30760 8974 30788 9982
rect 30840 9104 30892 9110
rect 30838 9072 30840 9081
rect 30892 9072 30894 9081
rect 30838 9007 30894 9016
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30840 8900 30892 8906
rect 30840 8842 30892 8848
rect 30852 8634 30880 8842
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 30852 8498 30880 8570
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 30208 8090 30236 8434
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 30484 7818 30512 8230
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30944 6882 30972 11070
rect 31036 10810 31064 11698
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31036 8498 31064 9658
rect 31128 8922 31156 13670
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 31220 12238 31248 13398
rect 31300 12708 31352 12714
rect 31300 12650 31352 12656
rect 31312 12288 31340 12650
rect 31496 12424 31524 14758
rect 31588 14618 31616 15370
rect 31576 14612 31628 14618
rect 31576 14554 31628 14560
rect 31588 13462 31616 14554
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31772 13682 31800 14418
rect 31864 14346 31892 15846
rect 34072 15706 34100 15846
rect 34060 15700 34112 15706
rect 34060 15642 34112 15648
rect 32312 15428 32364 15434
rect 32312 15370 32364 15376
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31680 13654 31800 13682
rect 31576 13456 31628 13462
rect 31576 13398 31628 13404
rect 31588 12646 31616 13398
rect 31680 13326 31708 13654
rect 31864 13462 31892 14282
rect 32140 14074 32168 14350
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31852 13456 31904 13462
rect 31852 13398 31904 13404
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 31680 12764 31708 13262
rect 31772 12918 31800 13262
rect 31864 12986 31892 13398
rect 31956 13258 31984 13874
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31760 12912 31812 12918
rect 31760 12854 31812 12860
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 31760 12776 31812 12782
rect 31680 12736 31760 12764
rect 31576 12640 31628 12646
rect 31576 12582 31628 12588
rect 31496 12396 31616 12424
rect 31392 12300 31444 12306
rect 31312 12260 31392 12288
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 10198 31248 12038
rect 31312 11286 31340 12260
rect 31392 12242 31444 12248
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31404 11354 31432 12106
rect 31496 11762 31524 12174
rect 31588 11812 31616 12396
rect 31680 12238 31708 12736
rect 31760 12718 31812 12724
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31772 12238 31800 12582
rect 31864 12434 31892 12786
rect 32140 12434 32168 13262
rect 31864 12406 32076 12434
rect 32140 12406 32260 12434
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31588 11784 31708 11812
rect 31484 11756 31536 11762
rect 31536 11716 31616 11744
rect 31484 11698 31536 11704
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31300 11280 31352 11286
rect 31300 11222 31352 11228
rect 31404 11150 31432 11290
rect 31300 11144 31352 11150
rect 31392 11144 31444 11150
rect 31300 11086 31352 11092
rect 31390 11112 31392 11121
rect 31444 11112 31446 11121
rect 31312 10266 31340 11086
rect 31390 11047 31446 11056
rect 31588 10742 31616 11716
rect 31680 11286 31708 11784
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31668 11280 31720 11286
rect 31668 11222 31720 11228
rect 31680 10742 31708 11222
rect 31576 10736 31628 10742
rect 31576 10678 31628 10684
rect 31668 10736 31720 10742
rect 31668 10678 31720 10684
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31404 10266 31432 10610
rect 31484 10532 31536 10538
rect 31484 10474 31536 10480
rect 31300 10260 31352 10266
rect 31300 10202 31352 10208
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31208 10192 31260 10198
rect 31208 10134 31260 10140
rect 31300 10056 31352 10062
rect 31352 10004 31432 10010
rect 31300 9998 31432 10004
rect 31312 9982 31432 9998
rect 31300 9920 31352 9926
rect 31300 9862 31352 9868
rect 31312 9586 31340 9862
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 31404 9382 31432 9982
rect 31496 9722 31524 10474
rect 31588 10266 31616 10678
rect 31668 10464 31720 10470
rect 31668 10406 31720 10412
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31404 9178 31432 9318
rect 31392 9172 31444 9178
rect 31392 9114 31444 9120
rect 31588 9042 31616 10202
rect 31680 9926 31708 10406
rect 31772 10062 31800 11630
rect 31864 11218 31892 11698
rect 32048 11234 32076 12406
rect 32232 12238 32260 12406
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32140 11762 32168 12174
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 32232 11354 32260 11494
rect 32220 11348 32272 11354
rect 32220 11290 32272 11296
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 31956 11206 32076 11234
rect 32126 11248 32182 11257
rect 31850 11112 31906 11121
rect 31850 11047 31906 11056
rect 31864 10742 31892 11047
rect 31852 10736 31904 10742
rect 31852 10678 31904 10684
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31668 9920 31720 9926
rect 31668 9862 31720 9868
rect 31666 9752 31722 9761
rect 31772 9738 31800 9998
rect 31722 9710 31800 9738
rect 31666 9687 31722 9696
rect 31772 9382 31800 9710
rect 31852 9580 31904 9586
rect 31956 9568 31984 11206
rect 32126 11183 32182 11192
rect 32140 11150 32168 11183
rect 32128 11144 32180 11150
rect 32048 11104 32128 11132
rect 32048 10674 32076 11104
rect 32128 11086 32180 11092
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32128 11008 32180 11014
rect 32128 10950 32180 10956
rect 32036 10668 32088 10674
rect 32036 10610 32088 10616
rect 32140 10062 32168 10950
rect 32232 10470 32260 11086
rect 32220 10464 32272 10470
rect 32220 10406 32272 10412
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32140 9722 32168 9998
rect 32128 9716 32180 9722
rect 32128 9658 32180 9664
rect 31904 9540 31984 9568
rect 31852 9522 31904 9528
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31772 9178 31800 9318
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 31128 8894 31432 8922
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 31128 8634 31156 8774
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 31036 8090 31064 8434
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 30944 6866 31064 6882
rect 30944 6860 31076 6866
rect 30944 6854 31024 6860
rect 31024 6802 31076 6808
rect 31208 6724 31260 6730
rect 31208 6666 31260 6672
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 31024 6656 31076 6662
rect 31024 6598 31076 6604
rect 30208 6254 30236 6598
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 29472 5914 29500 6190
rect 29552 6112 29604 6118
rect 29552 6054 29604 6060
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29564 5710 29592 6054
rect 29932 5778 29960 6054
rect 29920 5772 29972 5778
rect 29920 5714 29972 5720
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29564 5166 29592 5646
rect 30392 5642 30420 6258
rect 31036 5914 31064 6598
rect 31220 5914 31248 6666
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31220 5710 31248 5850
rect 31404 5794 31432 8894
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31496 8294 31524 8842
rect 31576 8832 31628 8838
rect 31576 8774 31628 8780
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31588 8498 31616 8774
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31484 8288 31536 8294
rect 31484 8230 31536 8236
rect 31496 7886 31524 8230
rect 31588 7886 31616 8434
rect 31680 8362 31708 8774
rect 31772 8498 31800 9114
rect 31864 8974 31892 9522
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 32140 8634 32168 8910
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 31668 6248 31720 6254
rect 31668 6190 31720 6196
rect 31680 5914 31708 6190
rect 32232 6118 32260 6598
rect 32220 6112 32272 6118
rect 32220 6054 32272 6060
rect 31668 5908 31720 5914
rect 31668 5850 31720 5856
rect 31404 5766 31708 5794
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 30380 5636 30432 5642
rect 30380 5578 30432 5584
rect 30392 5522 30420 5578
rect 30300 5494 30420 5522
rect 30300 5302 30328 5494
rect 29736 5296 29788 5302
rect 29736 5238 29788 5244
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 29564 4622 29592 5102
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29368 3188 29420 3194
rect 29368 3130 29420 3136
rect 29748 3126 29776 5238
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 29840 3738 29868 5102
rect 31312 4622 31340 5102
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 31404 4078 31432 5766
rect 31680 5710 31708 5766
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31588 5370 31616 5646
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 32232 4146 32260 6054
rect 32324 5914 32352 15370
rect 34532 15162 34560 16594
rect 34520 15156 34572 15162
rect 34520 15098 34572 15104
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 33140 14340 33192 14346
rect 33140 14282 33192 14288
rect 33152 14006 33180 14282
rect 33140 14000 33192 14006
rect 33140 13942 33192 13948
rect 34440 13938 34468 15030
rect 34532 14482 34560 15098
rect 34520 14476 34572 14482
rect 34520 14418 34572 14424
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34612 13728 34664 13734
rect 34612 13670 34664 13676
rect 34152 13524 34204 13530
rect 34152 13466 34204 13472
rect 34164 13326 34192 13466
rect 34624 13326 34652 13670
rect 32680 13320 32732 13326
rect 32680 13262 32732 13268
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 32692 12850 32720 13262
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32508 12442 32536 12786
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32404 12368 32456 12374
rect 32404 12310 32456 12316
rect 32416 11150 32444 12310
rect 32508 11762 32536 12378
rect 34624 12374 34652 13262
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34716 12986 34744 13126
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34704 12844 34756 12850
rect 34704 12786 34756 12792
rect 34612 12368 34664 12374
rect 34612 12310 34664 12316
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32416 9178 32444 11086
rect 32508 11082 32536 11698
rect 34428 11620 34480 11626
rect 34428 11562 34480 11568
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 34440 10742 34468 11562
rect 34428 10736 34480 10742
rect 34428 10678 34480 10684
rect 33968 9920 34020 9926
rect 33968 9862 34020 9868
rect 34244 9920 34296 9926
rect 34244 9862 34296 9868
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33152 9178 33180 9318
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33600 8288 33652 8294
rect 33600 8230 33652 8236
rect 33612 7002 33640 8230
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33060 5914 33088 6598
rect 33980 6458 34008 9862
rect 34256 9518 34284 9862
rect 34440 9722 34468 10678
rect 34624 10130 34652 12038
rect 34716 11558 34744 12786
rect 34704 11552 34756 11558
rect 34704 11494 34756 11500
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34716 10810 34744 11086
rect 34704 10804 34756 10810
rect 34704 10746 34756 10752
rect 34704 10464 34756 10470
rect 34704 10406 34756 10412
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34428 9716 34480 9722
rect 34428 9658 34480 9664
rect 34716 9654 34744 10406
rect 34704 9648 34756 9654
rect 34704 9590 34756 9596
rect 34244 9512 34296 9518
rect 34244 9454 34296 9460
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34164 8634 34192 8774
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 34256 8362 34284 9454
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 34716 7954 34744 9590
rect 34704 7948 34756 7954
rect 34704 7890 34756 7896
rect 34520 6792 34572 6798
rect 34520 6734 34572 6740
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 33968 6452 34020 6458
rect 33968 6394 34020 6400
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 33152 5914 33180 6054
rect 33888 5914 33916 6394
rect 34532 6322 34560 6734
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 33140 5908 33192 5914
rect 33140 5850 33192 5856
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 34532 4690 34560 6258
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34520 4684 34572 4690
rect 34520 4626 34572 4632
rect 32772 4616 32824 4622
rect 34624 4570 34652 5170
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34716 4826 34744 4966
rect 34704 4820 34756 4826
rect 34704 4762 34756 4768
rect 32772 4558 32824 4564
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 31392 4072 31444 4078
rect 31392 4014 31444 4020
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30472 3596 30524 3602
rect 30472 3538 30524 3544
rect 30484 3194 30512 3538
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 30576 3194 30604 3470
rect 30852 3194 30880 3470
rect 31864 3466 31892 3878
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31852 3460 31904 3466
rect 31852 3402 31904 3408
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 29736 3120 29788 3126
rect 29736 3062 29788 3068
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 17644 2944 18000 2972
rect 29000 2984 29052 2990
rect 17592 2926 17644 2932
rect 29000 2926 29052 2932
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 30838 2952 30894 2961
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 25872 2916 25924 2922
rect 25872 2858 25924 2864
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 18064 2582 18092 2858
rect 25884 2650 25912 2858
rect 26620 2650 26648 2858
rect 29012 2774 29040 2926
rect 29012 2746 29224 2774
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 29196 2514 29224 2746
rect 30300 2650 30328 2926
rect 30838 2887 30840 2896
rect 30892 2887 30894 2896
rect 30840 2858 30892 2864
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 32232 2514 32260 2790
rect 32692 2650 32720 3674
rect 32784 3602 32812 4558
rect 33784 4548 33836 4554
rect 33784 4490 33836 4496
rect 34532 4542 34652 4570
rect 33048 4480 33100 4486
rect 33048 4422 33100 4428
rect 33060 4146 33088 4422
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33244 3602 33272 3878
rect 32772 3596 32824 3602
rect 32772 3538 32824 3544
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 32784 3074 32812 3538
rect 32784 3058 32904 3074
rect 32784 3052 32916 3058
rect 32784 3046 32864 3052
rect 32864 2994 32916 3000
rect 32680 2644 32732 2650
rect 32680 2586 32732 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 29184 2508 29236 2514
rect 29184 2450 29236 2456
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 33244 2446 33272 3538
rect 33796 3126 33824 4490
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 33980 4146 34192 4162
rect 34256 4146 34284 4218
rect 33980 4140 34204 4146
rect 33980 4134 34152 4140
rect 33980 4078 34008 4134
rect 34152 4082 34204 4088
rect 34244 4140 34296 4146
rect 34244 4082 34296 4088
rect 33968 4072 34020 4078
rect 34532 4026 34560 4542
rect 34612 4480 34664 4486
rect 34612 4422 34664 4428
rect 34624 4146 34652 4422
rect 34704 4276 34756 4282
rect 34704 4218 34756 4224
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 33968 4014 34020 4020
rect 34072 4010 34560 4026
rect 34060 4004 34560 4010
rect 34112 3998 34560 4004
rect 34060 3946 34112 3952
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 34428 3936 34480 3942
rect 34428 3878 34480 3884
rect 34520 3936 34572 3942
rect 34520 3878 34572 3884
rect 33980 3670 34008 3878
rect 33968 3664 34020 3670
rect 33968 3606 34020 3612
rect 34164 3398 34192 3878
rect 34440 3466 34468 3878
rect 34532 3738 34560 3878
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 34624 3482 34652 3674
rect 34716 3602 34744 4218
rect 34704 3596 34756 3602
rect 34704 3538 34756 3544
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34532 3454 34652 3482
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 33784 3120 33836 3126
rect 33784 3062 33836 3068
rect 33796 2938 33824 3062
rect 33796 2922 34284 2938
rect 33796 2916 34296 2922
rect 33796 2910 34244 2916
rect 34244 2858 34296 2864
rect 34440 2854 34468 3402
rect 34532 3126 34560 3454
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 3126 34652 3334
rect 34716 3194 34744 3538
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34520 3120 34572 3126
rect 34520 3062 34572 3068
rect 34612 3120 34664 3126
rect 34612 3062 34664 3068
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 8576 2440 8628 2446
rect 17500 2440 17552 2446
rect 8576 2382 8628 2388
rect 17420 2400 17500 2428
rect 32 800 60 2382
rect 8588 1306 8616 2382
rect 8404 1278 8616 1306
rect 8404 800 8432 1278
rect 17420 800 17448 2400
rect 17500 2382 17552 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 26528 1306 26556 2382
rect 26436 1278 26556 1306
rect 26436 800 26464 1278
rect 34808 800 34836 23802
rect 35452 23730 35480 24822
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35636 22982 35664 26998
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 35820 26586 35848 26930
rect 35912 26874 35940 26930
rect 36004 26874 36032 28358
rect 36096 27878 36124 28562
rect 36728 28008 36780 28014
rect 36728 27950 36780 27956
rect 36084 27872 36136 27878
rect 36084 27814 36136 27820
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 36096 27470 36124 27814
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36188 26994 36216 27814
rect 36740 27674 36768 27950
rect 36728 27668 36780 27674
rect 36728 27610 36780 27616
rect 36820 27668 36872 27674
rect 36820 27610 36872 27616
rect 36360 27328 36412 27334
rect 36360 27270 36412 27276
rect 36372 27062 36400 27270
rect 36832 27130 36860 27610
rect 36924 27470 36952 31726
rect 37752 31346 37780 31726
rect 38016 31680 38068 31686
rect 38016 31622 38068 31628
rect 38028 31414 38056 31622
rect 38016 31408 38068 31414
rect 38016 31350 38068 31356
rect 37740 31340 37792 31346
rect 37740 31282 37792 31288
rect 38120 30326 38148 31726
rect 38108 30320 38160 30326
rect 38108 30262 38160 30268
rect 38764 30190 38792 31726
rect 39132 31346 39160 33374
rect 39224 33318 39252 33510
rect 39488 33516 39540 33522
rect 39488 33458 39540 33464
rect 39212 33312 39264 33318
rect 39212 33254 39264 33260
rect 39856 33312 39908 33318
rect 39856 33254 39908 33260
rect 39868 33114 39896 33254
rect 39856 33108 39908 33114
rect 39856 33050 39908 33056
rect 39488 31680 39540 31686
rect 39488 31622 39540 31628
rect 39500 31482 39528 31622
rect 39488 31476 39540 31482
rect 39488 31418 39540 31424
rect 39120 31340 39172 31346
rect 39040 31300 39120 31328
rect 38108 30184 38160 30190
rect 38108 30126 38160 30132
rect 38752 30184 38804 30190
rect 38752 30126 38804 30132
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37096 29504 37148 29510
rect 37096 29446 37148 29452
rect 37280 29504 37332 29510
rect 37280 29446 37332 29452
rect 37108 29306 37136 29446
rect 37096 29300 37148 29306
rect 37096 29242 37148 29248
rect 37292 29102 37320 29446
rect 37476 29238 37504 29990
rect 37464 29232 37516 29238
rect 37464 29174 37516 29180
rect 37280 29096 37332 29102
rect 37280 29038 37332 29044
rect 36912 27464 36964 27470
rect 36912 27406 36964 27412
rect 36820 27124 36872 27130
rect 36820 27066 36872 27072
rect 36360 27056 36412 27062
rect 36360 26998 36412 27004
rect 36176 26988 36228 26994
rect 36176 26930 36228 26936
rect 35912 26846 36216 26874
rect 35808 26580 35860 26586
rect 35808 26522 35860 26528
rect 35808 24132 35860 24138
rect 35808 24074 35860 24080
rect 35820 23866 35848 24074
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35624 22976 35676 22982
rect 35624 22918 35676 22924
rect 35636 22710 35664 22918
rect 35348 22704 35400 22710
rect 35624 22704 35676 22710
rect 35400 22652 35572 22658
rect 35348 22646 35572 22652
rect 35624 22646 35676 22652
rect 35360 22630 35572 22646
rect 35440 22568 35492 22574
rect 35440 22510 35492 22516
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22030 35480 22510
rect 35544 22030 35572 22630
rect 35624 22568 35676 22574
rect 35624 22510 35676 22516
rect 35636 22438 35664 22510
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 36004 22234 36032 22986
rect 36188 22658 36216 26846
rect 36924 26382 36952 27406
rect 37292 26382 37320 29038
rect 38120 26790 38148 30126
rect 39040 29170 39068 31300
rect 39120 31282 39172 31288
rect 39500 30394 39528 31418
rect 39488 30388 39540 30394
rect 39488 30330 39540 30336
rect 39120 30252 39172 30258
rect 39120 30194 39172 30200
rect 39028 29164 39080 29170
rect 39028 29106 39080 29112
rect 38752 29096 38804 29102
rect 38752 29038 38804 29044
rect 38764 28626 38792 29038
rect 39132 28694 39160 30194
rect 39212 30184 39264 30190
rect 39212 30126 39264 30132
rect 39224 29306 39252 30126
rect 39304 30048 39356 30054
rect 39304 29990 39356 29996
rect 39316 29850 39344 29990
rect 39304 29844 39356 29850
rect 39304 29786 39356 29792
rect 39212 29300 39264 29306
rect 39212 29242 39264 29248
rect 39396 29300 39448 29306
rect 39396 29242 39448 29248
rect 39120 28688 39172 28694
rect 39120 28630 39172 28636
rect 38752 28620 38804 28626
rect 38752 28562 38804 28568
rect 39408 28558 39436 29242
rect 39500 29170 39528 30330
rect 39580 30252 39632 30258
rect 39632 30212 39804 30240
rect 39580 30194 39632 30200
rect 39672 30048 39724 30054
rect 39672 29990 39724 29996
rect 39684 29850 39712 29990
rect 39672 29844 39724 29850
rect 39672 29786 39724 29792
rect 39580 29504 39632 29510
rect 39580 29446 39632 29452
rect 39488 29164 39540 29170
rect 39488 29106 39540 29112
rect 38936 28552 38988 28558
rect 38936 28494 38988 28500
rect 39396 28552 39448 28558
rect 39396 28494 39448 28500
rect 38948 28218 38976 28494
rect 38936 28212 38988 28218
rect 38936 28154 38988 28160
rect 38844 28076 38896 28082
rect 38844 28018 38896 28024
rect 39304 28076 39356 28082
rect 39304 28018 39356 28024
rect 39488 28076 39540 28082
rect 39488 28018 39540 28024
rect 38856 27402 38884 28018
rect 39316 27606 39344 28018
rect 39500 27674 39528 28018
rect 39488 27668 39540 27674
rect 39488 27610 39540 27616
rect 39304 27600 39356 27606
rect 39304 27542 39356 27548
rect 38844 27396 38896 27402
rect 38844 27338 38896 27344
rect 38108 26784 38160 26790
rect 38108 26726 38160 26732
rect 36912 26376 36964 26382
rect 36912 26318 36964 26324
rect 37280 26376 37332 26382
rect 37280 26318 37332 26324
rect 36268 25492 36320 25498
rect 36268 25434 36320 25440
rect 36280 23730 36308 25434
rect 36924 25294 36952 26318
rect 37292 25362 37320 26318
rect 37740 26308 37792 26314
rect 37740 26250 37792 26256
rect 37752 26042 37780 26250
rect 38752 26240 38804 26246
rect 38752 26182 38804 26188
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 38384 25832 38436 25838
rect 38384 25774 38436 25780
rect 38396 25498 38424 25774
rect 38660 25696 38712 25702
rect 38660 25638 38712 25644
rect 38672 25498 38700 25638
rect 38384 25492 38436 25498
rect 38384 25434 38436 25440
rect 38660 25492 38712 25498
rect 38660 25434 38712 25440
rect 37280 25356 37332 25362
rect 37280 25298 37332 25304
rect 38476 25356 38528 25362
rect 38476 25298 38528 25304
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 38488 24750 38516 25298
rect 38476 24744 38528 24750
rect 38476 24686 38528 24692
rect 38764 24614 38792 26182
rect 37740 24608 37792 24614
rect 37740 24550 37792 24556
rect 38752 24608 38804 24614
rect 38752 24550 38804 24556
rect 37752 24410 37780 24550
rect 37740 24404 37792 24410
rect 37740 24346 37792 24352
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 37924 24132 37976 24138
rect 37924 24074 37976 24080
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36464 23526 36492 24006
rect 37292 23662 37320 24006
rect 37936 23866 37964 24074
rect 37924 23860 37976 23866
rect 37924 23802 37976 23808
rect 38568 23860 38620 23866
rect 38568 23802 38620 23808
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 37280 23656 37332 23662
rect 37280 23598 37332 23604
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 36360 23112 36412 23118
rect 36360 23054 36412 23060
rect 36372 22778 36400 23054
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36084 22636 36136 22642
rect 36188 22630 36400 22658
rect 36084 22578 36136 22584
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 35360 21690 35388 21966
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 35452 21418 35480 21966
rect 35544 21622 35572 21966
rect 35808 21888 35860 21894
rect 35808 21830 35860 21836
rect 35532 21616 35584 21622
rect 35532 21558 35584 21564
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35532 21480 35584 21486
rect 35532 21422 35584 21428
rect 35440 21412 35492 21418
rect 35440 21354 35492 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35544 20942 35572 21422
rect 35728 21350 35756 21490
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35728 20942 35756 21286
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35440 20868 35492 20874
rect 35440 20810 35492 20816
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35452 19854 35480 20810
rect 35820 20466 35848 21830
rect 36096 21690 36124 22578
rect 36176 22500 36228 22506
rect 36176 22442 36228 22448
rect 36084 21684 36136 21690
rect 36084 21626 36136 21632
rect 36084 21548 36136 21554
rect 36188 21536 36216 22442
rect 36268 22432 36320 22438
rect 36268 22374 36320 22380
rect 36280 22234 36308 22374
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 36136 21508 36216 21536
rect 36084 21490 36136 21496
rect 35808 20460 35860 20466
rect 35808 20402 35860 20408
rect 35624 20052 35676 20058
rect 35624 19994 35676 20000
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 35532 19848 35584 19854
rect 35532 19790 35584 19796
rect 34888 19780 34940 19786
rect 34888 19722 34940 19728
rect 34900 19514 34928 19722
rect 35544 19514 35572 19790
rect 34888 19508 34940 19514
rect 34888 19450 34940 19456
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34888 18760 34940 18766
rect 35256 18760 35308 18766
rect 34940 18708 35256 18714
rect 34888 18702 35308 18708
rect 34900 18686 35296 18702
rect 35360 18426 35388 19314
rect 35544 18902 35572 19450
rect 35636 19378 35664 19994
rect 35820 19990 35848 20402
rect 35808 19984 35860 19990
rect 35808 19926 35860 19932
rect 35900 19916 35952 19922
rect 35900 19858 35952 19864
rect 35716 19712 35768 19718
rect 35716 19654 35768 19660
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35624 19372 35676 19378
rect 35624 19314 35676 19320
rect 35532 18896 35584 18902
rect 35532 18838 35584 18844
rect 35636 18766 35664 19314
rect 35728 18970 35756 19654
rect 35820 19417 35848 19654
rect 35806 19408 35862 19417
rect 35912 19378 35940 19858
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 35806 19343 35862 19352
rect 35900 19372 35952 19378
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 35624 18760 35676 18766
rect 35624 18702 35676 18708
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35820 17610 35848 19343
rect 35900 19314 35952 19320
rect 35912 19174 35940 19314
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35912 18766 35940 19110
rect 36188 18970 36216 19790
rect 36372 19360 36400 22630
rect 36464 21690 36492 23462
rect 36556 23322 36584 23598
rect 36544 23316 36596 23322
rect 36544 23258 36596 23264
rect 36636 23044 36688 23050
rect 36636 22986 36688 22992
rect 36544 22976 36596 22982
rect 36544 22918 36596 22924
rect 36452 21684 36504 21690
rect 36452 21626 36504 21632
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36464 20942 36492 21490
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36464 20466 36492 20878
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36556 19378 36584 22918
rect 36648 19718 36676 22986
rect 36820 20256 36872 20262
rect 36820 20198 36872 20204
rect 36636 19712 36688 19718
rect 36636 19654 36688 19660
rect 36728 19712 36780 19718
rect 36728 19654 36780 19660
rect 36740 19378 36768 19654
rect 36832 19378 36860 20198
rect 37292 19854 37320 23598
rect 38580 23526 38608 23802
rect 38672 23730 38700 24210
rect 38764 24206 38792 24550
rect 38752 24200 38804 24206
rect 38752 24142 38804 24148
rect 38660 23724 38712 23730
rect 38660 23666 38712 23672
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 37740 22568 37792 22574
rect 37740 22510 37792 22516
rect 37752 22234 37780 22510
rect 37740 22228 37792 22234
rect 37740 22170 37792 22176
rect 38200 22092 38252 22098
rect 38200 22034 38252 22040
rect 38108 21956 38160 21962
rect 38108 21898 38160 21904
rect 38120 21690 38148 21898
rect 38108 21684 38160 21690
rect 38108 21626 38160 21632
rect 38212 20466 38240 22034
rect 38580 21962 38608 23462
rect 38672 23322 38700 23666
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38672 22094 38700 23258
rect 38752 22094 38804 22098
rect 38672 22092 38804 22094
rect 38672 22066 38752 22092
rect 38752 22034 38804 22040
rect 38568 21956 38620 21962
rect 38568 21898 38620 21904
rect 38200 20460 38252 20466
rect 38200 20402 38252 20408
rect 38580 20346 38608 21898
rect 38856 21350 38884 27338
rect 39396 26444 39448 26450
rect 39396 26386 39448 26392
rect 39408 26042 39436 26386
rect 39592 26314 39620 29446
rect 39776 28626 39804 30212
rect 39856 29640 39908 29646
rect 39856 29582 39908 29588
rect 39868 29306 39896 29582
rect 39960 29578 39988 33866
rect 40224 33516 40276 33522
rect 40224 33458 40276 33464
rect 40236 33114 40264 33458
rect 40224 33108 40276 33114
rect 40224 33050 40276 33056
rect 40132 32428 40184 32434
rect 40132 32370 40184 32376
rect 40144 32026 40172 32370
rect 40132 32020 40184 32026
rect 40132 31962 40184 31968
rect 40236 30734 40264 33050
rect 40420 32842 40448 33934
rect 40500 33448 40552 33454
rect 40500 33390 40552 33396
rect 40408 32836 40460 32842
rect 40408 32778 40460 32784
rect 40420 32366 40448 32778
rect 40408 32360 40460 32366
rect 40408 32302 40460 32308
rect 40512 31890 40540 33390
rect 40604 32842 40632 34614
rect 41616 34610 41644 35686
rect 41708 34746 41736 35866
rect 41892 35866 42012 35894
rect 41696 34740 41748 34746
rect 41696 34682 41748 34688
rect 41604 34604 41656 34610
rect 41604 34546 41656 34552
rect 40684 34400 40736 34406
rect 40684 34342 40736 34348
rect 40776 34400 40828 34406
rect 40776 34342 40828 34348
rect 40696 33658 40724 34342
rect 40788 34066 40816 34342
rect 40776 34060 40828 34066
rect 40776 34002 40828 34008
rect 41328 34060 41380 34066
rect 41328 34002 41380 34008
rect 40684 33652 40736 33658
rect 40684 33594 40736 33600
rect 41340 33522 41368 34002
rect 41328 33516 41380 33522
rect 41328 33458 41380 33464
rect 41512 33312 41564 33318
rect 41512 33254 41564 33260
rect 40684 32972 40736 32978
rect 40684 32914 40736 32920
rect 40592 32836 40644 32842
rect 40592 32778 40644 32784
rect 40696 32230 40724 32914
rect 41144 32768 41196 32774
rect 41144 32710 41196 32716
rect 41156 32502 41184 32710
rect 41144 32496 41196 32502
rect 41144 32438 41196 32444
rect 40684 32224 40736 32230
rect 40684 32166 40736 32172
rect 41236 32224 41288 32230
rect 41236 32166 41288 32172
rect 40500 31884 40552 31890
rect 40500 31826 40552 31832
rect 41248 31822 41276 32166
rect 41524 31890 41552 33254
rect 41512 31884 41564 31890
rect 41512 31826 41564 31832
rect 41236 31816 41288 31822
rect 41236 31758 41288 31764
rect 40316 30796 40368 30802
rect 40316 30738 40368 30744
rect 40224 30728 40276 30734
rect 40224 30670 40276 30676
rect 40132 30252 40184 30258
rect 40132 30194 40184 30200
rect 40040 30184 40092 30190
rect 40040 30126 40092 30132
rect 39948 29572 40000 29578
rect 39948 29514 40000 29520
rect 39856 29300 39908 29306
rect 39856 29242 39908 29248
rect 39948 29232 40000 29238
rect 40052 29186 40080 30126
rect 40144 29850 40172 30194
rect 40132 29844 40184 29850
rect 40132 29786 40184 29792
rect 40144 29306 40172 29786
rect 40236 29714 40264 30670
rect 40328 30394 40356 30738
rect 40592 30592 40644 30598
rect 40592 30534 40644 30540
rect 40316 30388 40368 30394
rect 40316 30330 40368 30336
rect 40500 30048 40552 30054
rect 40500 29990 40552 29996
rect 40224 29708 40276 29714
rect 40224 29650 40276 29656
rect 40236 29306 40264 29650
rect 40512 29646 40540 29990
rect 40500 29640 40552 29646
rect 40500 29582 40552 29588
rect 40132 29300 40184 29306
rect 40132 29242 40184 29248
rect 40224 29300 40276 29306
rect 40224 29242 40276 29248
rect 40000 29180 40080 29186
rect 39948 29174 40080 29180
rect 39960 29158 40080 29174
rect 40408 29164 40460 29170
rect 39960 29102 39988 29158
rect 40408 29106 40460 29112
rect 39948 29096 40000 29102
rect 39948 29038 40000 29044
rect 40040 29028 40092 29034
rect 40040 28970 40092 28976
rect 39764 28620 39816 28626
rect 39764 28562 39816 28568
rect 39776 28218 39804 28562
rect 40052 28558 40080 28970
rect 40420 28694 40448 29106
rect 40408 28688 40460 28694
rect 40408 28630 40460 28636
rect 40604 28558 40632 30534
rect 41248 30326 41276 31758
rect 41236 30320 41288 30326
rect 41236 30262 41288 30268
rect 41248 29850 41276 30262
rect 41512 30252 41564 30258
rect 41512 30194 41564 30200
rect 41328 30116 41380 30122
rect 41328 30058 41380 30064
rect 41340 29850 41368 30058
rect 41420 30048 41472 30054
rect 41420 29990 41472 29996
rect 41236 29844 41288 29850
rect 41236 29786 41288 29792
rect 41328 29844 41380 29850
rect 41328 29786 41380 29792
rect 41340 29646 41368 29786
rect 41432 29714 41460 29990
rect 41524 29714 41552 30194
rect 41420 29708 41472 29714
rect 41420 29650 41472 29656
rect 41512 29708 41564 29714
rect 41512 29650 41564 29656
rect 40776 29640 40828 29646
rect 40776 29582 40828 29588
rect 41328 29640 41380 29646
rect 41328 29582 41380 29588
rect 40788 29306 40816 29582
rect 40960 29504 41012 29510
rect 40960 29446 41012 29452
rect 41696 29504 41748 29510
rect 41696 29446 41748 29452
rect 41788 29504 41840 29510
rect 41788 29446 41840 29452
rect 40776 29300 40828 29306
rect 40776 29242 40828 29248
rect 40868 29164 40920 29170
rect 40868 29106 40920 29112
rect 40880 29034 40908 29106
rect 40868 29028 40920 29034
rect 40868 28970 40920 28976
rect 40880 28558 40908 28970
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 40316 28552 40368 28558
rect 40316 28494 40368 28500
rect 40592 28552 40644 28558
rect 40592 28494 40644 28500
rect 40868 28552 40920 28558
rect 40868 28494 40920 28500
rect 39948 28484 40000 28490
rect 39948 28426 40000 28432
rect 39764 28212 39816 28218
rect 39764 28154 39816 28160
rect 39764 27600 39816 27606
rect 39764 27542 39816 27548
rect 39776 27402 39804 27542
rect 39764 27396 39816 27402
rect 39764 27338 39816 27344
rect 39488 26308 39540 26314
rect 39488 26250 39540 26256
rect 39580 26308 39632 26314
rect 39580 26250 39632 26256
rect 39396 26036 39448 26042
rect 39396 25978 39448 25984
rect 39500 25906 39528 26250
rect 39592 26042 39620 26250
rect 39580 26036 39632 26042
rect 39580 25978 39632 25984
rect 39488 25900 39540 25906
rect 39488 25842 39540 25848
rect 39028 25696 39080 25702
rect 39028 25638 39080 25644
rect 38844 21344 38896 21350
rect 38844 21286 38896 21292
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 38764 20602 38792 20742
rect 38752 20596 38804 20602
rect 38752 20538 38804 20544
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38856 20346 38884 20538
rect 38580 20318 38884 20346
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 36912 19712 36964 19718
rect 36912 19654 36964 19660
rect 36924 19378 36952 19654
rect 36452 19372 36504 19378
rect 36372 19332 36452 19360
rect 36268 19236 36320 19242
rect 36268 19178 36320 19184
rect 36176 18964 36228 18970
rect 36176 18906 36228 18912
rect 35900 18760 35952 18766
rect 35900 18702 35952 18708
rect 36188 18426 36216 18906
rect 36280 18766 36308 19178
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36372 18222 36400 19332
rect 36452 19314 36504 19320
rect 36544 19372 36596 19378
rect 36544 19314 36596 19320
rect 36728 19372 36780 19378
rect 36728 19314 36780 19320
rect 36820 19372 36872 19378
rect 36820 19314 36872 19320
rect 36912 19372 36964 19378
rect 36912 19314 36964 19320
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 36556 18970 36584 19314
rect 36832 19258 36860 19314
rect 37384 19258 37412 19314
rect 36832 19230 37412 19258
rect 37280 19168 37332 19174
rect 37280 19110 37332 19116
rect 36544 18964 36596 18970
rect 36544 18906 36596 18912
rect 37292 18698 37320 19110
rect 37464 18828 37516 18834
rect 37464 18770 37516 18776
rect 37280 18692 37332 18698
rect 37280 18634 37332 18640
rect 37476 18222 37504 18770
rect 38580 18698 38608 20318
rect 38948 20058 38976 20878
rect 38936 20052 38988 20058
rect 38936 19994 38988 20000
rect 38568 18692 38620 18698
rect 38568 18634 38620 18640
rect 38200 18624 38252 18630
rect 38200 18566 38252 18572
rect 38212 18426 38240 18566
rect 38200 18420 38252 18426
rect 38200 18362 38252 18368
rect 36360 18216 36412 18222
rect 36360 18158 36412 18164
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 35808 17604 35860 17610
rect 35808 17546 35860 17552
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35452 16454 35480 17070
rect 35440 16448 35492 16454
rect 35440 16390 35492 16396
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35452 15434 35480 16390
rect 35820 15910 35848 17546
rect 37476 17542 37504 18158
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35912 16250 35940 16934
rect 35992 16788 36044 16794
rect 35992 16730 36044 16736
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 36004 16250 36032 16730
rect 36820 16516 36872 16522
rect 36820 16458 36872 16464
rect 36728 16448 36780 16454
rect 36728 16390 36780 16396
rect 36740 16250 36768 16390
rect 35900 16244 35952 16250
rect 35900 16186 35952 16192
rect 35992 16244 36044 16250
rect 35992 16186 36044 16192
rect 36728 16244 36780 16250
rect 36728 16186 36780 16192
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 36832 15434 36860 16458
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 35440 15428 35492 15434
rect 35440 15370 35492 15376
rect 36820 15428 36872 15434
rect 36820 15370 36872 15376
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35360 15094 35388 15302
rect 35348 15088 35400 15094
rect 35348 15030 35400 15036
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14482 35388 14758
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35452 13190 35480 15370
rect 35900 15360 35952 15366
rect 35900 15302 35952 15308
rect 35912 15162 35940 15302
rect 35900 15156 35952 15162
rect 35900 15098 35952 15104
rect 35716 14952 35768 14958
rect 35716 14894 35768 14900
rect 35728 14618 35756 14894
rect 36360 14816 36412 14822
rect 36360 14758 36412 14764
rect 35716 14612 35768 14618
rect 35716 14554 35768 14560
rect 35992 14408 36044 14414
rect 35992 14350 36044 14356
rect 36004 14006 36032 14350
rect 36372 14006 36400 14758
rect 36832 14414 36860 15370
rect 36820 14408 36872 14414
rect 36820 14350 36872 14356
rect 36832 14006 36860 14350
rect 37200 14056 37228 15846
rect 37292 15162 37320 16730
rect 37476 16658 37504 17478
rect 37844 17338 37872 18158
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 38028 16250 38056 17138
rect 38212 16590 38240 18362
rect 38200 16584 38252 16590
rect 38200 16526 38252 16532
rect 38384 16448 38436 16454
rect 38384 16390 38436 16396
rect 38016 16244 38068 16250
rect 38016 16186 38068 16192
rect 37464 16176 37516 16182
rect 37464 16118 37516 16124
rect 37476 15706 37504 16118
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 37280 15156 37332 15162
rect 37280 15098 37332 15104
rect 37280 14068 37332 14074
rect 37200 14028 37280 14056
rect 37280 14010 37332 14016
rect 35992 14000 36044 14006
rect 35992 13942 36044 13948
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36004 13870 36032 13942
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 35624 13320 35676 13326
rect 35624 13262 35676 13268
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 36728 13320 36780 13326
rect 36728 13262 36780 13268
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 34888 13184 34940 13190
rect 34888 13126 34940 13132
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 34900 12850 34928 13126
rect 35636 12986 35664 13262
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 34888 12844 34940 12850
rect 34888 12786 34940 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 11830 35388 12922
rect 36096 12442 36124 13262
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 35348 11824 35400 11830
rect 35348 11766 35400 11772
rect 36740 11558 36768 13262
rect 37108 12986 37136 13262
rect 37096 12980 37148 12986
rect 37096 12922 37148 12928
rect 37004 12164 37056 12170
rect 37004 12106 37056 12112
rect 37016 11626 37044 12106
rect 37004 11620 37056 11626
rect 37004 11562 37056 11568
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 36452 11552 36504 11558
rect 36452 11494 36504 11500
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10266 35388 10406
rect 35348 10260 35400 10266
rect 35348 10202 35400 10208
rect 35452 10198 35480 10950
rect 35440 10192 35492 10198
rect 35440 10134 35492 10140
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34980 7812 35032 7818
rect 34980 7754 35032 7760
rect 34992 7546 35020 7754
rect 34980 7540 35032 7546
rect 34980 7482 35032 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35348 5364 35400 5370
rect 35348 5306 35400 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4690 35388 5306
rect 35440 5228 35492 5234
rect 35440 5170 35492 5176
rect 35348 4684 35400 4690
rect 35348 4626 35400 4632
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35360 3058 35388 4626
rect 35452 4282 35480 5170
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 35532 3936 35584 3942
rect 35532 3878 35584 3884
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35452 3194 35480 3538
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 35544 3126 35572 3878
rect 35636 3738 35664 11494
rect 36360 11144 36412 11150
rect 36360 11086 36412 11092
rect 36372 10266 36400 11086
rect 36464 10742 36492 11494
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36648 10810 36676 11018
rect 37016 11014 37044 11562
rect 37188 11212 37240 11218
rect 37188 11154 37240 11160
rect 37004 11008 37056 11014
rect 37004 10950 37056 10956
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36452 10736 36504 10742
rect 36452 10678 36504 10684
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 36832 8838 36860 9522
rect 36924 8906 36952 9522
rect 36912 8900 36964 8906
rect 36912 8842 36964 8848
rect 36820 8832 36872 8838
rect 36820 8774 36872 8780
rect 36360 8288 36412 8294
rect 36360 8230 36412 8236
rect 36372 7818 36400 8230
rect 36636 8016 36688 8022
rect 36636 7958 36688 7964
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36372 6730 36400 7754
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36360 6724 36412 6730
rect 36360 6666 36412 6672
rect 36556 6118 36584 7686
rect 36648 7546 36676 7958
rect 36924 7886 36952 8842
rect 37016 8566 37044 10950
rect 37200 9586 37228 11154
rect 37292 9994 37320 14010
rect 37752 13938 37780 15438
rect 37844 14958 37872 16050
rect 38396 15910 38424 16390
rect 38580 15910 38608 18634
rect 37924 15904 37976 15910
rect 37924 15846 37976 15852
rect 38384 15904 38436 15910
rect 38384 15846 38436 15852
rect 38568 15904 38620 15910
rect 38568 15846 38620 15852
rect 37936 15706 37964 15846
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 37832 14952 37884 14958
rect 37832 14894 37884 14900
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37464 13320 37516 13326
rect 37464 13262 37516 13268
rect 37476 12306 37504 13262
rect 37752 12434 37780 13874
rect 37844 13530 37872 14894
rect 38672 14414 38700 15370
rect 39040 15366 39068 25638
rect 39500 24954 39528 25842
rect 39488 24948 39540 24954
rect 39488 24890 39540 24896
rect 39120 24812 39172 24818
rect 39120 24754 39172 24760
rect 39132 24410 39160 24754
rect 39396 24744 39448 24750
rect 39396 24686 39448 24692
rect 39120 24404 39172 24410
rect 39120 24346 39172 24352
rect 39408 24206 39436 24686
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39212 24064 39264 24070
rect 39212 24006 39264 24012
rect 39224 23866 39252 24006
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39776 22098 39804 27338
rect 39960 26382 39988 28426
rect 40328 28082 40356 28494
rect 40316 28076 40368 28082
rect 40316 28018 40368 28024
rect 40328 27470 40356 28018
rect 40316 27464 40368 27470
rect 40316 27406 40368 27412
rect 40972 26450 41000 29446
rect 41512 29232 41564 29238
rect 41512 29174 41564 29180
rect 41328 29164 41380 29170
rect 41328 29106 41380 29112
rect 41236 29096 41288 29102
rect 41236 29038 41288 29044
rect 41248 28966 41276 29038
rect 41236 28960 41288 28966
rect 41236 28902 41288 28908
rect 41340 28082 41368 29106
rect 41328 28076 41380 28082
rect 41328 28018 41380 28024
rect 40500 26444 40552 26450
rect 40500 26386 40552 26392
rect 40960 26444 41012 26450
rect 40960 26386 41012 26392
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 40224 26376 40276 26382
rect 40224 26318 40276 26324
rect 39960 26042 39988 26318
rect 40236 26042 40264 26318
rect 39948 26036 40000 26042
rect 39948 25978 40000 25984
rect 40224 26036 40276 26042
rect 40224 25978 40276 25984
rect 40512 25906 40540 26386
rect 41524 26382 41552 29174
rect 41708 28558 41736 29446
rect 41800 29306 41828 29446
rect 41788 29300 41840 29306
rect 41788 29242 41840 29248
rect 41800 29209 41828 29242
rect 41786 29200 41842 29209
rect 41786 29135 41842 29144
rect 41696 28552 41748 28558
rect 41696 28494 41748 28500
rect 40868 26376 40920 26382
rect 40868 26318 40920 26324
rect 41420 26376 41472 26382
rect 41420 26318 41472 26324
rect 41512 26376 41564 26382
rect 41512 26318 41564 26324
rect 40592 26308 40644 26314
rect 40592 26250 40644 26256
rect 40500 25900 40552 25906
rect 40500 25842 40552 25848
rect 40408 25832 40460 25838
rect 40408 25774 40460 25780
rect 40040 24812 40092 24818
rect 40040 24754 40092 24760
rect 40052 24070 40080 24754
rect 40132 24608 40184 24614
rect 40132 24550 40184 24556
rect 40144 24206 40172 24550
rect 40420 24206 40448 25774
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 40052 23594 40080 24006
rect 40420 23866 40448 24142
rect 40408 23860 40460 23866
rect 40408 23802 40460 23808
rect 40040 23588 40092 23594
rect 40040 23530 40092 23536
rect 40052 22574 40080 23530
rect 40500 23044 40552 23050
rect 40500 22986 40552 22992
rect 40512 22778 40540 22986
rect 40500 22772 40552 22778
rect 40500 22714 40552 22720
rect 40040 22568 40092 22574
rect 40040 22510 40092 22516
rect 39764 22092 39816 22098
rect 39764 22034 39816 22040
rect 39856 21888 39908 21894
rect 39856 21830 39908 21836
rect 39868 21690 39896 21830
rect 39856 21684 39908 21690
rect 39856 21626 39908 21632
rect 39396 21480 39448 21486
rect 39396 21422 39448 21428
rect 39408 21146 39436 21422
rect 39488 21344 39540 21350
rect 39488 21286 39540 21292
rect 39396 21140 39448 21146
rect 39396 21082 39448 21088
rect 39500 21010 39528 21286
rect 39488 21004 39540 21010
rect 39488 20946 39540 20952
rect 39304 20800 39356 20806
rect 39304 20742 39356 20748
rect 39316 19786 39344 20742
rect 39500 20602 39528 20946
rect 39488 20596 39540 20602
rect 39488 20538 39540 20544
rect 39500 19854 39528 20538
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 39304 19780 39356 19786
rect 39304 19722 39356 19728
rect 39316 18426 39344 19722
rect 39304 18420 39356 18426
rect 39304 18362 39356 18368
rect 40604 17338 40632 26250
rect 40880 25974 40908 26318
rect 41144 26240 41196 26246
rect 41144 26182 41196 26188
rect 41156 25974 41184 26182
rect 41432 26042 41460 26318
rect 41420 26036 41472 26042
rect 41420 25978 41472 25984
rect 41524 25974 41552 26318
rect 41788 26308 41840 26314
rect 41788 26250 41840 26256
rect 40868 25968 40920 25974
rect 40868 25910 40920 25916
rect 41144 25968 41196 25974
rect 41144 25910 41196 25916
rect 41512 25968 41564 25974
rect 41512 25910 41564 25916
rect 40684 24812 40736 24818
rect 40684 24754 40736 24760
rect 40776 24812 40828 24818
rect 40776 24754 40828 24760
rect 40696 23866 40724 24754
rect 40788 24342 40816 24754
rect 41604 24744 41656 24750
rect 41604 24686 41656 24692
rect 40776 24336 40828 24342
rect 40776 24278 40828 24284
rect 41420 24268 41472 24274
rect 41420 24210 41472 24216
rect 40684 23860 40736 23866
rect 40684 23802 40736 23808
rect 41432 23730 41460 24210
rect 41616 23866 41644 24686
rect 41696 24608 41748 24614
rect 41696 24550 41748 24556
rect 41708 23866 41736 24550
rect 41800 24410 41828 26250
rect 41788 24404 41840 24410
rect 41788 24346 41840 24352
rect 41604 23860 41656 23866
rect 41604 23802 41656 23808
rect 41696 23860 41748 23866
rect 41696 23802 41748 23808
rect 41420 23724 41472 23730
rect 41420 23666 41472 23672
rect 41800 23662 41828 24346
rect 41788 23656 41840 23662
rect 41788 23598 41840 23604
rect 41604 23520 41656 23526
rect 41604 23462 41656 23468
rect 41616 23118 41644 23462
rect 41800 23322 41828 23598
rect 41788 23316 41840 23322
rect 41788 23258 41840 23264
rect 41604 23112 41656 23118
rect 41604 23054 41656 23060
rect 41800 22642 41828 23258
rect 41788 22636 41840 22642
rect 41788 22578 41840 22584
rect 39120 17332 39172 17338
rect 39120 17274 39172 17280
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 39132 15570 39160 17274
rect 41892 16182 41920 35866
rect 41972 34944 42024 34950
rect 41972 34886 42024 34892
rect 41984 34610 42012 34886
rect 41972 34604 42024 34610
rect 41972 34546 42024 34552
rect 41984 33930 42012 34546
rect 41972 33924 42024 33930
rect 41972 33866 42024 33872
rect 42076 33522 42104 35974
rect 42812 35894 42840 36790
rect 42812 35866 42932 35894
rect 42524 34604 42576 34610
rect 42524 34546 42576 34552
rect 42536 34202 42564 34546
rect 42800 34536 42852 34542
rect 42800 34478 42852 34484
rect 42812 34202 42840 34478
rect 42524 34196 42576 34202
rect 42524 34138 42576 34144
rect 42800 34196 42852 34202
rect 42800 34138 42852 34144
rect 42904 33658 42932 35866
rect 43076 34536 43128 34542
rect 43076 34478 43128 34484
rect 43088 33930 43116 34478
rect 42984 33924 43036 33930
rect 42984 33866 43036 33872
rect 43076 33924 43128 33930
rect 43076 33866 43128 33872
rect 42996 33658 43024 33866
rect 42892 33652 42944 33658
rect 42892 33594 42944 33600
rect 42984 33652 43036 33658
rect 42984 33594 43036 33600
rect 42064 33516 42116 33522
rect 42064 33458 42116 33464
rect 42892 33448 42944 33454
rect 42892 33390 42944 33396
rect 42524 31816 42576 31822
rect 42524 31758 42576 31764
rect 42800 31816 42852 31822
rect 42800 31758 42852 31764
rect 42536 31482 42564 31758
rect 42524 31476 42576 31482
rect 42524 31418 42576 31424
rect 42156 30796 42208 30802
rect 42156 30738 42208 30744
rect 41972 30048 42024 30054
rect 41972 29990 42024 29996
rect 41984 29782 42012 29990
rect 41972 29776 42024 29782
rect 41972 29718 42024 29724
rect 41972 29504 42024 29510
rect 41972 29446 42024 29452
rect 41984 29170 42012 29446
rect 42168 29170 42196 30738
rect 42708 29640 42760 29646
rect 42708 29582 42760 29588
rect 42720 29238 42748 29582
rect 42708 29232 42760 29238
rect 42708 29174 42760 29180
rect 41972 29164 42024 29170
rect 41972 29106 42024 29112
rect 42156 29164 42208 29170
rect 42156 29106 42208 29112
rect 42248 29164 42300 29170
rect 42300 29124 42380 29152
rect 42248 29106 42300 29112
rect 42352 28994 42380 29124
rect 42260 28966 42380 28994
rect 42616 29028 42668 29034
rect 42616 28970 42668 28976
rect 42260 28626 42288 28966
rect 42248 28620 42300 28626
rect 42248 28562 42300 28568
rect 42432 26988 42484 26994
rect 42432 26930 42484 26936
rect 42444 26042 42472 26930
rect 42628 26586 42656 28970
rect 42812 28762 42840 31758
rect 42904 31278 42932 33390
rect 42892 31272 42944 31278
rect 42892 31214 42944 31220
rect 43088 31210 43116 33866
rect 43168 33584 43220 33590
rect 43168 33526 43220 33532
rect 43076 31204 43128 31210
rect 43076 31146 43128 31152
rect 43088 30122 43116 31146
rect 43180 30734 43208 33526
rect 43272 31482 43300 37810
rect 44180 37800 44232 37806
rect 44180 37742 44232 37748
rect 43720 37120 43772 37126
rect 43720 37062 43772 37068
rect 43732 36854 43760 37062
rect 44192 36922 44220 37742
rect 44180 36916 44232 36922
rect 44180 36858 44232 36864
rect 43720 36848 43772 36854
rect 43720 36790 43772 36796
rect 43732 36378 43760 36790
rect 43720 36372 43772 36378
rect 43720 36314 43772 36320
rect 44376 35894 44404 44270
rect 45282 44231 45338 44240
rect 44456 37800 44508 37806
rect 44456 37742 44508 37748
rect 44468 37466 44496 37742
rect 44456 37460 44508 37466
rect 44456 37402 44508 37408
rect 44284 35866 44404 35894
rect 44088 34944 44140 34950
rect 44088 34886 44140 34892
rect 43536 34672 43588 34678
rect 43536 34614 43588 34620
rect 43548 34406 43576 34614
rect 43536 34400 43588 34406
rect 43536 34342 43588 34348
rect 43444 33924 43496 33930
rect 43444 33866 43496 33872
rect 43456 32774 43484 33866
rect 43628 33856 43680 33862
rect 43628 33798 43680 33804
rect 43640 33658 43668 33798
rect 43628 33652 43680 33658
rect 43628 33594 43680 33600
rect 44100 33386 44128 34886
rect 44284 33454 44312 35866
rect 45284 34944 45336 34950
rect 45284 34886 45336 34892
rect 45296 34785 45324 34886
rect 45282 34776 45338 34785
rect 45282 34711 45338 34720
rect 44272 33448 44324 33454
rect 44272 33390 44324 33396
rect 44088 33380 44140 33386
rect 44088 33322 44140 33328
rect 43904 33312 43956 33318
rect 43904 33254 43956 33260
rect 43444 32768 43496 32774
rect 43444 32710 43496 32716
rect 43456 31770 43484 32710
rect 43916 32570 43944 33254
rect 43904 32564 43956 32570
rect 43904 32506 43956 32512
rect 43812 32224 43864 32230
rect 43812 32166 43864 32172
rect 43456 31754 43576 31770
rect 43824 31754 43852 32166
rect 43456 31748 43588 31754
rect 43456 31742 43536 31748
rect 43536 31690 43588 31696
rect 43640 31726 43852 31754
rect 43548 31659 43576 31690
rect 43260 31476 43312 31482
rect 43260 31418 43312 31424
rect 43352 31408 43404 31414
rect 43352 31350 43404 31356
rect 43364 30870 43392 31350
rect 43536 31272 43588 31278
rect 43536 31214 43588 31220
rect 43444 31136 43496 31142
rect 43444 31078 43496 31084
rect 43456 30938 43484 31078
rect 43444 30932 43496 30938
rect 43444 30874 43496 30880
rect 43352 30864 43404 30870
rect 43352 30806 43404 30812
rect 43168 30728 43220 30734
rect 43168 30670 43220 30676
rect 43180 30258 43208 30670
rect 43364 30258 43392 30806
rect 43548 30326 43576 31214
rect 43536 30320 43588 30326
rect 43536 30262 43588 30268
rect 43168 30252 43220 30258
rect 43168 30194 43220 30200
rect 43352 30252 43404 30258
rect 43352 30194 43404 30200
rect 43076 30116 43128 30122
rect 43076 30058 43128 30064
rect 43088 29850 43116 30058
rect 42984 29844 43036 29850
rect 42984 29786 43036 29792
rect 43076 29844 43128 29850
rect 43076 29786 43128 29792
rect 42892 29572 42944 29578
rect 42892 29514 42944 29520
rect 42904 29170 42932 29514
rect 42996 29306 43024 29786
rect 42984 29300 43036 29306
rect 42984 29242 43036 29248
rect 43180 29170 43208 30194
rect 43364 29578 43392 30194
rect 43548 29866 43576 30262
rect 43456 29838 43576 29866
rect 43456 29646 43484 29838
rect 43536 29776 43588 29782
rect 43536 29718 43588 29724
rect 43444 29640 43496 29646
rect 43444 29582 43496 29588
rect 43352 29572 43404 29578
rect 43352 29514 43404 29520
rect 43364 29306 43392 29514
rect 43260 29300 43312 29306
rect 43260 29242 43312 29248
rect 43352 29300 43404 29306
rect 43352 29242 43404 29248
rect 42892 29164 42944 29170
rect 42892 29106 42944 29112
rect 43168 29164 43220 29170
rect 43168 29106 43220 29112
rect 42800 28756 42852 28762
rect 42800 28698 42852 28704
rect 42812 27538 42840 28698
rect 42904 28506 42932 29106
rect 43272 28642 43300 29242
rect 43444 29096 43496 29102
rect 43444 29038 43496 29044
rect 43272 28614 43392 28642
rect 43456 28626 43484 29038
rect 42904 28478 43024 28506
rect 42892 28416 42944 28422
rect 42892 28358 42944 28364
rect 42904 28218 42932 28358
rect 42996 28218 43024 28478
rect 43260 28484 43312 28490
rect 43260 28426 43312 28432
rect 42892 28212 42944 28218
rect 42892 28154 42944 28160
rect 42984 28212 43036 28218
rect 42984 28154 43036 28160
rect 42984 28076 43036 28082
rect 42984 28018 43036 28024
rect 42996 27962 43024 28018
rect 43272 28014 43300 28426
rect 43364 28218 43392 28614
rect 43444 28620 43496 28626
rect 43444 28562 43496 28568
rect 43352 28212 43404 28218
rect 43352 28154 43404 28160
rect 43260 28008 43312 28014
rect 42996 27934 43116 27962
rect 43260 27950 43312 27956
rect 43456 27946 43484 28562
rect 43548 28558 43576 29718
rect 43536 28552 43588 28558
rect 43536 28494 43588 28500
rect 42984 27872 43036 27878
rect 42984 27814 43036 27820
rect 42800 27532 42852 27538
rect 42800 27474 42852 27480
rect 42708 26988 42760 26994
rect 42708 26930 42760 26936
rect 42616 26580 42668 26586
rect 42616 26522 42668 26528
rect 42524 26308 42576 26314
rect 42524 26250 42576 26256
rect 42432 26036 42484 26042
rect 42432 25978 42484 25984
rect 42064 25832 42116 25838
rect 42064 25774 42116 25780
rect 42076 25430 42104 25774
rect 42536 25770 42564 26250
rect 42720 26246 42748 26930
rect 42812 26450 42840 27474
rect 42996 26994 43024 27814
rect 43088 27674 43116 27934
rect 43168 27940 43220 27946
rect 43168 27882 43220 27888
rect 43444 27940 43496 27946
rect 43444 27882 43496 27888
rect 43076 27668 43128 27674
rect 43076 27610 43128 27616
rect 43180 27130 43208 27882
rect 43456 27674 43484 27882
rect 43444 27668 43496 27674
rect 43444 27610 43496 27616
rect 43168 27124 43220 27130
rect 43168 27066 43220 27072
rect 42984 26988 43036 26994
rect 42984 26930 43036 26936
rect 42892 26784 42944 26790
rect 42892 26726 42944 26732
rect 42800 26444 42852 26450
rect 42800 26386 42852 26392
rect 42904 26382 42932 26726
rect 42996 26586 43024 26930
rect 43076 26784 43128 26790
rect 43076 26726 43128 26732
rect 42984 26580 43036 26586
rect 42984 26522 43036 26528
rect 42892 26376 42944 26382
rect 42892 26318 42944 26324
rect 42708 26240 42760 26246
rect 42708 26182 42760 26188
rect 42524 25764 42576 25770
rect 42524 25706 42576 25712
rect 42064 25424 42116 25430
rect 42064 25366 42116 25372
rect 42340 25152 42392 25158
rect 42340 25094 42392 25100
rect 42352 24818 42380 25094
rect 42720 24886 42748 26182
rect 43088 25906 43116 26726
rect 43180 26042 43208 27066
rect 43536 26920 43588 26926
rect 43536 26862 43588 26868
rect 43260 26308 43312 26314
rect 43260 26250 43312 26256
rect 43272 26042 43300 26250
rect 43352 26240 43404 26246
rect 43352 26182 43404 26188
rect 43168 26036 43220 26042
rect 43168 25978 43220 25984
rect 43260 26036 43312 26042
rect 43260 25978 43312 25984
rect 42984 25900 43036 25906
rect 42984 25842 43036 25848
rect 43076 25900 43128 25906
rect 43076 25842 43128 25848
rect 42892 25764 42944 25770
rect 42892 25706 42944 25712
rect 42800 25696 42852 25702
rect 42800 25638 42852 25644
rect 42812 25294 42840 25638
rect 42904 25294 42932 25706
rect 42800 25288 42852 25294
rect 42800 25230 42852 25236
rect 42892 25288 42944 25294
rect 42892 25230 42944 25236
rect 42800 25152 42852 25158
rect 42800 25094 42852 25100
rect 42812 24886 42840 25094
rect 42708 24880 42760 24886
rect 42708 24822 42760 24828
rect 42800 24880 42852 24886
rect 42800 24822 42852 24828
rect 42340 24812 42392 24818
rect 42340 24754 42392 24760
rect 42720 24410 42748 24822
rect 42708 24404 42760 24410
rect 42708 24346 42760 24352
rect 42616 24132 42668 24138
rect 42616 24074 42668 24080
rect 42064 24064 42116 24070
rect 42064 24006 42116 24012
rect 42076 23866 42104 24006
rect 42064 23860 42116 23866
rect 42064 23802 42116 23808
rect 42628 23798 42656 24074
rect 42812 23866 42840 24822
rect 42904 24274 42932 25230
rect 42996 25226 43024 25842
rect 43364 25838 43392 26182
rect 43352 25832 43404 25838
rect 43352 25774 43404 25780
rect 43168 25764 43220 25770
rect 43168 25706 43220 25712
rect 42984 25220 43036 25226
rect 42984 25162 43036 25168
rect 43076 24812 43128 24818
rect 43076 24754 43128 24760
rect 42892 24268 42944 24274
rect 42892 24210 42944 24216
rect 42800 23860 42852 23866
rect 42800 23802 42852 23808
rect 42616 23792 42668 23798
rect 42616 23734 42668 23740
rect 43088 22982 43116 24754
rect 43180 24614 43208 25706
rect 43548 25498 43576 26862
rect 43536 25492 43588 25498
rect 43536 25434 43588 25440
rect 43260 25220 43312 25226
rect 43260 25162 43312 25168
rect 43272 24954 43300 25162
rect 43260 24948 43312 24954
rect 43260 24890 43312 24896
rect 43168 24608 43220 24614
rect 43168 24550 43220 24556
rect 43260 23656 43312 23662
rect 43260 23598 43312 23604
rect 43272 23322 43300 23598
rect 43260 23316 43312 23322
rect 43260 23258 43312 23264
rect 43548 23118 43576 25434
rect 43536 23112 43588 23118
rect 43536 23054 43588 23060
rect 43076 22976 43128 22982
rect 43076 22918 43128 22924
rect 41880 16176 41932 16182
rect 41880 16118 41932 16124
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 39764 15904 39816 15910
rect 39764 15846 39816 15852
rect 39120 15564 39172 15570
rect 39120 15506 39172 15512
rect 39776 15366 39804 15846
rect 41616 15706 41644 15982
rect 42248 15904 42300 15910
rect 42248 15846 42300 15852
rect 41604 15700 41656 15706
rect 41604 15642 41656 15648
rect 42260 15570 42288 15846
rect 40684 15564 40736 15570
rect 40684 15506 40736 15512
rect 42248 15564 42300 15570
rect 42248 15506 42300 15512
rect 38752 15360 38804 15366
rect 38752 15302 38804 15308
rect 39028 15360 39080 15366
rect 39028 15302 39080 15308
rect 39764 15360 39816 15366
rect 39764 15302 39816 15308
rect 38660 14408 38712 14414
rect 38660 14350 38712 14356
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 38764 13394 38792 15302
rect 40696 13802 40724 15506
rect 43640 13802 43668 31726
rect 43904 31340 43956 31346
rect 43904 31282 43956 31288
rect 43916 29782 43944 31282
rect 43996 29844 44048 29850
rect 43996 29786 44048 29792
rect 43904 29776 43956 29782
rect 43904 29718 43956 29724
rect 43904 29640 43956 29646
rect 43904 29582 43956 29588
rect 43812 29504 43864 29510
rect 43812 29446 43864 29452
rect 43824 29306 43852 29446
rect 43916 29306 43944 29582
rect 43812 29300 43864 29306
rect 43812 29242 43864 29248
rect 43904 29300 43956 29306
rect 43904 29242 43956 29248
rect 43718 29200 43774 29209
rect 43718 29135 43720 29144
rect 43772 29135 43774 29144
rect 43720 29106 43772 29112
rect 43812 29096 43864 29102
rect 43812 29038 43864 29044
rect 43904 29096 43956 29102
rect 44008 29084 44036 29786
rect 44088 29708 44140 29714
rect 44088 29650 44140 29656
rect 44100 29102 44128 29650
rect 43956 29056 44036 29084
rect 43904 29038 43956 29044
rect 43824 28422 43852 29038
rect 43904 28960 43956 28966
rect 43904 28902 43956 28908
rect 43812 28416 43864 28422
rect 43812 28358 43864 28364
rect 43916 28082 43944 28902
rect 44008 28558 44036 29056
rect 44088 29096 44140 29102
rect 44088 29038 44140 29044
rect 44088 28688 44140 28694
rect 44088 28630 44140 28636
rect 43996 28552 44048 28558
rect 43996 28494 44048 28500
rect 44100 28218 44128 28630
rect 44180 28416 44232 28422
rect 44180 28358 44232 28364
rect 44192 28218 44220 28358
rect 44088 28212 44140 28218
rect 44088 28154 44140 28160
rect 44180 28212 44232 28218
rect 44180 28154 44232 28160
rect 43904 28076 43956 28082
rect 43904 28018 43956 28024
rect 44180 27872 44232 27878
rect 44180 27814 44232 27820
rect 43996 26988 44048 26994
rect 43996 26930 44048 26936
rect 44008 26586 44036 26930
rect 43996 26580 44048 26586
rect 43996 26522 44048 26528
rect 43720 26308 43772 26314
rect 43720 26250 43772 26256
rect 43732 24682 43760 26250
rect 44008 25786 44036 26522
rect 44192 25906 44220 27814
rect 44180 25900 44232 25906
rect 44180 25842 44232 25848
rect 43916 25770 44036 25786
rect 43904 25764 44036 25770
rect 43956 25758 44036 25764
rect 43904 25706 43956 25712
rect 43720 24676 43772 24682
rect 43720 24618 43772 24624
rect 43732 24138 43760 24618
rect 43720 24132 43772 24138
rect 43720 24074 43772 24080
rect 44284 16574 44312 33390
rect 44548 31680 44600 31686
rect 44548 31622 44600 31628
rect 44560 31346 44588 31622
rect 44548 31340 44600 31346
rect 44548 31282 44600 31288
rect 45282 25256 45338 25265
rect 45282 25191 45338 25200
rect 44364 25152 44416 25158
rect 44364 25094 44416 25100
rect 44376 24274 44404 25094
rect 44548 24608 44600 24614
rect 44548 24550 44600 24556
rect 44560 24410 44588 24550
rect 44548 24404 44600 24410
rect 44548 24346 44600 24352
rect 44364 24268 44416 24274
rect 44364 24210 44416 24216
rect 44560 23866 44588 24346
rect 45296 23866 45324 25191
rect 44548 23860 44600 23866
rect 44548 23802 44600 23808
rect 45284 23860 45336 23866
rect 45284 23802 45336 23808
rect 44640 23520 44692 23526
rect 44640 23462 44692 23468
rect 44652 17066 44680 23462
rect 44640 17060 44692 17066
rect 44640 17002 44692 17008
rect 44548 16584 44600 16590
rect 44284 16546 44404 16574
rect 44376 16046 44404 16546
rect 44548 16526 44600 16532
rect 44364 16040 44416 16046
rect 44364 15982 44416 15988
rect 43812 15972 43864 15978
rect 43812 15914 43864 15920
rect 43824 15706 43852 15914
rect 43996 15904 44048 15910
rect 43996 15846 44048 15852
rect 43812 15700 43864 15706
rect 43812 15642 43864 15648
rect 44008 15162 44036 15846
rect 43996 15156 44048 15162
rect 43996 15098 44048 15104
rect 40684 13796 40736 13802
rect 40684 13738 40736 13744
rect 41236 13796 41288 13802
rect 41236 13738 41288 13744
rect 43628 13796 43680 13802
rect 43628 13738 43680 13744
rect 39580 13728 39632 13734
rect 39580 13670 39632 13676
rect 39592 13394 39620 13670
rect 38752 13388 38804 13394
rect 38752 13330 38804 13336
rect 39580 13388 39632 13394
rect 39580 13330 39632 13336
rect 37924 13320 37976 13326
rect 37924 13262 37976 13268
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 37936 12986 37964 13262
rect 37924 12980 37976 12986
rect 37924 12922 37976 12928
rect 37752 12406 37872 12434
rect 37844 12306 37872 12406
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37832 12300 37884 12306
rect 37832 12242 37884 12248
rect 37476 11762 37504 12242
rect 39040 12170 39068 13262
rect 40500 13184 40552 13190
rect 40500 13126 40552 13132
rect 40512 12986 40540 13126
rect 40500 12980 40552 12986
rect 40500 12922 40552 12928
rect 40696 12782 40724 13738
rect 41248 13394 41276 13738
rect 41236 13388 41288 13394
rect 41236 13330 41288 13336
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 40684 12776 40736 12782
rect 40684 12718 40736 12724
rect 39028 12164 39080 12170
rect 39028 12106 39080 12112
rect 37464 11756 37516 11762
rect 37384 11716 37464 11744
rect 37384 11354 37412 11716
rect 37464 11698 37516 11704
rect 37372 11348 37424 11354
rect 37372 11290 37424 11296
rect 38568 11280 38620 11286
rect 38568 11222 38620 11228
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 37188 9580 37240 9586
rect 37188 9522 37240 9528
rect 37096 8832 37148 8838
rect 37096 8774 37148 8780
rect 37004 8560 37056 8566
rect 37004 8502 37056 8508
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36912 7880 36964 7886
rect 36912 7822 36964 7828
rect 36740 7546 36768 7822
rect 37108 7818 37136 8774
rect 37096 7812 37148 7818
rect 37096 7754 37148 7760
rect 36820 7744 36872 7750
rect 36820 7686 36872 7692
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36832 7002 36860 7686
rect 36912 7404 36964 7410
rect 36912 7346 36964 7352
rect 37004 7404 37056 7410
rect 37004 7346 37056 7352
rect 36820 6996 36872 7002
rect 36820 6938 36872 6944
rect 36728 6724 36780 6730
rect 36728 6666 36780 6672
rect 36544 6112 36596 6118
rect 36544 6054 36596 6060
rect 36556 5234 36584 6054
rect 36740 5234 36768 6666
rect 36924 6458 36952 7346
rect 37016 6730 37044 7346
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 36912 6452 36964 6458
rect 36912 6394 36964 6400
rect 37108 6390 37136 7754
rect 37292 7546 37320 9930
rect 37384 9722 37412 10610
rect 37832 10600 37884 10606
rect 37832 10542 37884 10548
rect 37556 9988 37608 9994
rect 37556 9930 37608 9936
rect 37372 9716 37424 9722
rect 37372 9658 37424 9664
rect 37384 9178 37412 9658
rect 37568 9518 37596 9930
rect 37844 9518 37872 10542
rect 38384 10464 38436 10470
rect 38384 10406 38436 10412
rect 38396 9518 38424 10406
rect 38580 9518 38608 11222
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 38844 11076 38896 11082
rect 38844 11018 38896 11024
rect 38856 10674 38884 11018
rect 38844 10668 38896 10674
rect 38844 10610 38896 10616
rect 38856 9994 38884 10610
rect 38844 9988 38896 9994
rect 38844 9930 38896 9936
rect 38842 9616 38898 9625
rect 38842 9551 38844 9560
rect 38896 9551 38898 9560
rect 38844 9522 38896 9528
rect 37556 9512 37608 9518
rect 37556 9454 37608 9460
rect 37832 9512 37884 9518
rect 37832 9454 37884 9460
rect 38384 9512 38436 9518
rect 38384 9454 38436 9460
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 38396 8974 38424 9454
rect 38580 9178 38608 9454
rect 38948 9178 38976 11086
rect 39120 11008 39172 11014
rect 39120 10950 39172 10956
rect 39132 10810 39160 10950
rect 39120 10804 39172 10810
rect 39120 10746 39172 10752
rect 40696 10674 40724 12718
rect 41340 12714 41368 13262
rect 43812 13252 43864 13258
rect 43812 13194 43864 13200
rect 43824 12986 43852 13194
rect 44376 13190 44404 15982
rect 44560 15162 44588 16526
rect 44732 16448 44784 16454
rect 44730 16416 44732 16425
rect 44784 16416 44786 16425
rect 44730 16351 44786 16360
rect 44548 15156 44600 15162
rect 44548 15098 44600 15104
rect 44364 13184 44416 13190
rect 44364 13126 44416 13132
rect 43812 12980 43864 12986
rect 43812 12922 43864 12928
rect 44376 12918 44404 13126
rect 44364 12912 44416 12918
rect 44364 12854 44416 12860
rect 41328 12708 41380 12714
rect 41328 12650 41380 12656
rect 44640 12708 44692 12714
rect 44640 12650 44692 12656
rect 40684 10668 40736 10674
rect 40684 10610 40736 10616
rect 40224 10600 40276 10606
rect 40224 10542 40276 10548
rect 40236 10266 40264 10542
rect 41236 10464 41288 10470
rect 41236 10406 41288 10412
rect 40224 10260 40276 10266
rect 40224 10202 40276 10208
rect 41248 10130 41276 10406
rect 39212 10124 39264 10130
rect 39212 10066 39264 10072
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 43628 10124 43680 10130
rect 43628 10066 43680 10072
rect 39028 9920 39080 9926
rect 39028 9862 39080 9868
rect 39040 9450 39068 9862
rect 39120 9648 39172 9654
rect 39118 9616 39120 9625
rect 39172 9616 39174 9625
rect 39118 9551 39174 9560
rect 39028 9444 39080 9450
rect 39028 9386 39080 9392
rect 38568 9172 38620 9178
rect 38568 9114 38620 9120
rect 38936 9172 38988 9178
rect 38936 9114 38988 9120
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 39040 8906 39068 9386
rect 39120 9376 39172 9382
rect 39120 9318 39172 9324
rect 39028 8900 39080 8906
rect 39028 8842 39080 8848
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37556 7744 37608 7750
rect 37556 7686 37608 7692
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37096 6384 37148 6390
rect 37096 6326 37148 6332
rect 37292 5302 37320 7482
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37384 7002 37412 7346
rect 37372 6996 37424 7002
rect 37372 6938 37424 6944
rect 37476 6866 37504 7686
rect 37568 7342 37596 7686
rect 37556 7336 37608 7342
rect 37556 7278 37608 7284
rect 37568 6866 37596 7278
rect 37648 7268 37700 7274
rect 37648 7210 37700 7216
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 37556 6860 37608 6866
rect 37556 6802 37608 6808
rect 37476 6254 37504 6802
rect 37464 6248 37516 6254
rect 37464 6190 37516 6196
rect 37568 6118 37596 6802
rect 37660 6390 37688 7210
rect 37752 7206 37780 7822
rect 38660 7812 38712 7818
rect 38660 7754 38712 7760
rect 37740 7200 37792 7206
rect 37740 7142 37792 7148
rect 37648 6384 37700 6390
rect 37648 6326 37700 6332
rect 37660 6254 37688 6326
rect 37752 6322 37780 7142
rect 37924 6792 37976 6798
rect 37924 6734 37976 6740
rect 37936 6458 37964 6734
rect 38200 6656 38252 6662
rect 38200 6598 38252 6604
rect 38292 6656 38344 6662
rect 38292 6598 38344 6604
rect 38212 6458 38240 6598
rect 38304 6458 38332 6598
rect 37924 6452 37976 6458
rect 37924 6394 37976 6400
rect 38200 6452 38252 6458
rect 38200 6394 38252 6400
rect 38292 6452 38344 6458
rect 38292 6394 38344 6400
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 38672 6254 38700 7754
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38764 7478 38792 7686
rect 38752 7472 38804 7478
rect 38752 7414 38804 7420
rect 39132 7410 39160 9318
rect 39224 8838 39252 10066
rect 39304 10056 39356 10062
rect 39304 9998 39356 10004
rect 39316 9722 39344 9998
rect 40868 9988 40920 9994
rect 40868 9930 40920 9936
rect 43168 9988 43220 9994
rect 43168 9930 43220 9936
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 39304 9716 39356 9722
rect 39304 9658 39356 9664
rect 39868 9518 39896 9862
rect 40880 9674 40908 9930
rect 41696 9920 41748 9926
rect 41696 9862 41748 9868
rect 42156 9920 42208 9926
rect 42156 9862 42208 9868
rect 40604 9646 40908 9674
rect 39856 9512 39908 9518
rect 39856 9454 39908 9460
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 39316 9178 39344 9318
rect 39304 9172 39356 9178
rect 39304 9114 39356 9120
rect 39488 8900 39540 8906
rect 39488 8842 39540 8848
rect 39212 8832 39264 8838
rect 39212 8774 39264 8780
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39212 7472 39264 7478
rect 39212 7414 39264 7420
rect 39120 7404 39172 7410
rect 39120 7346 39172 7352
rect 38752 7336 38804 7342
rect 38752 7278 38804 7284
rect 39028 7336 39080 7342
rect 39028 7278 39080 7284
rect 38764 6254 38792 7278
rect 37648 6248 37700 6254
rect 37648 6190 37700 6196
rect 38660 6248 38712 6254
rect 38660 6190 38712 6196
rect 38752 6248 38804 6254
rect 38752 6190 38804 6196
rect 37556 6112 37608 6118
rect 37556 6054 37608 6060
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 37280 5296 37332 5302
rect 37280 5238 37332 5244
rect 36544 5228 36596 5234
rect 36544 5170 36596 5176
rect 36728 5228 36780 5234
rect 36728 5170 36780 5176
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 35716 4072 35768 4078
rect 35716 4014 35768 4020
rect 35624 3732 35676 3738
rect 35624 3674 35676 3680
rect 35532 3120 35584 3126
rect 35532 3062 35584 3068
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35728 2854 35756 4014
rect 35912 3602 35940 4082
rect 36096 4010 36124 5102
rect 36452 5092 36504 5098
rect 36452 5034 36504 5040
rect 36176 5024 36228 5030
rect 36176 4966 36228 4972
rect 36188 4826 36216 4966
rect 36176 4820 36228 4826
rect 36176 4762 36228 4768
rect 36266 4312 36322 4321
rect 36188 4270 36266 4298
rect 36188 4214 36216 4270
rect 36266 4247 36322 4256
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 36464 4078 36492 5034
rect 36740 4554 36768 5170
rect 36728 4548 36780 4554
rect 36728 4490 36780 4496
rect 36544 4480 36596 4486
rect 36544 4422 36596 4428
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 36084 4004 36136 4010
rect 36084 3946 36136 3952
rect 36556 3942 36584 4422
rect 36634 4312 36690 4321
rect 36634 4247 36636 4256
rect 36688 4247 36690 4256
rect 36636 4218 36688 4224
rect 36740 4010 36768 4490
rect 37188 4480 37240 4486
rect 37188 4422 37240 4428
rect 37200 4298 37228 4422
rect 37200 4270 37320 4298
rect 37188 4208 37240 4214
rect 37188 4150 37240 4156
rect 37096 4140 37148 4146
rect 37096 4082 37148 4088
rect 36728 4004 36780 4010
rect 36728 3946 36780 3952
rect 36912 4004 36964 4010
rect 36912 3946 36964 3952
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36740 3058 36768 3946
rect 36924 3602 36952 3946
rect 37108 3738 37136 4082
rect 37096 3732 37148 3738
rect 37096 3674 37148 3680
rect 37200 3602 37228 4150
rect 37292 4078 37320 4270
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 37384 3670 37412 5646
rect 38028 4826 38056 5646
rect 38672 5114 38700 6190
rect 38752 5364 38804 5370
rect 38752 5306 38804 5312
rect 38764 5234 38792 5306
rect 39040 5234 39068 7278
rect 39132 6798 39160 7346
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 39224 6662 39252 7414
rect 39316 7002 39344 7822
rect 39500 7206 39528 8842
rect 40604 8498 40632 9646
rect 41708 9042 41736 9862
rect 41880 9648 41932 9654
rect 41880 9590 41932 9596
rect 41892 9178 41920 9590
rect 42168 9586 42196 9862
rect 43180 9722 43208 9930
rect 43168 9716 43220 9722
rect 43168 9658 43220 9664
rect 42156 9580 42208 9586
rect 42156 9522 42208 9528
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 42064 9444 42116 9450
rect 42064 9386 42116 9392
rect 41880 9172 41932 9178
rect 41880 9114 41932 9120
rect 41696 9036 41748 9042
rect 41696 8978 41748 8984
rect 41708 8566 41736 8978
rect 41972 8968 42024 8974
rect 41972 8910 42024 8916
rect 41984 8566 42012 8910
rect 42076 8906 42104 9386
rect 42720 9042 42748 9522
rect 42708 9036 42760 9042
rect 42708 8978 42760 8984
rect 42248 8968 42300 8974
rect 42248 8910 42300 8916
rect 42616 8968 42668 8974
rect 42616 8910 42668 8916
rect 42064 8900 42116 8906
rect 42064 8842 42116 8848
rect 42260 8634 42288 8910
rect 42628 8634 42656 8910
rect 42248 8628 42300 8634
rect 42248 8570 42300 8576
rect 42616 8628 42668 8634
rect 42616 8570 42668 8576
rect 41696 8560 41748 8566
rect 41696 8502 41748 8508
rect 41972 8560 42024 8566
rect 41972 8502 42024 8508
rect 40408 8492 40460 8498
rect 40408 8434 40460 8440
rect 40592 8492 40644 8498
rect 40592 8434 40644 8440
rect 40316 8288 40368 8294
rect 40316 8230 40368 8236
rect 40328 8090 40356 8230
rect 40316 8084 40368 8090
rect 40316 8026 40368 8032
rect 40224 7744 40276 7750
rect 40224 7686 40276 7692
rect 40236 7478 40264 7686
rect 40224 7472 40276 7478
rect 40224 7414 40276 7420
rect 40420 7410 40448 8434
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 41236 8288 41288 8294
rect 41236 8230 41288 8236
rect 41248 7886 41276 8230
rect 41236 7880 41288 7886
rect 41236 7822 41288 7828
rect 41432 7750 41460 8366
rect 41420 7744 41472 7750
rect 41420 7686 41472 7692
rect 39580 7404 39632 7410
rect 39580 7346 39632 7352
rect 40408 7404 40460 7410
rect 40408 7346 40460 7352
rect 41328 7404 41380 7410
rect 41328 7346 41380 7352
rect 39488 7200 39540 7206
rect 39488 7142 39540 7148
rect 39304 6996 39356 7002
rect 39304 6938 39356 6944
rect 39212 6656 39264 6662
rect 39212 6598 39264 6604
rect 38752 5228 38804 5234
rect 38752 5170 38804 5176
rect 39028 5228 39080 5234
rect 39028 5170 39080 5176
rect 39212 5228 39264 5234
rect 39212 5170 39264 5176
rect 38672 5086 38884 5114
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37844 4282 37872 4558
rect 37936 4536 37964 4762
rect 38752 4752 38804 4758
rect 38752 4694 38804 4700
rect 38016 4548 38068 4554
rect 37936 4508 38016 4536
rect 38016 4490 38068 4496
rect 37832 4276 37884 4282
rect 37832 4218 37884 4224
rect 38028 4078 38056 4490
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4146 38240 4422
rect 38764 4282 38792 4694
rect 38856 4690 38884 5086
rect 38844 4684 38896 4690
rect 38844 4626 38896 4632
rect 38752 4276 38804 4282
rect 38752 4218 38804 4224
rect 38200 4140 38252 4146
rect 38200 4082 38252 4088
rect 38016 4072 38068 4078
rect 38016 4014 38068 4020
rect 39120 4072 39172 4078
rect 39224 4060 39252 5170
rect 39500 4706 39528 7142
rect 39592 6730 39620 7346
rect 39672 7268 39724 7274
rect 39672 7210 39724 7216
rect 39684 6798 39712 7210
rect 39672 6792 39724 6798
rect 39672 6734 39724 6740
rect 39580 6724 39632 6730
rect 39580 6666 39632 6672
rect 39592 5914 39620 6666
rect 39580 5908 39632 5914
rect 39580 5850 39632 5856
rect 41340 5370 41368 7346
rect 41432 7342 41460 7686
rect 41708 7546 41736 8502
rect 42064 8288 42116 8294
rect 42064 8230 42116 8236
rect 42432 8288 42484 8294
rect 42432 8230 42484 8236
rect 42076 8090 42104 8230
rect 42064 8084 42116 8090
rect 42064 8026 42116 8032
rect 41696 7540 41748 7546
rect 41696 7482 41748 7488
rect 42076 7410 42104 8026
rect 42248 7540 42300 7546
rect 42248 7482 42300 7488
rect 42260 7410 42288 7482
rect 42444 7410 42472 8230
rect 42720 7410 42748 8978
rect 42892 8968 42944 8974
rect 42892 8910 42944 8916
rect 41788 7404 41840 7410
rect 41788 7346 41840 7352
rect 42064 7404 42116 7410
rect 42064 7346 42116 7352
rect 42248 7404 42300 7410
rect 42248 7346 42300 7352
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 42708 7404 42760 7410
rect 42708 7346 42760 7352
rect 41420 7336 41472 7342
rect 41420 7278 41472 7284
rect 41800 6458 41828 7346
rect 42720 6866 42748 7346
rect 42800 6928 42852 6934
rect 42800 6870 42852 6876
rect 42708 6860 42760 6866
rect 42708 6802 42760 6808
rect 42720 6458 42748 6802
rect 42812 6458 42840 6870
rect 42904 6866 42932 8910
rect 43076 8900 43128 8906
rect 43076 8842 43128 8848
rect 43088 7818 43116 8842
rect 43352 8832 43404 8838
rect 43352 8774 43404 8780
rect 43076 7812 43128 7818
rect 43076 7754 43128 7760
rect 43364 6866 43392 8774
rect 43640 7886 43668 10066
rect 43720 8424 43772 8430
rect 43720 8366 43772 8372
rect 43628 7880 43680 7886
rect 43628 7822 43680 7828
rect 43444 7812 43496 7818
rect 43444 7754 43496 7760
rect 42892 6860 42944 6866
rect 42892 6802 42944 6808
rect 43076 6860 43128 6866
rect 43076 6802 43128 6808
rect 43352 6860 43404 6866
rect 43352 6802 43404 6808
rect 41788 6452 41840 6458
rect 41788 6394 41840 6400
rect 42708 6452 42760 6458
rect 42708 6394 42760 6400
rect 42800 6452 42852 6458
rect 42800 6394 42852 6400
rect 42248 6316 42300 6322
rect 42248 6258 42300 6264
rect 42892 6316 42944 6322
rect 42892 6258 42944 6264
rect 41328 5364 41380 5370
rect 41328 5306 41380 5312
rect 42156 5364 42208 5370
rect 42156 5306 42208 5312
rect 41512 5228 41564 5234
rect 41512 5170 41564 5176
rect 39580 5160 39632 5166
rect 39580 5102 39632 5108
rect 41052 5160 41104 5166
rect 41052 5102 41104 5108
rect 39592 4826 39620 5102
rect 41064 4826 41092 5102
rect 39580 4820 39632 4826
rect 39580 4762 39632 4768
rect 40868 4820 40920 4826
rect 40868 4762 40920 4768
rect 41052 4820 41104 4826
rect 41052 4762 41104 4768
rect 39500 4690 39620 4706
rect 39500 4684 39632 4690
rect 39500 4678 39580 4684
rect 39580 4626 39632 4632
rect 39304 4480 39356 4486
rect 39304 4422 39356 4428
rect 39172 4032 39252 4060
rect 39120 4014 39172 4020
rect 37372 3664 37424 3670
rect 37372 3606 37424 3612
rect 36912 3596 36964 3602
rect 36912 3538 36964 3544
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 37200 3194 37228 3538
rect 38028 3534 38056 4014
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 38396 3738 38424 3878
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 37556 3528 37608 3534
rect 37556 3470 37608 3476
rect 38016 3528 38068 3534
rect 38016 3470 38068 3476
rect 37568 3194 37596 3470
rect 38568 3392 38620 3398
rect 38568 3334 38620 3340
rect 37188 3188 37240 3194
rect 37188 3130 37240 3136
rect 37556 3188 37608 3194
rect 37556 3130 37608 3136
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 38580 2990 38608 3334
rect 39224 3194 39252 4032
rect 39316 3534 39344 4422
rect 39592 3602 39620 4626
rect 40040 4616 40092 4622
rect 40040 4558 40092 4564
rect 40052 4282 40080 4558
rect 40776 4548 40828 4554
rect 40880 4536 40908 4762
rect 41064 4622 41092 4762
rect 41052 4616 41104 4622
rect 40828 4508 40908 4536
rect 40776 4490 40828 4496
rect 40684 4480 40736 4486
rect 40684 4422 40736 4428
rect 40040 4276 40092 4282
rect 40040 4218 40092 4224
rect 40696 4146 40724 4422
rect 40880 4146 40908 4508
rect 40972 4576 41052 4604
rect 40972 4146 41000 4576
rect 41052 4558 41104 4564
rect 41328 4616 41380 4622
rect 41328 4558 41380 4564
rect 41420 4616 41472 4622
rect 41420 4558 41472 4564
rect 41340 4146 41368 4558
rect 41432 4282 41460 4558
rect 41524 4554 41552 5170
rect 41696 5092 41748 5098
rect 41696 5034 41748 5040
rect 41512 4548 41564 4554
rect 41512 4490 41564 4496
rect 41708 4486 41736 5034
rect 42168 4826 42196 5306
rect 42260 5234 42288 6258
rect 42248 5228 42300 5234
rect 42248 5170 42300 5176
rect 42156 4820 42208 4826
rect 42156 4762 42208 4768
rect 42260 4622 42288 5170
rect 42904 5166 42932 6258
rect 42984 6180 43036 6186
rect 42984 6122 43036 6128
rect 42892 5160 42944 5166
rect 42892 5102 42944 5108
rect 42248 4616 42300 4622
rect 42248 4558 42300 4564
rect 42904 4554 42932 5102
rect 42996 5030 43024 6122
rect 43088 5778 43116 6802
rect 43456 6730 43484 7754
rect 43640 7546 43668 7822
rect 43628 7540 43680 7546
rect 43628 7482 43680 7488
rect 43640 7018 43668 7482
rect 43732 7274 43760 8366
rect 43720 7268 43772 7274
rect 43720 7210 43772 7216
rect 43548 7002 43668 7018
rect 43536 6996 43668 7002
rect 43588 6990 43668 6996
rect 43536 6938 43588 6944
rect 43444 6724 43496 6730
rect 43444 6666 43496 6672
rect 43076 5772 43128 5778
rect 43076 5714 43128 5720
rect 42984 5024 43036 5030
rect 42984 4966 43036 4972
rect 41972 4548 42024 4554
rect 41972 4490 42024 4496
rect 42892 4548 42944 4554
rect 42892 4490 42944 4496
rect 41696 4480 41748 4486
rect 41696 4422 41748 4428
rect 41984 4434 42012 4490
rect 42800 4480 42852 4486
rect 41984 4406 42104 4434
rect 42800 4422 42852 4428
rect 41420 4276 41472 4282
rect 41420 4218 41472 4224
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 40684 4140 40736 4146
rect 40684 4082 40736 4088
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 40960 4140 41012 4146
rect 40960 4082 41012 4088
rect 41328 4140 41380 4146
rect 41328 4082 41380 4088
rect 40512 3738 40540 4082
rect 42076 4078 42104 4406
rect 42340 4140 42392 4146
rect 42340 4082 42392 4088
rect 42064 4072 42116 4078
rect 42064 4014 42116 4020
rect 41236 3936 41288 3942
rect 41236 3878 41288 3884
rect 40500 3732 40552 3738
rect 40500 3674 40552 3680
rect 39580 3596 39632 3602
rect 39580 3538 39632 3544
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 41248 3194 41276 3878
rect 42076 3194 42104 4014
rect 39212 3188 39264 3194
rect 39212 3130 39264 3136
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 42064 3188 42116 3194
rect 42064 3130 42116 3136
rect 42352 3126 42380 4082
rect 42812 4078 42840 4422
rect 42800 4072 42852 4078
rect 42800 4014 42852 4020
rect 43088 3942 43116 5714
rect 43456 5642 43484 6666
rect 44652 6458 44680 12650
rect 45282 6896 45338 6905
rect 45282 6831 45338 6840
rect 44640 6452 44692 6458
rect 44640 6394 44692 6400
rect 45296 6390 45324 6831
rect 45284 6384 45336 6390
rect 45284 6326 45336 6332
rect 43352 5636 43404 5642
rect 43352 5578 43404 5584
rect 43444 5636 43496 5642
rect 43444 5578 43496 5584
rect 43364 5370 43392 5578
rect 43352 5364 43404 5370
rect 43352 5306 43404 5312
rect 43168 4548 43220 4554
rect 43168 4490 43220 4496
rect 43180 4078 43208 4490
rect 43456 4282 43484 5578
rect 44824 5568 44876 5574
rect 44824 5510 44876 5516
rect 44836 5166 44864 5510
rect 44824 5160 44876 5166
rect 44824 5102 44876 5108
rect 43444 4276 43496 4282
rect 43444 4218 43496 4224
rect 43168 4072 43220 4078
rect 43168 4014 43220 4020
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42340 3120 42392 3126
rect 42340 3062 42392 3068
rect 38568 2984 38620 2990
rect 38568 2926 38620 2932
rect 43902 2952 43958 2961
rect 43902 2887 43958 2896
rect 35716 2848 35768 2854
rect 35716 2790 35768 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 43916 2650 43944 2887
rect 43904 2644 43956 2650
rect 43904 2586 43956 2592
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 26422 0 26478 800
rect 34794 0 34850 800
rect 43810 0 43866 800
<< via2 >>
rect 938 46280 994 46336
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 938 36760 994 36816
rect 938 27920 994 27976
rect 938 18400 994 18456
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 5814 28484 5870 28520
rect 5814 28464 5816 28484
rect 5816 28464 5868 28484
rect 5868 28464 5870 28484
rect 6550 30368 6606 30424
rect 6826 28600 6882 28656
rect 6458 28056 6514 28112
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 8114 27920 8170 27976
rect 8942 28484 8998 28520
rect 8942 28464 8944 28484
rect 8944 28464 8996 28484
rect 8996 28464 8998 28484
rect 10230 33904 10286 33960
rect 12162 33652 12218 33688
rect 12162 33632 12164 33652
rect 12164 33632 12216 33652
rect 12216 33632 12218 33652
rect 12346 31728 12402 31784
rect 12254 30676 12256 30696
rect 12256 30676 12308 30696
rect 12308 30676 12310 30696
rect 12254 30640 12310 30676
rect 11334 30368 11390 30424
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 11242 23604 11244 23624
rect 11244 23604 11296 23624
rect 11296 23604 11298 23624
rect 11242 23568 11298 23604
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 13174 31900 13176 31920
rect 13176 31900 13228 31920
rect 13228 31900 13230 31920
rect 13174 31864 13230 31900
rect 12530 28600 12586 28656
rect 12438 27920 12494 27976
rect 13726 34040 13782 34096
rect 13174 28872 13230 28928
rect 13634 28076 13690 28112
rect 13634 28056 13636 28076
rect 13636 28056 13688 28076
rect 13688 28056 13690 28076
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 10690 15700 10746 15736
rect 10690 15680 10692 15700
rect 10692 15680 10744 15700
rect 10744 15680 10746 15700
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 10690 14320 10746 14376
rect 11426 15428 11482 15464
rect 11426 15408 11428 15428
rect 11428 15408 11480 15428
rect 11480 15408 11482 15428
rect 11978 14864 12034 14920
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 14278 31728 14334 31784
rect 15474 31728 15530 31784
rect 14830 30660 14886 30696
rect 14830 30640 14832 30660
rect 14832 30640 14884 30660
rect 14884 30640 14886 30660
rect 15290 23568 15346 23624
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 17130 33632 17186 33688
rect 16578 28872 16634 28928
rect 11518 11056 11574 11112
rect 11058 10260 11114 10296
rect 11058 10240 11060 10260
rect 11060 10240 11112 10260
rect 11112 10240 11114 10260
rect 12530 12416 12586 12472
rect 12530 12044 12532 12064
rect 12532 12044 12584 12064
rect 12584 12044 12586 12064
rect 12530 12008 12586 12044
rect 11794 11464 11850 11520
rect 12346 9424 12402 9480
rect 13266 13776 13322 13832
rect 13266 10376 13322 10432
rect 12714 9560 12770 9616
rect 12990 9424 13046 9480
rect 12346 6568 12402 6624
rect 12530 5616 12586 5672
rect 13726 12144 13782 12200
rect 14278 15816 14334 15872
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 18050 31864 18106 31920
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19338 31728 19394 31784
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 21178 33924 21234 33960
rect 21178 33904 21180 33924
rect 21180 33904 21232 33924
rect 21232 33904 21234 33924
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 14830 15816 14886 15872
rect 14554 15544 14610 15600
rect 14002 13812 14004 13832
rect 14004 13812 14056 13832
rect 14056 13812 14058 13832
rect 14002 13776 14058 13812
rect 14002 12552 14058 12608
rect 14278 13932 14334 13968
rect 14278 13912 14280 13932
rect 14280 13912 14332 13932
rect 14332 13912 14334 13932
rect 14738 14184 14794 14240
rect 13818 11600 13874 11656
rect 13818 10784 13874 10840
rect 14094 9968 14150 10024
rect 13542 6840 13598 6896
rect 15566 14592 15622 14648
rect 15198 12688 15254 12744
rect 15198 12008 15254 12064
rect 15014 11328 15070 11384
rect 15290 11756 15346 11792
rect 15290 11736 15292 11756
rect 15292 11736 15344 11756
rect 15344 11736 15346 11756
rect 15382 10920 15438 10976
rect 15658 12724 15660 12744
rect 15660 12724 15712 12744
rect 15712 12724 15714 12744
rect 15658 12688 15714 12724
rect 15658 12552 15714 12608
rect 16118 15816 16174 15872
rect 15842 13776 15898 13832
rect 15750 9560 15806 9616
rect 15474 6316 15530 6352
rect 16670 13912 16726 13968
rect 16486 11600 16542 11656
rect 17038 14764 17040 14784
rect 17040 14764 17092 14784
rect 17092 14764 17094 14784
rect 17038 14728 17094 14764
rect 17222 15272 17278 15328
rect 17130 14456 17186 14512
rect 17682 15000 17738 15056
rect 17590 14864 17646 14920
rect 17590 14764 17592 14784
rect 17592 14764 17644 14784
rect 17644 14764 17646 14784
rect 17590 14728 17646 14764
rect 17314 13812 17316 13832
rect 17316 13812 17368 13832
rect 17368 13812 17370 13832
rect 17314 13776 17370 13812
rect 16486 9560 16542 9616
rect 17038 10240 17094 10296
rect 16670 8900 16726 8936
rect 16670 8880 16672 8900
rect 16672 8880 16724 8900
rect 16724 8880 16726 8900
rect 16486 6840 16542 6896
rect 17958 14592 18014 14648
rect 17682 12552 17738 12608
rect 17222 11056 17278 11112
rect 17314 10784 17370 10840
rect 17222 10376 17278 10432
rect 17222 9580 17278 9616
rect 17222 9560 17224 9580
rect 17224 9560 17276 9580
rect 17276 9560 17278 9580
rect 17222 8880 17278 8936
rect 15474 6296 15476 6316
rect 15476 6296 15528 6316
rect 15528 6296 15530 6316
rect 17130 6568 17186 6624
rect 17958 11092 17960 11112
rect 17960 11092 18012 11112
rect 18012 11092 18014 11112
rect 17958 11056 18014 11092
rect 18602 15680 18658 15736
rect 18602 14184 18658 14240
rect 18326 11192 18382 11248
rect 17866 9968 17922 10024
rect 18602 10920 18658 10976
rect 18418 9424 18474 9480
rect 18326 6840 18382 6896
rect 18602 9152 18658 9208
rect 18970 11328 19026 11384
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19154 14456 19210 14512
rect 18970 11056 19026 11112
rect 19154 11076 19210 11112
rect 19154 11056 19156 11076
rect 19156 11056 19208 11076
rect 19208 11056 19210 11076
rect 19798 15680 19854 15736
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19522 15000 19578 15056
rect 24398 34040 24454 34096
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19522 12688 19578 12744
rect 20074 12280 20130 12336
rect 19706 12180 19708 12200
rect 19708 12180 19760 12200
rect 19760 12180 19762 12200
rect 19706 12144 19762 12180
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20074 12008 20130 12064
rect 19706 11600 19762 11656
rect 19614 11464 19670 11520
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19430 10140 19432 10160
rect 19432 10140 19484 10160
rect 19484 10140 19486 10160
rect 19430 10104 19486 10140
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19522 9632 19578 9688
rect 19338 9152 19394 9208
rect 19614 9288 19670 9344
rect 19982 9424 20038 9480
rect 20074 9152 20130 9208
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19062 6296 19118 6352
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 21178 19216 21234 19272
rect 21914 19216 21970 19272
rect 21638 15564 21694 15600
rect 21638 15544 21640 15564
rect 21640 15544 21692 15564
rect 21692 15544 21694 15564
rect 20442 11328 20498 11384
rect 20626 12144 20682 12200
rect 20626 11600 20682 11656
rect 20350 10004 20352 10024
rect 20352 10004 20404 10024
rect 20404 10004 20406 10024
rect 20350 9968 20406 10004
rect 20350 9832 20406 9888
rect 20350 8200 20406 8256
rect 20994 11736 21050 11792
rect 20718 9832 20774 9888
rect 17590 5636 17646 5672
rect 17590 5616 17592 5636
rect 17592 5616 17644 5636
rect 17644 5616 17646 5636
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 22466 17992 22522 18048
rect 22650 16632 22706 16688
rect 22098 15444 22100 15464
rect 22100 15444 22152 15464
rect 22152 15444 22154 15464
rect 22098 15408 22154 15444
rect 22374 15680 22430 15736
rect 22742 15408 22798 15464
rect 22374 12824 22430 12880
rect 22650 13776 22706 13832
rect 22558 10920 22614 10976
rect 22558 9988 22614 10024
rect 22558 9968 22560 9988
rect 22560 9968 22612 9988
rect 22612 9968 22614 9988
rect 22558 9560 22614 9616
rect 23386 15428 23442 15464
rect 23386 15408 23388 15428
rect 23388 15408 23440 15428
rect 23440 15408 23442 15428
rect 24122 15680 24178 15736
rect 23294 8084 23350 8120
rect 23294 8064 23296 8084
rect 23296 8064 23348 8084
rect 23348 8064 23350 8084
rect 26698 42064 26754 42120
rect 27066 37168 27122 37224
rect 27342 36252 27344 36272
rect 27344 36252 27396 36272
rect 27396 36252 27398 36272
rect 27342 36216 27398 36252
rect 28814 42064 28870 42120
rect 29642 41248 29698 41304
rect 30102 41676 30158 41712
rect 30102 41656 30104 41676
rect 30104 41656 30156 41676
rect 30156 41656 30158 41676
rect 31114 41012 31116 41032
rect 31116 41012 31168 41032
rect 31168 41012 31170 41032
rect 31114 40976 31170 41012
rect 31574 41148 31576 41168
rect 31576 41148 31628 41168
rect 31628 41148 31630 41168
rect 31574 41112 31630 41148
rect 30102 33088 30158 33144
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 32126 40976 32182 41032
rect 32586 41656 32642 41712
rect 32494 41148 32496 41168
rect 32496 41148 32548 41168
rect 32548 41148 32550 41168
rect 32494 41112 32550 41148
rect 33598 41540 33654 41576
rect 33598 41520 33600 41540
rect 33600 41520 33652 41540
rect 33652 41520 33654 41540
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34334 41540 34390 41576
rect 34334 41520 34336 41540
rect 34336 41520 34388 41540
rect 34388 41520 34390 41540
rect 35070 41268 35126 41304
rect 35070 41248 35072 41268
rect 35072 41248 35124 41268
rect 35124 41248 35126 41268
rect 31666 19916 31722 19952
rect 31666 19896 31668 19916
rect 31668 19896 31720 19916
rect 31720 19896 31722 19916
rect 33598 34604 33654 34640
rect 33598 34584 33600 34604
rect 33600 34584 33652 34604
rect 33652 34584 33654 34604
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34334 36216 34390 36272
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 36174 37168 36230 37224
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 38658 38528 38714 38584
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 39302 38528 39358 38584
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 32310 19896 32366 19952
rect 33874 19372 33930 19408
rect 33874 19352 33876 19372
rect 33876 19352 33928 19372
rect 33928 19352 33930 19372
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 29550 9152 29606 9208
rect 30378 14356 30380 14376
rect 30380 14356 30432 14376
rect 30432 14356 30434 14376
rect 30378 14320 30434 14356
rect 29918 9696 29974 9752
rect 30746 11192 30802 11248
rect 30102 9052 30104 9072
rect 30104 9052 30156 9072
rect 30156 9052 30158 9072
rect 30102 9016 30158 9052
rect 30286 9172 30342 9208
rect 30286 9152 30288 9172
rect 30288 9152 30340 9172
rect 30340 9152 30342 9172
rect 30838 9052 30840 9072
rect 30840 9052 30892 9072
rect 30892 9052 30894 9072
rect 30838 9016 30894 9052
rect 31390 11092 31392 11112
rect 31392 11092 31444 11112
rect 31444 11092 31446 11112
rect 31390 11056 31446 11092
rect 31850 11056 31906 11112
rect 31666 9696 31722 9752
rect 32126 11192 32182 11248
rect 30838 2916 30894 2952
rect 30838 2896 30840 2916
rect 30840 2896 30892 2916
rect 30892 2896 30894 2916
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35806 19352 35862 19408
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 41786 29144 41842 29200
rect 45282 44240 45338 44296
rect 45282 34720 45338 34776
rect 43718 29164 43774 29200
rect 43718 29144 43720 29164
rect 43720 29144 43772 29164
rect 43772 29144 43774 29164
rect 45282 25200 45338 25256
rect 38842 9580 38898 9616
rect 38842 9560 38844 9580
rect 38844 9560 38896 9580
rect 38896 9560 38898 9580
rect 44730 16396 44732 16416
rect 44732 16396 44784 16416
rect 44784 16396 44786 16416
rect 44730 16360 44786 16396
rect 39118 9596 39120 9616
rect 39120 9596 39172 9616
rect 39172 9596 39174 9616
rect 39118 9560 39174 9596
rect 36266 4256 36322 4312
rect 36634 4276 36690 4312
rect 36634 4256 36636 4276
rect 36636 4256 36688 4276
rect 36688 4256 36690 4276
rect 45282 6840 45338 6896
rect 43902 2896 43958 2952
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 0 46338 800 46368
rect 933 46338 999 46341
rect 0 46336 999 46338
rect 0 46280 938 46336
rect 994 46280 999 46336
rect 0 46278 999 46280
rect 0 46248 800 46278
rect 933 46275 999 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 45277 44298 45343 44301
rect 45537 44298 46337 44328
rect 45277 44296 46337 44298
rect 45277 44240 45282 44296
rect 45338 44240 46337 44296
rect 45277 44238 46337 44240
rect 45277 44235 45343 44238
rect 45537 44208 46337 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 26693 42122 26759 42125
rect 28809 42122 28875 42125
rect 26693 42120 28875 42122
rect 26693 42064 26698 42120
rect 26754 42064 28814 42120
rect 28870 42064 28875 42120
rect 26693 42062 28875 42064
rect 26693 42059 26759 42062
rect 28809 42059 28875 42062
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 30097 41714 30163 41717
rect 32581 41714 32647 41717
rect 30097 41712 32647 41714
rect 30097 41656 30102 41712
rect 30158 41656 32586 41712
rect 32642 41656 32647 41712
rect 30097 41654 32647 41656
rect 30097 41651 30163 41654
rect 32581 41651 32647 41654
rect 33593 41578 33659 41581
rect 34329 41578 34395 41581
rect 33593 41576 34395 41578
rect 33593 41520 33598 41576
rect 33654 41520 34334 41576
rect 34390 41520 34395 41576
rect 33593 41518 34395 41520
rect 33593 41515 33659 41518
rect 34329 41515 34395 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 29637 41306 29703 41309
rect 35065 41306 35131 41309
rect 29637 41304 35131 41306
rect 29637 41248 29642 41304
rect 29698 41248 35070 41304
rect 35126 41248 35131 41304
rect 29637 41246 35131 41248
rect 29637 41243 29703 41246
rect 35065 41243 35131 41246
rect 31569 41170 31635 41173
rect 32489 41170 32555 41173
rect 31569 41168 32555 41170
rect 31569 41112 31574 41168
rect 31630 41112 32494 41168
rect 32550 41112 32555 41168
rect 31569 41110 32555 41112
rect 31569 41107 31635 41110
rect 32489 41107 32555 41110
rect 31109 41034 31175 41037
rect 32121 41034 32187 41037
rect 31109 41032 32187 41034
rect 31109 40976 31114 41032
rect 31170 40976 32126 41032
rect 32182 40976 32187 41032
rect 31109 40974 32187 40976
rect 31109 40971 31175 40974
rect 32121 40971 32187 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 38653 38586 38719 38589
rect 39297 38586 39363 38589
rect 38653 38584 39363 38586
rect 38653 38528 38658 38584
rect 38714 38528 39302 38584
rect 39358 38528 39363 38584
rect 38653 38526 39363 38528
rect 38653 38523 38719 38526
rect 39297 38523 39363 38526
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 27061 37226 27127 37229
rect 36169 37226 36235 37229
rect 27061 37224 36235 37226
rect 27061 37168 27066 37224
rect 27122 37168 36174 37224
rect 36230 37168 36235 37224
rect 27061 37166 36235 37168
rect 27061 37163 27127 37166
rect 36169 37163 36235 37166
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 27337 36274 27403 36277
rect 34329 36274 34395 36277
rect 27337 36272 34395 36274
rect 27337 36216 27342 36272
rect 27398 36216 34334 36272
rect 34390 36216 34395 36272
rect 27337 36214 34395 36216
rect 27337 36211 27403 36214
rect 34329 36211 34395 36214
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 45277 34778 45343 34781
rect 45537 34778 46337 34808
rect 45277 34776 46337 34778
rect 45277 34720 45282 34776
rect 45338 34720 46337 34776
rect 45277 34718 46337 34720
rect 45277 34715 45343 34718
rect 45537 34688 46337 34718
rect 33174 34580 33180 34644
rect 33244 34642 33250 34644
rect 33593 34642 33659 34645
rect 33244 34640 33659 34642
rect 33244 34584 33598 34640
rect 33654 34584 33659 34640
rect 33244 34582 33659 34584
rect 33244 34580 33250 34582
rect 33593 34579 33659 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 13721 34098 13787 34101
rect 24393 34098 24459 34101
rect 13721 34096 24459 34098
rect 13721 34040 13726 34096
rect 13782 34040 24398 34096
rect 24454 34040 24459 34096
rect 13721 34038 24459 34040
rect 13721 34035 13787 34038
rect 24393 34035 24459 34038
rect 10225 33962 10291 33965
rect 21173 33962 21239 33965
rect 10225 33960 21239 33962
rect 10225 33904 10230 33960
rect 10286 33904 21178 33960
rect 21234 33904 21239 33960
rect 10225 33902 21239 33904
rect 10225 33899 10291 33902
rect 21173 33899 21239 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 12157 33690 12223 33693
rect 17125 33690 17191 33693
rect 12157 33688 17191 33690
rect 12157 33632 12162 33688
rect 12218 33632 17130 33688
rect 17186 33632 17191 33688
rect 12157 33630 17191 33632
rect 12157 33627 12223 33630
rect 17125 33627 17191 33630
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 30097 33146 30163 33149
rect 33174 33146 33180 33148
rect 30097 33144 33180 33146
rect 30097 33088 30102 33144
rect 30158 33088 33180 33144
rect 30097 33086 33180 33088
rect 30097 33083 30163 33086
rect 33174 33084 33180 33086
rect 33244 33084 33250 33148
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 13169 31922 13235 31925
rect 18045 31922 18111 31925
rect 13169 31920 18111 31922
rect 13169 31864 13174 31920
rect 13230 31864 18050 31920
rect 18106 31864 18111 31920
rect 13169 31862 18111 31864
rect 13169 31859 13235 31862
rect 18045 31859 18111 31862
rect 12341 31786 12407 31789
rect 14273 31786 14339 31789
rect 12341 31784 14339 31786
rect 12341 31728 12346 31784
rect 12402 31728 14278 31784
rect 14334 31728 14339 31784
rect 12341 31726 14339 31728
rect 12341 31723 12407 31726
rect 14273 31723 14339 31726
rect 15469 31786 15535 31789
rect 19333 31786 19399 31789
rect 15469 31784 19399 31786
rect 15469 31728 15474 31784
rect 15530 31728 19338 31784
rect 19394 31728 19399 31784
rect 15469 31726 19399 31728
rect 15469 31723 15535 31726
rect 19333 31723 19399 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 12249 30698 12315 30701
rect 14825 30698 14891 30701
rect 12249 30696 14891 30698
rect 12249 30640 12254 30696
rect 12310 30640 14830 30696
rect 14886 30640 14891 30696
rect 12249 30638 14891 30640
rect 12249 30635 12315 30638
rect 14825 30635 14891 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 6545 30426 6611 30429
rect 11329 30426 11395 30429
rect 6545 30424 11395 30426
rect 6545 30368 6550 30424
rect 6606 30368 11334 30424
rect 11390 30368 11395 30424
rect 6545 30366 11395 30368
rect 6545 30363 6611 30366
rect 11329 30363 11395 30366
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 41781 29202 41847 29205
rect 43713 29202 43779 29205
rect 41781 29200 43779 29202
rect 41781 29144 41786 29200
rect 41842 29144 43718 29200
rect 43774 29144 43779 29200
rect 41781 29142 43779 29144
rect 41781 29139 41847 29142
rect 43713 29139 43779 29142
rect 13169 28930 13235 28933
rect 16573 28930 16639 28933
rect 13169 28928 16639 28930
rect 13169 28872 13174 28928
rect 13230 28872 16578 28928
rect 16634 28872 16639 28928
rect 13169 28870 16639 28872
rect 13169 28867 13235 28870
rect 16573 28867 16639 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 6821 28658 6887 28661
rect 12525 28658 12591 28661
rect 6821 28656 12591 28658
rect 6821 28600 6826 28656
rect 6882 28600 12530 28656
rect 12586 28600 12591 28656
rect 6821 28598 12591 28600
rect 6821 28595 6887 28598
rect 12525 28595 12591 28598
rect 5809 28522 5875 28525
rect 8937 28522 9003 28525
rect 5809 28520 9003 28522
rect 5809 28464 5814 28520
rect 5870 28464 8942 28520
rect 8998 28464 9003 28520
rect 5809 28462 9003 28464
rect 5809 28459 5875 28462
rect 8937 28459 9003 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 6453 28114 6519 28117
rect 13629 28114 13695 28117
rect 6453 28112 13695 28114
rect 6453 28056 6458 28112
rect 6514 28056 13634 28112
rect 13690 28056 13695 28112
rect 6453 28054 13695 28056
rect 6453 28051 6519 28054
rect 13629 28051 13695 28054
rect 0 27978 800 28008
rect 933 27978 999 27981
rect 0 27976 999 27978
rect 0 27920 938 27976
rect 994 27920 999 27976
rect 0 27918 999 27920
rect 0 27888 800 27918
rect 933 27915 999 27918
rect 8109 27978 8175 27981
rect 12433 27978 12499 27981
rect 8109 27976 12499 27978
rect 8109 27920 8114 27976
rect 8170 27920 12438 27976
rect 12494 27920 12499 27976
rect 8109 27918 12499 27920
rect 8109 27915 8175 27918
rect 12433 27915 12499 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 45277 25258 45343 25261
rect 45537 25258 46337 25288
rect 45277 25256 46337 25258
rect 45277 25200 45282 25256
rect 45338 25200 46337 25256
rect 45277 25198 46337 25200
rect 45277 25195 45343 25198
rect 45537 25168 46337 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 11237 23626 11303 23629
rect 15285 23626 15351 23629
rect 11237 23624 15351 23626
rect 11237 23568 11242 23624
rect 11298 23568 15290 23624
rect 15346 23568 15351 23624
rect 11237 23566 15351 23568
rect 11237 23563 11303 23566
rect 15285 23563 15351 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 31661 19954 31727 19957
rect 32305 19954 32371 19957
rect 31661 19952 32371 19954
rect 31661 19896 31666 19952
rect 31722 19896 32310 19952
rect 32366 19896 32371 19952
rect 31661 19894 32371 19896
rect 31661 19891 31727 19894
rect 32305 19891 32371 19894
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 33869 19410 33935 19413
rect 35801 19410 35867 19413
rect 33869 19408 35867 19410
rect 33869 19352 33874 19408
rect 33930 19352 35806 19408
rect 35862 19352 35867 19408
rect 33869 19350 35867 19352
rect 33869 19347 33935 19350
rect 35801 19347 35867 19350
rect 21173 19274 21239 19277
rect 21909 19274 21975 19277
rect 21173 19272 21975 19274
rect 21173 19216 21178 19272
rect 21234 19216 21914 19272
rect 21970 19216 21975 19272
rect 21173 19214 21975 19216
rect 21173 19211 21239 19214
rect 21909 19211 21975 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 22461 18052 22527 18053
rect 22461 18048 22508 18052
rect 22572 18050 22578 18052
rect 22461 17992 22466 18048
rect 22461 17988 22508 17992
rect 22572 17990 22618 18050
rect 22572 17988 22578 17990
rect 22461 17987 22527 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 22645 16692 22711 16693
rect 22645 16688 22692 16692
rect 22756 16690 22762 16692
rect 22645 16632 22650 16688
rect 22645 16628 22692 16632
rect 22756 16630 22802 16690
rect 22756 16628 22762 16630
rect 22645 16627 22711 16628
rect 44725 16418 44791 16421
rect 45537 16418 46337 16448
rect 44725 16416 46337 16418
rect 44725 16360 44730 16416
rect 44786 16360 46337 16416
rect 44725 16358 46337 16360
rect 44725 16355 44791 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 45537 16328 46337 16358
rect 19570 16287 19886 16288
rect 14273 15874 14339 15877
rect 14825 15874 14891 15877
rect 16113 15874 16179 15877
rect 14273 15872 19350 15874
rect 14273 15816 14278 15872
rect 14334 15816 14830 15872
rect 14886 15816 16118 15872
rect 16174 15816 19350 15872
rect 14273 15814 19350 15816
rect 14273 15811 14339 15814
rect 14825 15811 14891 15814
rect 16113 15811 16179 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 10685 15738 10751 15741
rect 18597 15738 18663 15741
rect 10685 15736 18663 15738
rect 10685 15680 10690 15736
rect 10746 15680 18602 15736
rect 18658 15680 18663 15736
rect 10685 15678 18663 15680
rect 19290 15738 19350 15814
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19793 15738 19859 15741
rect 20478 15738 20484 15740
rect 19290 15736 20484 15738
rect 19290 15680 19798 15736
rect 19854 15680 20484 15736
rect 19290 15678 20484 15680
rect 10685 15675 10751 15678
rect 18597 15675 18663 15678
rect 19793 15675 19859 15678
rect 20478 15676 20484 15678
rect 20548 15676 20554 15740
rect 22369 15738 22435 15741
rect 24117 15738 24183 15741
rect 22369 15736 24183 15738
rect 22369 15680 22374 15736
rect 22430 15680 24122 15736
rect 24178 15680 24183 15736
rect 22369 15678 24183 15680
rect 22369 15675 22435 15678
rect 24117 15675 24183 15678
rect 14549 15602 14615 15605
rect 21633 15602 21699 15605
rect 14549 15600 21699 15602
rect 14549 15544 14554 15600
rect 14610 15544 21638 15600
rect 21694 15544 21699 15600
rect 14549 15542 21699 15544
rect 14549 15539 14615 15542
rect 21633 15539 21699 15542
rect 11421 15466 11487 15469
rect 22093 15466 22159 15469
rect 11421 15464 22159 15466
rect 11421 15408 11426 15464
rect 11482 15408 22098 15464
rect 22154 15408 22159 15464
rect 11421 15406 22159 15408
rect 11421 15403 11487 15406
rect 22093 15403 22159 15406
rect 22737 15466 22803 15469
rect 23381 15466 23447 15469
rect 22737 15464 23447 15466
rect 22737 15408 22742 15464
rect 22798 15408 23386 15464
rect 23442 15408 23447 15464
rect 22737 15406 23447 15408
rect 22737 15403 22803 15406
rect 23381 15403 23447 15406
rect 17217 15332 17283 15333
rect 17166 15330 17172 15332
rect 17126 15270 17172 15330
rect 17236 15328 17283 15332
rect 17278 15272 17283 15328
rect 17166 15268 17172 15270
rect 17236 15268 17283 15272
rect 17217 15267 17283 15268
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 17677 15058 17743 15061
rect 19517 15058 19583 15061
rect 17677 15056 19583 15058
rect 17677 15000 17682 15056
rect 17738 15000 19522 15056
rect 19578 15000 19583 15056
rect 17677 14998 19583 15000
rect 17677 14995 17743 14998
rect 19517 14995 19583 14998
rect 11973 14922 12039 14925
rect 17585 14922 17651 14925
rect 11973 14920 17651 14922
rect 11973 14864 11978 14920
rect 12034 14864 17590 14920
rect 17646 14864 17651 14920
rect 11973 14862 17651 14864
rect 11973 14859 12039 14862
rect 17585 14859 17651 14862
rect 17033 14786 17099 14789
rect 17585 14786 17651 14789
rect 17033 14784 17651 14786
rect 17033 14728 17038 14784
rect 17094 14728 17590 14784
rect 17646 14728 17651 14784
rect 17033 14726 17651 14728
rect 17033 14723 17099 14726
rect 17585 14723 17651 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 15561 14650 15627 14653
rect 17953 14650 18019 14653
rect 15561 14648 18019 14650
rect 15561 14592 15566 14648
rect 15622 14592 17958 14648
rect 18014 14592 18019 14648
rect 15561 14590 18019 14592
rect 15561 14587 15627 14590
rect 17953 14587 18019 14590
rect 17125 14514 17191 14517
rect 19149 14514 19215 14517
rect 17125 14512 19215 14514
rect 17125 14456 17130 14512
rect 17186 14456 19154 14512
rect 19210 14456 19215 14512
rect 17125 14454 19215 14456
rect 17125 14451 17191 14454
rect 19149 14451 19215 14454
rect 10685 14378 10751 14381
rect 30373 14378 30439 14381
rect 10685 14376 30439 14378
rect 10685 14320 10690 14376
rect 10746 14320 30378 14376
rect 30434 14320 30439 14376
rect 10685 14318 30439 14320
rect 10685 14315 10751 14318
rect 30373 14315 30439 14318
rect 14733 14242 14799 14245
rect 18597 14242 18663 14245
rect 14733 14240 18663 14242
rect 14733 14184 14738 14240
rect 14794 14184 18602 14240
rect 18658 14184 18663 14240
rect 14733 14182 18663 14184
rect 14733 14179 14799 14182
rect 18597 14179 18663 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 14273 13970 14339 13973
rect 16665 13970 16731 13973
rect 14273 13968 16731 13970
rect 14273 13912 14278 13968
rect 14334 13912 16670 13968
rect 16726 13912 16731 13968
rect 14273 13910 16731 13912
rect 14273 13907 14339 13910
rect 16665 13907 16731 13910
rect 13261 13834 13327 13837
rect 13997 13834 14063 13837
rect 15837 13834 15903 13837
rect 13261 13832 15903 13834
rect 13261 13776 13266 13832
rect 13322 13776 14002 13832
rect 14058 13776 15842 13832
rect 15898 13776 15903 13832
rect 13261 13774 15903 13776
rect 13261 13771 13327 13774
rect 13997 13771 14063 13774
rect 15837 13771 15903 13774
rect 17309 13834 17375 13837
rect 22645 13834 22711 13837
rect 17309 13832 22711 13834
rect 17309 13776 17314 13832
rect 17370 13776 22650 13832
rect 22706 13776 22711 13832
rect 17309 13774 22711 13776
rect 17309 13771 17375 13774
rect 22645 13771 22711 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 22369 12882 22435 12885
rect 23054 12882 23060 12884
rect 22369 12880 23060 12882
rect 22369 12824 22374 12880
rect 22430 12824 23060 12880
rect 22369 12822 23060 12824
rect 22369 12819 22435 12822
rect 23054 12820 23060 12822
rect 23124 12820 23130 12884
rect 15193 12746 15259 12749
rect 15653 12746 15719 12749
rect 15193 12744 15719 12746
rect 15193 12688 15198 12744
rect 15254 12688 15658 12744
rect 15714 12688 15719 12744
rect 15193 12686 15719 12688
rect 15193 12683 15259 12686
rect 15653 12683 15719 12686
rect 19374 12684 19380 12748
rect 19444 12746 19450 12748
rect 19517 12746 19583 12749
rect 19444 12744 19583 12746
rect 19444 12688 19522 12744
rect 19578 12688 19583 12744
rect 19444 12686 19583 12688
rect 19444 12684 19450 12686
rect 19517 12683 19583 12686
rect 13997 12610 14063 12613
rect 15653 12610 15719 12613
rect 17677 12610 17743 12613
rect 13997 12608 17743 12610
rect 13997 12552 14002 12608
rect 14058 12552 15658 12608
rect 15714 12552 17682 12608
rect 17738 12552 17743 12608
rect 13997 12550 17743 12552
rect 13997 12547 14063 12550
rect 15653 12547 15719 12550
rect 17677 12547 17743 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 12382 12412 12388 12476
rect 12452 12474 12458 12476
rect 12525 12474 12591 12477
rect 12452 12472 12591 12474
rect 12452 12416 12530 12472
rect 12586 12416 12591 12472
rect 12452 12414 12591 12416
rect 12452 12412 12458 12414
rect 12525 12411 12591 12414
rect 20069 12338 20135 12341
rect 20069 12336 20178 12338
rect 20069 12280 20074 12336
rect 20130 12280 20178 12336
rect 20069 12275 20178 12280
rect 13721 12202 13787 12205
rect 19701 12202 19767 12205
rect 13721 12200 19767 12202
rect 13721 12144 13726 12200
rect 13782 12144 19706 12200
rect 19762 12144 19767 12200
rect 13721 12142 19767 12144
rect 13721 12139 13787 12142
rect 19701 12139 19767 12142
rect 20118 12069 20178 12275
rect 20478 12140 20484 12204
rect 20548 12202 20554 12204
rect 20621 12202 20687 12205
rect 20548 12200 20687 12202
rect 20548 12144 20626 12200
rect 20682 12144 20687 12200
rect 20548 12142 20687 12144
rect 20548 12140 20554 12142
rect 20621 12139 20687 12142
rect 12525 12066 12591 12069
rect 15193 12066 15259 12069
rect 12525 12064 15259 12066
rect 12525 12008 12530 12064
rect 12586 12008 15198 12064
rect 15254 12008 15259 12064
rect 12525 12006 15259 12008
rect 12525 12003 12591 12006
rect 15193 12003 15259 12006
rect 20069 12064 20178 12069
rect 20069 12008 20074 12064
rect 20130 12008 20178 12064
rect 20069 12006 20178 12008
rect 20069 12003 20135 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 15285 11794 15351 11797
rect 20989 11794 21055 11797
rect 15285 11792 21055 11794
rect 15285 11736 15290 11792
rect 15346 11736 20994 11792
rect 21050 11736 21055 11792
rect 15285 11734 21055 11736
rect 15285 11731 15351 11734
rect 20989 11731 21055 11734
rect 13486 11596 13492 11660
rect 13556 11658 13562 11660
rect 13813 11658 13879 11661
rect 16481 11658 16547 11661
rect 13556 11656 16547 11658
rect 13556 11600 13818 11656
rect 13874 11600 16486 11656
rect 16542 11600 16547 11656
rect 13556 11598 16547 11600
rect 13556 11596 13562 11598
rect 13813 11595 13879 11598
rect 16481 11595 16547 11598
rect 19701 11658 19767 11661
rect 20621 11658 20687 11661
rect 19701 11656 20687 11658
rect 19701 11600 19706 11656
rect 19762 11600 20626 11656
rect 20682 11600 20687 11656
rect 19701 11598 20687 11600
rect 19701 11595 19767 11598
rect 20621 11595 20687 11598
rect 11789 11522 11855 11525
rect 19609 11522 19675 11525
rect 11789 11520 19675 11522
rect 11789 11464 11794 11520
rect 11850 11464 19614 11520
rect 19670 11464 19675 11520
rect 11789 11462 19675 11464
rect 11789 11459 11855 11462
rect 19609 11459 19675 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 15009 11386 15075 11389
rect 18965 11386 19031 11389
rect 20437 11386 20503 11389
rect 15009 11384 20503 11386
rect 15009 11328 15014 11384
rect 15070 11328 18970 11384
rect 19026 11328 20442 11384
rect 20498 11328 20503 11384
rect 15009 11326 20503 11328
rect 15009 11323 15075 11326
rect 18965 11323 19031 11326
rect 20437 11323 20503 11326
rect 18321 11250 18387 11253
rect 30741 11250 30807 11253
rect 32121 11250 32187 11253
rect 18321 11248 19258 11250
rect 18321 11192 18326 11248
rect 18382 11192 19258 11248
rect 18321 11190 19258 11192
rect 18321 11187 18387 11190
rect 19198 11117 19258 11190
rect 30741 11248 32187 11250
rect 30741 11192 30746 11248
rect 30802 11192 32126 11248
rect 32182 11192 32187 11248
rect 30741 11190 32187 11192
rect 30741 11187 30807 11190
rect 32121 11187 32187 11190
rect 11513 11114 11579 11117
rect 17217 11114 17283 11117
rect 17953 11114 18019 11117
rect 18965 11114 19031 11117
rect 11513 11112 19031 11114
rect 11513 11056 11518 11112
rect 11574 11056 17222 11112
rect 17278 11056 17958 11112
rect 18014 11056 18970 11112
rect 19026 11056 19031 11112
rect 11513 11054 19031 11056
rect 11513 11051 11579 11054
rect 17217 11051 17283 11054
rect 17953 11051 18019 11054
rect 18965 11051 19031 11054
rect 19149 11112 19258 11117
rect 19149 11056 19154 11112
rect 19210 11056 19258 11112
rect 19149 11054 19258 11056
rect 31385 11114 31451 11117
rect 31845 11114 31911 11117
rect 31385 11112 31911 11114
rect 31385 11056 31390 11112
rect 31446 11056 31850 11112
rect 31906 11056 31911 11112
rect 31385 11054 31911 11056
rect 19149 11051 19215 11054
rect 31385 11051 31451 11054
rect 31845 11051 31911 11054
rect 15377 10978 15443 10981
rect 18597 10978 18663 10981
rect 22553 10980 22619 10981
rect 15377 10976 18663 10978
rect 15377 10920 15382 10976
rect 15438 10920 18602 10976
rect 18658 10920 18663 10976
rect 15377 10918 18663 10920
rect 15377 10915 15443 10918
rect 18597 10915 18663 10918
rect 22502 10916 22508 10980
rect 22572 10978 22619 10980
rect 22572 10976 22664 10978
rect 22614 10920 22664 10976
rect 22572 10918 22664 10920
rect 22572 10916 22619 10918
rect 22553 10915 22619 10916
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 13813 10842 13879 10845
rect 17309 10842 17375 10845
rect 13813 10840 17375 10842
rect 13813 10784 13818 10840
rect 13874 10784 17314 10840
rect 17370 10784 17375 10840
rect 13813 10782 17375 10784
rect 13813 10779 13879 10782
rect 17309 10779 17375 10782
rect 13261 10434 13327 10437
rect 17217 10434 17283 10437
rect 13261 10432 17283 10434
rect 13261 10376 13266 10432
rect 13322 10376 17222 10432
rect 17278 10376 17283 10432
rect 13261 10374 17283 10376
rect 13261 10371 13327 10374
rect 17217 10371 17283 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 11053 10298 11119 10301
rect 17033 10298 17099 10301
rect 11053 10296 17099 10298
rect 11053 10240 11058 10296
rect 11114 10240 17038 10296
rect 17094 10240 17099 10296
rect 11053 10238 17099 10240
rect 11053 10235 11119 10238
rect 17033 10235 17099 10238
rect 19425 10162 19491 10165
rect 19382 10160 19491 10162
rect 19382 10104 19430 10160
rect 19486 10104 19491 10160
rect 19382 10099 19491 10104
rect 14089 10026 14155 10029
rect 17861 10026 17927 10029
rect 14089 10024 17927 10026
rect 14089 9968 14094 10024
rect 14150 9968 17866 10024
rect 17922 9968 17927 10024
rect 14089 9966 17927 9968
rect 14089 9963 14155 9966
rect 17861 9963 17927 9966
rect 19382 9690 19442 10099
rect 20345 10026 20411 10029
rect 22553 10026 22619 10029
rect 20345 10024 22619 10026
rect 20345 9968 20350 10024
rect 20406 9968 22558 10024
rect 22614 9968 22619 10024
rect 20345 9966 22619 9968
rect 20345 9963 20411 9966
rect 22553 9963 22619 9966
rect 20345 9890 20411 9893
rect 20713 9890 20779 9893
rect 20345 9888 20779 9890
rect 20345 9832 20350 9888
rect 20406 9832 20718 9888
rect 20774 9832 20779 9888
rect 20345 9830 20779 9832
rect 20345 9827 20411 9830
rect 20713 9827 20779 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 29913 9754 29979 9757
rect 31661 9754 31727 9757
rect 29913 9752 31727 9754
rect 29913 9696 29918 9752
rect 29974 9696 31666 9752
rect 31722 9696 31727 9752
rect 29913 9694 31727 9696
rect 19517 9690 19583 9693
rect 29913 9691 29979 9694
rect 31661 9691 31727 9694
rect 19382 9688 19583 9690
rect 19382 9632 19522 9688
rect 19578 9632 19583 9688
rect 19382 9630 19583 9632
rect 19517 9627 19583 9630
rect 12709 9618 12775 9621
rect 15745 9618 15811 9621
rect 16481 9618 16547 9621
rect 17217 9620 17283 9621
rect 12709 9616 16547 9618
rect 12709 9560 12714 9616
rect 12770 9560 15750 9616
rect 15806 9560 16486 9616
rect 16542 9560 16547 9616
rect 12709 9558 16547 9560
rect 12709 9555 12775 9558
rect 15745 9555 15811 9558
rect 16481 9555 16547 9558
rect 17166 9556 17172 9620
rect 17236 9618 17283 9620
rect 22553 9618 22619 9621
rect 22686 9618 22692 9620
rect 17236 9616 17328 9618
rect 17278 9560 17328 9616
rect 17236 9558 17328 9560
rect 22553 9616 22692 9618
rect 22553 9560 22558 9616
rect 22614 9560 22692 9616
rect 22553 9558 22692 9560
rect 17236 9556 17283 9558
rect 17217 9555 17283 9556
rect 22553 9555 22619 9558
rect 22686 9556 22692 9558
rect 22756 9556 22762 9620
rect 38837 9618 38903 9621
rect 39113 9618 39179 9621
rect 38837 9616 39179 9618
rect 38837 9560 38842 9616
rect 38898 9560 39118 9616
rect 39174 9560 39179 9616
rect 38837 9558 39179 9560
rect 38837 9555 38903 9558
rect 39113 9555 39179 9558
rect 12341 9482 12407 9485
rect 12566 9482 12572 9484
rect 12341 9480 12572 9482
rect 12341 9424 12346 9480
rect 12402 9424 12572 9480
rect 12341 9422 12572 9424
rect 12341 9419 12407 9422
rect 12566 9420 12572 9422
rect 12636 9420 12642 9484
rect 12985 9482 13051 9485
rect 18413 9482 18479 9485
rect 19977 9482 20043 9485
rect 12985 9480 20043 9482
rect 12985 9424 12990 9480
rect 13046 9424 18418 9480
rect 18474 9424 19982 9480
rect 20038 9424 20043 9480
rect 12985 9422 20043 9424
rect 12985 9419 13051 9422
rect 18413 9419 18479 9422
rect 19977 9419 20043 9422
rect 19374 9284 19380 9348
rect 19444 9346 19450 9348
rect 19609 9346 19675 9349
rect 19444 9344 19675 9346
rect 19444 9288 19614 9344
rect 19670 9288 19675 9344
rect 19444 9286 19675 9288
rect 19444 9284 19450 9286
rect 19609 9283 19675 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 18597 9210 18663 9213
rect 19333 9210 19399 9213
rect 20069 9210 20135 9213
rect 18597 9208 20135 9210
rect 18597 9152 18602 9208
rect 18658 9152 19338 9208
rect 19394 9152 20074 9208
rect 20130 9152 20135 9208
rect 18597 9150 20135 9152
rect 18597 9147 18663 9150
rect 19333 9147 19399 9150
rect 20069 9147 20135 9150
rect 29545 9210 29611 9213
rect 30281 9210 30347 9213
rect 29545 9208 30347 9210
rect 29545 9152 29550 9208
rect 29606 9152 30286 9208
rect 30342 9152 30347 9208
rect 29545 9150 30347 9152
rect 29545 9147 29611 9150
rect 30281 9147 30347 9150
rect 30097 9074 30163 9077
rect 30833 9074 30899 9077
rect 30097 9072 30899 9074
rect 30097 9016 30102 9072
rect 30158 9016 30838 9072
rect 30894 9016 30899 9072
rect 30097 9014 30899 9016
rect 30097 9011 30163 9014
rect 30833 9011 30899 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 16665 8938 16731 8941
rect 17217 8938 17283 8941
rect 16665 8936 17283 8938
rect 16665 8880 16670 8936
rect 16726 8880 17222 8936
rect 17278 8880 17283 8936
rect 16665 8878 17283 8880
rect 16665 8875 16731 8878
rect 17217 8875 17283 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 20345 8258 20411 8261
rect 20478 8258 20484 8260
rect 20345 8256 20484 8258
rect 20345 8200 20350 8256
rect 20406 8200 20484 8256
rect 20345 8198 20484 8200
rect 20345 8195 20411 8198
rect 20478 8196 20484 8198
rect 20548 8196 20554 8260
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 23054 8060 23060 8124
rect 23124 8122 23130 8124
rect 23289 8122 23355 8125
rect 23124 8120 23355 8122
rect 23124 8064 23294 8120
rect 23350 8064 23355 8120
rect 23124 8062 23355 8064
rect 23124 8060 23130 8062
rect 23289 8059 23355 8062
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 13537 6900 13603 6901
rect 13486 6898 13492 6900
rect 13446 6838 13492 6898
rect 13556 6896 13603 6900
rect 13598 6840 13603 6896
rect 13486 6836 13492 6838
rect 13556 6836 13603 6840
rect 13537 6835 13603 6836
rect 16481 6898 16547 6901
rect 18321 6898 18387 6901
rect 16481 6896 18387 6898
rect 16481 6840 16486 6896
rect 16542 6840 18326 6896
rect 18382 6840 18387 6896
rect 16481 6838 18387 6840
rect 16481 6835 16547 6838
rect 18321 6835 18387 6838
rect 45277 6898 45343 6901
rect 45537 6898 46337 6928
rect 45277 6896 46337 6898
rect 45277 6840 45282 6896
rect 45338 6840 46337 6896
rect 45277 6838 46337 6840
rect 45277 6835 45343 6838
rect 45537 6808 46337 6838
rect 12341 6626 12407 6629
rect 17125 6626 17191 6629
rect 12341 6624 17191 6626
rect 12341 6568 12346 6624
rect 12402 6568 17130 6624
rect 17186 6568 17191 6624
rect 12341 6566 17191 6568
rect 12341 6563 12407 6566
rect 17125 6563 17191 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 15469 6354 15535 6357
rect 19057 6354 19123 6357
rect 15469 6352 19123 6354
rect 15469 6296 15474 6352
rect 15530 6296 19062 6352
rect 19118 6296 19123 6352
rect 15469 6294 19123 6296
rect 15469 6291 15535 6294
rect 19057 6291 19123 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 12525 5674 12591 5677
rect 17585 5674 17651 5677
rect 12525 5672 17651 5674
rect 12525 5616 12530 5672
rect 12586 5616 17590 5672
rect 17646 5616 17651 5672
rect 12525 5614 17651 5616
rect 12525 5611 12591 5614
rect 17585 5611 17651 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 36261 4314 36327 4317
rect 36629 4314 36695 4317
rect 36261 4312 36695 4314
rect 36261 4256 36266 4312
rect 36322 4256 36634 4312
rect 36690 4256 36695 4312
rect 36261 4254 36695 4256
rect 36261 4251 36327 4254
rect 36629 4251 36695 4254
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 30833 2954 30899 2957
rect 43897 2954 43963 2957
rect 30833 2952 43963 2954
rect 30833 2896 30838 2952
rect 30894 2896 43902 2952
rect 43958 2896 43963 2952
rect 30833 2894 43963 2896
rect 30833 2891 30899 2894
rect 43897 2891 43963 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 33180 34580 33244 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 33180 33084 33244 33148
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 22508 18048 22572 18052
rect 22508 17992 22522 18048
rect 22522 17992 22572 18048
rect 22508 17988 22572 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 22692 16688 22756 16692
rect 22692 16632 22706 16688
rect 22706 16632 22756 16688
rect 22692 16628 22756 16632
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 20484 15676 20548 15740
rect 17172 15328 17236 15332
rect 17172 15272 17222 15328
rect 17222 15272 17236 15328
rect 17172 15268 17236 15272
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 23060 12820 23124 12884
rect 19380 12684 19444 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 12388 12412 12452 12476
rect 20484 12140 20548 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 13492 11596 13556 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 22508 10976 22572 10980
rect 22508 10920 22558 10976
rect 22558 10920 22572 10976
rect 22508 10916 22572 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 17172 9616 17236 9620
rect 17172 9560 17222 9616
rect 17222 9560 17236 9616
rect 17172 9556 17236 9560
rect 22692 9556 22756 9620
rect 12572 9420 12636 9484
rect 19380 9284 19444 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 20484 8196 20548 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 23060 8060 23124 8124
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 13492 6896 13556 6900
rect 13492 6840 13542 6896
rect 13542 6840 13556 6896
rect 13492 6836 13556 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 46272 4528 46288
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 19568 45728 19888 46288
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 34928 46272 35248 46288
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 33179 34644 33245 34645
rect 33179 34580 33180 34644
rect 33244 34580 33245 34644
rect 33179 34579 33245 34580
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 33182 33149 33242 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 33179 33148 33245 33149
rect 33179 33084 33180 33148
rect 33244 33084 33245 33148
rect 33179 33083 33245 33084
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 22507 18052 22573 18053
rect 22507 17988 22508 18052
rect 22572 17988 22573 18052
rect 22507 17987 22573 17988
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 17171 15332 17237 15333
rect 17171 15268 17172 15332
rect 17236 15268 17237 15332
rect 17171 15267 17237 15268
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 12387 12476 12453 12477
rect 12387 12412 12388 12476
rect 12452 12450 12453 12476
rect 12452 12412 12634 12450
rect 12387 12411 12634 12412
rect 12390 12390 12634 12411
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 12574 9485 12634 12390
rect 13491 11660 13557 11661
rect 13491 11596 13492 11660
rect 13556 11596 13557 11660
rect 13491 11595 13557 11596
rect 12571 9484 12637 9485
rect 12571 9420 12572 9484
rect 12636 9420 12637 9484
rect 12571 9419 12637 9420
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 13494 6901 13554 11595
rect 17174 9621 17234 15267
rect 19568 15264 19888 16288
rect 20483 15740 20549 15741
rect 20483 15676 20484 15740
rect 20548 15676 20549 15740
rect 20483 15675 20549 15676
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19379 12748 19445 12749
rect 19379 12684 19380 12748
rect 19444 12684 19445 12748
rect 19379 12683 19445 12684
rect 17171 9620 17237 9621
rect 17171 9556 17172 9620
rect 17236 9556 17237 9620
rect 17171 9555 17237 9556
rect 19382 9349 19442 12683
rect 19568 12000 19888 13024
rect 20486 12205 20546 15675
rect 20483 12204 20549 12205
rect 20483 12140 20484 12204
rect 20548 12140 20549 12204
rect 20483 12139 20549 12140
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19379 9348 19445 9349
rect 19379 9284 19380 9348
rect 19444 9284 19445 9348
rect 19379 9283 19445 9284
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 20486 8261 20546 12139
rect 22510 10981 22570 17987
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 22691 16692 22757 16693
rect 22691 16628 22692 16692
rect 22756 16628 22757 16692
rect 22691 16627 22757 16628
rect 22507 10980 22573 10981
rect 22507 10916 22508 10980
rect 22572 10916 22573 10980
rect 22507 10915 22573 10916
rect 22694 9621 22754 16627
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 23059 12884 23125 12885
rect 23059 12820 23060 12884
rect 23124 12820 23125 12884
rect 23059 12819 23125 12820
rect 22691 9620 22757 9621
rect 22691 9556 22692 9620
rect 22756 9556 22757 9620
rect 22691 9555 22757 9556
rect 20483 8260 20549 8261
rect 20483 8196 20484 8260
rect 20548 8196 20549 8260
rect 20483 8195 20549 8196
rect 23062 8125 23122 12819
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 23059 8124 23125 8125
rect 23059 8060 23060 8124
rect 23124 8060 23125 8124
rect 23059 8059 23125 8060
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 13491 6900 13557 6901
rect 13491 6836 13492 6900
rect 13556 6836 13557 6900
rect 13491 6835 13557 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__and3_1  _1295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28152 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25852 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1297_
timestamp 1688980957
transform -1 0 23920 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1298_
timestamp 1688980957
transform -1 0 22908 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27692 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28428 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1302_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1303_
timestamp 1688980957
transform -1 0 24472 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1304_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23460 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1305_
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1688980957
transform -1 0 26864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1307_
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1308_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1309_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1310_
timestamp 1688980957
transform 1 0 10212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1688980957
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1312_
timestamp 1688980957
transform -1 0 31188 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1688980957
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1314_
timestamp 1688980957
transform 1 0 25576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1315_
timestamp 1688980957
transform -1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1316_
timestamp 1688980957
transform 1 0 15088 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1317_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1318_
timestamp 1688980957
transform 1 0 34960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1688980957
transform 1 0 35972 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1320_
timestamp 1688980957
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1688980957
transform -1 0 11040 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1322_
timestamp 1688980957
transform 1 0 32384 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1688980957
transform 1 0 32936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1324_
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1688980957
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1326_
timestamp 1688980957
transform -1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1327_
timestamp 1688980957
transform -1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1328_
timestamp 1688980957
transform 1 0 24840 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1688980957
transform -1 0 25484 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1330_
timestamp 1688980957
transform 1 0 6624 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1688980957
transform -1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1332_
timestamp 1688980957
transform 1 0 6624 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1688980957
transform 1 0 7268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1334_
timestamp 1688980957
transform 1 0 6808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1688980957
transform -1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1336_
timestamp 1688980957
transform -1 0 44436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 1688980957
transform -1 0 43608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1338_
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 1688980957
transform -1 0 8372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1340_
timestamp 1688980957
transform -1 0 44436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1688980957
transform -1 0 44068 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1342_
timestamp 1688980957
transform 1 0 43516 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1688980957
transform -1 0 44344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1688980957
transform -1 0 31556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1345_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1346_
timestamp 1688980957
transform 1 0 34776 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1347_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1348_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1688980957
transform 1 0 34500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1350_
timestamp 1688980957
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1351_
timestamp 1688980957
transform 1 0 34684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1352_
timestamp 1688980957
transform -1 0 36064 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1353_
timestamp 1688980957
transform -1 0 36340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1354_
timestamp 1688980957
transform -1 0 36800 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1357_
timestamp 1688980957
transform 1 0 37812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1358_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42320 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1359_
timestamp 1688980957
transform -1 0 42044 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1360_
timestamp 1688980957
transform 1 0 41308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1361_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _1362_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1363_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 39652 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1364_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1365_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1366_
timestamp 1688980957
transform 1 0 37996 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1367_
timestamp 1688980957
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1688980957
transform 1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1369_
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _1370_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39100 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1371_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1688980957
transform 1 0 40480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1688980957
transform 1 0 40756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1374_
timestamp 1688980957
transform -1 0 40756 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1375_
timestamp 1688980957
transform -1 0 40204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1376_
timestamp 1688980957
transform -1 0 41216 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1377_
timestamp 1688980957
transform 1 0 41216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1378_
timestamp 1688980957
transform -1 0 41308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1688980957
transform -1 0 42320 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1380_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42780 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1381_
timestamp 1688980957
transform 1 0 41860 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1688980957
transform 1 0 42780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42596 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1384_
timestamp 1688980957
transform -1 0 43056 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1385_
timestamp 1688980957
transform 1 0 43056 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1386_
timestamp 1688980957
transform 1 0 42412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1387_
timestamp 1688980957
transform -1 0 43056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1388_
timestamp 1688980957
transform -1 0 42872 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1389_
timestamp 1688980957
transform -1 0 42044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1390_
timestamp 1688980957
transform -1 0 42136 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1688980957
transform -1 0 41676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1392_
timestamp 1688980957
transform 1 0 41860 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1393_
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1394_
timestamp 1688980957
transform -1 0 42688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1395_
timestamp 1688980957
transform -1 0 40664 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1688980957
transform 1 0 40296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1397_
timestamp 1688980957
transform -1 0 39744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1398_
timestamp 1688980957
transform -1 0 36064 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1399_
timestamp 1688980957
transform -1 0 38088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1400_
timestamp 1688980957
transform -1 0 37720 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1401_
timestamp 1688980957
transform 1 0 38088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1403_
timestamp 1688980957
transform 1 0 36708 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1404_
timestamp 1688980957
transform -1 0 36892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1405_
timestamp 1688980957
transform 1 0 35696 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1406_
timestamp 1688980957
transform -1 0 37812 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1407_
timestamp 1688980957
transform -1 0 37168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1408_
timestamp 1688980957
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1688980957
transform 1 0 38916 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1410_
timestamp 1688980957
transform 1 0 38088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1411_
timestamp 1688980957
transform -1 0 40296 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1412_
timestamp 1688980957
transform -1 0 39192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1413_
timestamp 1688980957
transform 1 0 39100 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1414_
timestamp 1688980957
transform -1 0 36984 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1415_
timestamp 1688980957
transform -1 0 35236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1688980957
transform 1 0 43148 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1418_
timestamp 1688980957
transform -1 0 43700 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1419_
timestamp 1688980957
transform 1 0 42596 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1420_
timestamp 1688980957
transform -1 0 42320 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1421_
timestamp 1688980957
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1422_
timestamp 1688980957
transform -1 0 41308 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1423_
timestamp 1688980957
transform 1 0 41676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1424_
timestamp 1688980957
transform 1 0 42044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1425_
timestamp 1688980957
transform 1 0 39928 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1426_
timestamp 1688980957
transform -1 0 40296 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1427_
timestamp 1688980957
transform -1 0 40848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1428_
timestamp 1688980957
transform -1 0 39652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1429_
timestamp 1688980957
transform -1 0 39376 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1688980957
transform -1 0 39100 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1431_
timestamp 1688980957
transform -1 0 38640 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1432_
timestamp 1688980957
transform 1 0 37904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1433_
timestamp 1688980957
transform -1 0 38364 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1434_
timestamp 1688980957
transform 1 0 23000 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1435_
timestamp 1688980957
transform -1 0 23460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1436_
timestamp 1688980957
transform -1 0 23828 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1437_
timestamp 1688980957
transform 1 0 24472 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1438_
timestamp 1688980957
transform -1 0 35788 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1439_
timestamp 1688980957
transform -1 0 27692 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1440_
timestamp 1688980957
transform 1 0 28796 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1441_
timestamp 1688980957
transform -1 0 26864 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1442_
timestamp 1688980957
transform -1 0 26128 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1443_
timestamp 1688980957
transform -1 0 24012 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1688980957
transform 1 0 24012 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1445_
timestamp 1688980957
transform -1 0 22448 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1446_
timestamp 1688980957
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1447_
timestamp 1688980957
transform 1 0 22172 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 1688980957
transform 1 0 23736 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1449_
timestamp 1688980957
transform 1 0 21896 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1450_
timestamp 1688980957
transform 1 0 22264 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1451_
timestamp 1688980957
transform 1 0 22356 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1452_
timestamp 1688980957
transform 1 0 22172 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1688980957
transform -1 0 21712 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1454_
timestamp 1688980957
transform -1 0 18400 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1455_
timestamp 1688980957
transform 1 0 11684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1456_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13616 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1457_
timestamp 1688980957
transform -1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1458_
timestamp 1688980957
transform -1 0 21712 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1459_
timestamp 1688980957
transform 1 0 7728 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1460_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1461_
timestamp 1688980957
transform -1 0 15824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1462_
timestamp 1688980957
transform -1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1463_
timestamp 1688980957
transform -1 0 15916 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1464_
timestamp 1688980957
transform -1 0 15272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1465_
timestamp 1688980957
transform 1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1466_
timestamp 1688980957
transform 1 0 11868 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1467_
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1468_
timestamp 1688980957
transform -1 0 15824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1469_
timestamp 1688980957
transform -1 0 13984 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1470_
timestamp 1688980957
transform -1 0 14536 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1471_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1472_
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1473_
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1474_
timestamp 1688980957
transform -1 0 15088 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1475_
timestamp 1688980957
transform -1 0 17940 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1476_
timestamp 1688980957
transform -1 0 13984 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1477_
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1478_
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1479_
timestamp 1688980957
transform 1 0 9936 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1480_
timestamp 1688980957
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1481_
timestamp 1688980957
transform -1 0 13892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1483_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12788 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1484_
timestamp 1688980957
transform -1 0 16468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1485_
timestamp 1688980957
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1486_
timestamp 1688980957
transform 1 0 12880 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1487_
timestamp 1688980957
transform 1 0 12144 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1488_
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1489_
timestamp 1688980957
transform 1 0 12604 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1490_
timestamp 1688980957
transform -1 0 11868 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1491_
timestamp 1688980957
transform 1 0 12328 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1492_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1493_
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1494_
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1495_
timestamp 1688980957
transform -1 0 18952 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1496_
timestamp 1688980957
transform 1 0 17664 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1497_
timestamp 1688980957
transform 1 0 17940 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1688980957
transform -1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1499_
timestamp 1688980957
transform 1 0 16100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17020 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1501_
timestamp 1688980957
transform -1 0 16560 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1688980957
transform -1 0 16100 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1503_
timestamp 1688980957
transform -1 0 15548 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1504_
timestamp 1688980957
transform 1 0 15732 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1688980957
transform -1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1506_
timestamp 1688980957
transform 1 0 15272 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1688980957
transform -1 0 16560 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1508_
timestamp 1688980957
transform -1 0 14444 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1509_
timestamp 1688980957
transform -1 0 15272 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1510_
timestamp 1688980957
transform -1 0 15088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1511_
timestamp 1688980957
transform -1 0 14904 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1512_
timestamp 1688980957
transform -1 0 13248 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1513_
timestamp 1688980957
transform -1 0 12880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1514_
timestamp 1688980957
transform -1 0 9476 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1515_
timestamp 1688980957
transform -1 0 8832 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1516_
timestamp 1688980957
transform 1 0 9384 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1517_
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1688980957
transform -1 0 10304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1519_
timestamp 1688980957
transform -1 0 8740 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1520_
timestamp 1688980957
transform 1 0 7912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1521_
timestamp 1688980957
transform -1 0 9108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 1688980957
transform -1 0 6164 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1524_
timestamp 1688980957
transform 1 0 5704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1525_
timestamp 1688980957
transform -1 0 5704 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 1688980957
transform -1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 1688980957
transform 1 0 5612 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1688980957
transform 1 0 6532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1530_
timestamp 1688980957
transform -1 0 6808 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1688980957
transform -1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1532_
timestamp 1688980957
transform -1 0 5612 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1688980957
transform 1 0 4968 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1688980957
transform -1 0 6624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1535_
timestamp 1688980957
transform 1 0 5612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1536_
timestamp 1688980957
transform 1 0 6808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1537_
timestamp 1688980957
transform 1 0 7360 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1538_
timestamp 1688980957
transform 1 0 6900 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1688980957
transform -1 0 8096 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1540_
timestamp 1688980957
transform 1 0 6440 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1688980957
transform 1 0 6808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1543_
timestamp 1688980957
transform 1 0 9384 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1544_
timestamp 1688980957
transform 1 0 9016 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1688980957
transform 1 0 9660 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1546_
timestamp 1688980957
transform -1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1547_
timestamp 1688980957
transform 1 0 10396 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1548_
timestamp 1688980957
transform -1 0 11224 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1688980957
transform 1 0 12880 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1551_
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1552_
timestamp 1688980957
transform 1 0 12420 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1688980957
transform 1 0 12420 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1554_
timestamp 1688980957
transform 1 0 14168 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1555_
timestamp 1688980957
transform -1 0 14168 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1556_
timestamp 1688980957
transform -1 0 13616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1557_
timestamp 1688980957
transform -1 0 13984 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1558_
timestamp 1688980957
transform -1 0 14168 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1559_
timestamp 1688980957
transform 1 0 39192 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1560_
timestamp 1688980957
transform -1 0 39284 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1561_
timestamp 1688980957
transform -1 0 39192 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1688980957
transform -1 0 38180 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1688980957
transform -1 0 39560 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1564_
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1565_
timestamp 1688980957
transform -1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1566_
timestamp 1688980957
transform 1 0 7912 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1567_
timestamp 1688980957
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38548 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1569_
timestamp 1688980957
transform 1 0 37996 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1570_
timestamp 1688980957
transform -1 0 34316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1688980957
transform -1 0 33672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1572_
timestamp 1688980957
transform -1 0 35972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1574_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43700 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1575_
timestamp 1688980957
transform 1 0 10764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 1688980957
transform -1 0 12972 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1577_
timestamp 1688980957
transform 1 0 13616 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1578_
timestamp 1688980957
transform -1 0 13800 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1579_
timestamp 1688980957
transform 1 0 12880 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1580_
timestamp 1688980957
transform -1 0 14168 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1581_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12788 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1582_
timestamp 1688980957
transform 1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1583_
timestamp 1688980957
transform 1 0 9384 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1584_
timestamp 1688980957
transform -1 0 10028 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1585_
timestamp 1688980957
transform 1 0 7084 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1586_
timestamp 1688980957
transform 1 0 10028 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1688980957
transform 1 0 7728 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1589_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1590_
timestamp 1688980957
transform 1 0 10120 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1688980957
transform 1 0 8372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1592_
timestamp 1688980957
transform -1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1593_
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1594_
timestamp 1688980957
transform 1 0 10028 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1595_
timestamp 1688980957
transform 1 0 10304 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1596_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1597_
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 1688980957
transform 1 0 11224 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1599_
timestamp 1688980957
transform -1 0 18032 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1600_
timestamp 1688980957
transform -1 0 20240 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1601_
timestamp 1688980957
transform 1 0 17296 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1602_
timestamp 1688980957
transform -1 0 18768 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1688980957
transform -1 0 18952 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1604_
timestamp 1688980957
transform -1 0 18768 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1605_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18216 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1606_
timestamp 1688980957
transform -1 0 16560 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1688980957
transform 1 0 16744 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1688980957
transform 1 0 17572 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1609_
timestamp 1688980957
transform -1 0 17572 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1610_
timestamp 1688980957
transform -1 0 15272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1611_
timestamp 1688980957
transform -1 0 14996 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1612_
timestamp 1688980957
transform 1 0 15640 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1613_
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1614_
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1615_
timestamp 1688980957
transform -1 0 11408 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1616_
timestamp 1688980957
transform 1 0 14812 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1618_
timestamp 1688980957
transform 1 0 10580 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1619_
timestamp 1688980957
transform 1 0 9292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1620_
timestamp 1688980957
transform -1 0 9292 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1621_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10304 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1622_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1623_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1624_
timestamp 1688980957
transform -1 0 18400 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1625_
timestamp 1688980957
transform -1 0 17388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1626_
timestamp 1688980957
transform 1 0 17480 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1627_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1628_
timestamp 1688980957
transform 1 0 16376 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1629_
timestamp 1688980957
transform 1 0 15640 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1630_
timestamp 1688980957
transform 1 0 17020 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1631_
timestamp 1688980957
transform 1 0 41768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_4  _1632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 40848 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1633_
timestamp 1688980957
transform -1 0 41216 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1634_
timestamp 1688980957
transform 1 0 41124 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1635_
timestamp 1688980957
transform 1 0 38916 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1636_
timestamp 1688980957
transform 1 0 39376 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1637_
timestamp 1688980957
transform -1 0 39100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1638_
timestamp 1688980957
transform -1 0 40572 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39100 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1641_
timestamp 1688980957
transform -1 0 40940 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40572 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1643_
timestamp 1688980957
transform 1 0 43516 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1644_
timestamp 1688980957
transform -1 0 44896 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1645_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42504 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1646_
timestamp 1688980957
transform -1 0 44252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1647_
timestamp 1688980957
transform -1 0 44252 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1648_
timestamp 1688980957
transform -1 0 43056 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1649_
timestamp 1688980957
transform 1 0 43516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_2  _1650_
timestamp 1688980957
transform -1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1651_
timestamp 1688980957
transform 1 0 43700 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1652_
timestamp 1688980957
transform 1 0 44068 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1653_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1655_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42964 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1656_
timestamp 1688980957
transform 1 0 43424 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1657_
timestamp 1688980957
transform -1 0 43424 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1658_
timestamp 1688980957
transform 1 0 41216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1688980957
transform -1 0 42136 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1660_
timestamp 1688980957
transform -1 0 41400 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1661_
timestamp 1688980957
transform -1 0 41492 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1662_
timestamp 1688980957
transform -1 0 41032 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1663_
timestamp 1688980957
transform 1 0 40020 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1664_
timestamp 1688980957
transform -1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1688980957
transform 1 0 39652 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1666_
timestamp 1688980957
transform 1 0 39652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1667_
timestamp 1688980957
transform 1 0 39836 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1668_
timestamp 1688980957
transform 1 0 39284 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1669_
timestamp 1688980957
transform 1 0 39008 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1670_
timestamp 1688980957
transform -1 0 39744 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1671_
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1672_
timestamp 1688980957
transform -1 0 39652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1673_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36984 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1674_
timestamp 1688980957
transform 1 0 29808 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1675_
timestamp 1688980957
transform 1 0 31188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1676_
timestamp 1688980957
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1677_
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1678_
timestamp 1688980957
transform 1 0 31924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1679_
timestamp 1688980957
transform -1 0 39192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1688980957
transform -1 0 39744 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1681_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1682_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1683_
timestamp 1688980957
transform -1 0 24932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1688980957
transform 1 0 23552 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1688980957
transform -1 0 24288 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1687_
timestamp 1688980957
transform -1 0 24380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1688980957
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1688980957
transform 1 0 26128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1688980957
transform -1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1692_
timestamp 1688980957
transform 1 0 23460 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1693_
timestamp 1688980957
transform -1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1694_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1688980957
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1696_
timestamp 1688980957
transform -1 0 26864 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1697_
timestamp 1688980957
transform -1 0 26680 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1698_
timestamp 1688980957
transform 1 0 24840 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1688980957
transform -1 0 24932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1700_
timestamp 1688980957
transform 1 0 23552 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 1688980957
transform -1 0 23460 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1702_
timestamp 1688980957
transform -1 0 23828 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1688980957
transform 1 0 26680 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1688980957
transform -1 0 26864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1688980957
transform 1 0 24196 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1688980957
transform -1 0 24288 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1708_
timestamp 1688980957
transform -1 0 26680 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1688980957
transform 1 0 26680 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1688980957
transform -1 0 26864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1688980957
transform 1 0 27140 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1688980957
transform -1 0 27416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1688980957
transform 1 0 27140 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1688980957
transform -1 0 26956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1715_
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1716_
timestamp 1688980957
transform -1 0 26312 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1688980957
transform 1 0 28152 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1688980957
transform -1 0 27876 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1719_
timestamp 1688980957
transform -1 0 24104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1720_
timestamp 1688980957
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1721_
timestamp 1688980957
transform 1 0 23920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1722_
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1723_
timestamp 1688980957
transform -1 0 24380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1724_
timestamp 1688980957
transform -1 0 33580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1725_
timestamp 1688980957
transform 1 0 33580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1726_
timestamp 1688980957
transform -1 0 25852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1727_
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1728_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27048 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1729_
timestamp 1688980957
transform 1 0 27232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1730_
timestamp 1688980957
transform -1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1731_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1732_
timestamp 1688980957
transform 1 0 24472 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1733_
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1734_
timestamp 1688980957
transform -1 0 24288 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1735_
timestamp 1688980957
transform -1 0 24472 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1736_
timestamp 1688980957
transform -1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1738_
timestamp 1688980957
transform 1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1739_
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1740_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1741_
timestamp 1688980957
transform 1 0 24656 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1742_
timestamp 1688980957
transform 1 0 23828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1743_
timestamp 1688980957
transform 1 0 25852 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1744_
timestamp 1688980957
transform 1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1745_
timestamp 1688980957
transform -1 0 28152 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1746_
timestamp 1688980957
transform -1 0 28060 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1747_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1748_
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1749_
timestamp 1688980957
transform -1 0 29900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1750_
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1751_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1752_
timestamp 1688980957
transform -1 0 29440 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1753_
timestamp 1688980957
transform 1 0 30176 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1754_
timestamp 1688980957
transform 1 0 30820 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1755_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1756_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1688980957
transform 1 0 33948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1758_
timestamp 1688980957
transform -1 0 29348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1759_
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1760_
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1761_
timestamp 1688980957
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1762_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1763_
timestamp 1688980957
transform 1 0 35144 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1764_
timestamp 1688980957
transform -1 0 36248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1765_
timestamp 1688980957
transform -1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1766_
timestamp 1688980957
transform 1 0 36340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1767_
timestamp 1688980957
transform 1 0 29348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1768_
timestamp 1688980957
transform 1 0 28704 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1769_
timestamp 1688980957
transform 1 0 35512 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1770_
timestamp 1688980957
transform -1 0 35788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1771_
timestamp 1688980957
transform -1 0 36524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1772_
timestamp 1688980957
transform 1 0 35144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1773_
timestamp 1688980957
transform 1 0 36064 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1774_
timestamp 1688980957
transform -1 0 36064 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1775_
timestamp 1688980957
transform 1 0 35420 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1776_
timestamp 1688980957
transform 1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1777_
timestamp 1688980957
transform -1 0 35880 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1778_
timestamp 1688980957
transform 1 0 35972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1779_
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1780_
timestamp 1688980957
transform -1 0 30912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1781_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1782_
timestamp 1688980957
transform -1 0 37536 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1783_
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1784_
timestamp 1688980957
transform -1 0 37076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1785_
timestamp 1688980957
transform 1 0 36064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1688980957
transform -1 0 36064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1787_
timestamp 1688980957
transform -1 0 35972 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp 1688980957
transform -1 0 36156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1789_
timestamp 1688980957
transform 1 0 28612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1790_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1791_
timestamp 1688980957
transform 1 0 34224 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1792_
timestamp 1688980957
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1793_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1794_
timestamp 1688980957
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1795_
timestamp 1688980957
transform -1 0 33580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1796_
timestamp 1688980957
transform 1 0 27784 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1797_
timestamp 1688980957
transform 1 0 30084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1798_
timestamp 1688980957
transform 1 0 29440 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1799_
timestamp 1688980957
transform 1 0 31556 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 1688980957
transform 1 0 31004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1801_
timestamp 1688980957
transform 1 0 31004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1802_
timestamp 1688980957
transform -1 0 35880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1803_
timestamp 1688980957
transform -1 0 35788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1804_
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1805_
timestamp 1688980957
transform -1 0 34224 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1807_
timestamp 1688980957
transform -1 0 33304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1808_
timestamp 1688980957
transform -1 0 33028 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1809_
timestamp 1688980957
transform 1 0 31648 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp 1688980957
transform -1 0 31556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1811_
timestamp 1688980957
transform -1 0 29440 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1812_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1688980957
transform 1 0 31188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1814_
timestamp 1688980957
transform 1 0 31280 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1815_
timestamp 1688980957
transform 1 0 32292 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1816_
timestamp 1688980957
transform -1 0 32016 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1817_
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1818_
timestamp 1688980957
transform 1 0 32660 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1819_
timestamp 1688980957
transform -1 0 32292 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1820_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp 1688980957
transform 1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1822_
timestamp 1688980957
transform -1 0 30636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1823_
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1824_
timestamp 1688980957
transform 1 0 29624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1825_
timestamp 1688980957
transform 1 0 29624 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1826_
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1827_
timestamp 1688980957
transform -1 0 33304 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1828_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32844 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1829_
timestamp 1688980957
transform -1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1830_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32476 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1831_
timestamp 1688980957
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1832_
timestamp 1688980957
transform 1 0 28980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1833_
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1834_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1835_
timestamp 1688980957
transform 1 0 32476 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1836_
timestamp 1688980957
transform 1 0 33120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1837_
timestamp 1688980957
transform 1 0 33304 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1838_
timestamp 1688980957
transform -1 0 33580 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1839_
timestamp 1688980957
transform 1 0 33672 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1840_
timestamp 1688980957
transform -1 0 29992 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1841_
timestamp 1688980957
transform -1 0 29716 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1842_
timestamp 1688980957
transform 1 0 29072 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1843_
timestamp 1688980957
transform 1 0 34132 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1688980957
transform 1 0 34040 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1845_
timestamp 1688980957
transform 1 0 33672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_4  _1846_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32568 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _1847_
timestamp 1688980957
transform 1 0 35328 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1848_
timestamp 1688980957
transform -1 0 36524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1849_
timestamp 1688980957
transform 1 0 35512 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1850_
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1851_
timestamp 1688980957
transform 1 0 28428 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1852_
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1853_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35144 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1854_
timestamp 1688980957
transform 1 0 35604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1855_
timestamp 1688980957
transform 1 0 35880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1856_
timestamp 1688980957
transform -1 0 36248 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1857_
timestamp 1688980957
transform -1 0 34592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1858_
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1859_
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1860_
timestamp 1688980957
transform -1 0 35604 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1861_
timestamp 1688980957
transform 1 0 34868 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1862_
timestamp 1688980957
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1863_
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1864_
timestamp 1688980957
transform -1 0 30636 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1865_
timestamp 1688980957
transform 1 0 29716 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1688980957
transform 1 0 33120 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1867_
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1868_
timestamp 1688980957
transform 1 0 33580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1869_
timestamp 1688980957
transform 1 0 34776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1870_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1871_
timestamp 1688980957
transform -1 0 34408 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1872_
timestamp 1688980957
transform 1 0 32752 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1873_
timestamp 1688980957
transform 1 0 33396 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp 1688980957
transform -1 0 32384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1875_
timestamp 1688980957
transform -1 0 29992 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1876_
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1877_
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1878_
timestamp 1688980957
transform 1 0 32016 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1879_
timestamp 1688980957
transform 1 0 32568 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1880_
timestamp 1688980957
transform -1 0 34040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1881_
timestamp 1688980957
transform 1 0 33028 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1882_
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1883_
timestamp 1688980957
transform -1 0 34040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1884_
timestamp 1688980957
transform 1 0 30176 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1885_
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 1688980957
transform -1 0 32752 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1887_
timestamp 1688980957
transform 1 0 32752 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1888_
timestamp 1688980957
transform -1 0 32568 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1889_
timestamp 1688980957
transform 1 0 32200 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 1688980957
transform 1 0 33120 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1891_
timestamp 1688980957
transform 1 0 32476 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1892_
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1893_
timestamp 1688980957
transform -1 0 32568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1894_
timestamp 1688980957
transform 1 0 31188 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1895_
timestamp 1688980957
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1896_
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1897_
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1688980957
transform 1 0 30820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1899_
timestamp 1688980957
transform 1 0 30912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1900_
timestamp 1688980957
transform 1 0 31556 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1688980957
transform -1 0 33672 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1902_
timestamp 1688980957
transform -1 0 33396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1903_
timestamp 1688980957
transform 1 0 32660 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1904_
timestamp 1688980957
transform 1 0 33764 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1906_
timestamp 1688980957
transform -1 0 29808 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1907_
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1908_
timestamp 1688980957
transform -1 0 33580 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1909_
timestamp 1688980957
transform 1 0 33580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1910_
timestamp 1688980957
transform -1 0 33396 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1911_
timestamp 1688980957
transform 1 0 32108 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1912_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1913_
timestamp 1688980957
transform 1 0 32384 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1914_
timestamp 1688980957
transform -1 0 33120 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1915_
timestamp 1688980957
transform -1 0 24012 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1916_
timestamp 1688980957
transform 1 0 32568 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1917_
timestamp 1688980957
transform -1 0 33304 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1918_
timestamp 1688980957
transform 1 0 30176 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1919_
timestamp 1688980957
transform 1 0 29900 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1920_
timestamp 1688980957
transform 1 0 30084 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1921_
timestamp 1688980957
transform 1 0 32384 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1922_
timestamp 1688980957
transform -1 0 34040 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1923_
timestamp 1688980957
transform 1 0 33304 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1924_
timestamp 1688980957
transform 1 0 33948 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1925_
timestamp 1688980957
transform 1 0 28704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _1926_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30084 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1927_
timestamp 1688980957
transform 1 0 35144 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1928_
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1929_
timestamp 1688980957
transform 1 0 35420 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1930_
timestamp 1688980957
transform 1 0 33948 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1931_
timestamp 1688980957
transform -1 0 33304 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1932_
timestamp 1688980957
transform -1 0 32936 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1933_
timestamp 1688980957
transform -1 0 34132 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1934_
timestamp 1688980957
transform 1 0 34776 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1935_
timestamp 1688980957
transform 1 0 35604 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1936_
timestamp 1688980957
transform -1 0 34500 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1937_
timestamp 1688980957
transform -1 0 35788 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1938_
timestamp 1688980957
transform 1 0 34684 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1939_
timestamp 1688980957
transform 1 0 35236 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1940_
timestamp 1688980957
transform -1 0 34132 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1941_
timestamp 1688980957
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1942_
timestamp 1688980957
transform -1 0 34500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1943_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1944_
timestamp 1688980957
transform -1 0 33672 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1945_
timestamp 1688980957
transform -1 0 34684 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1946_
timestamp 1688980957
transform 1 0 33672 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1947_
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1948_
timestamp 1688980957
transform -1 0 34408 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1949_
timestamp 1688980957
transform -1 0 33672 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1950_
timestamp 1688980957
transform -1 0 34040 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1951_
timestamp 1688980957
transform 1 0 34040 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1952_
timestamp 1688980957
transform 1 0 34684 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1953_
timestamp 1688980957
transform 1 0 33672 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1954_
timestamp 1688980957
transform 1 0 32752 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1955_
timestamp 1688980957
transform -1 0 33120 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1956_
timestamp 1688980957
transform -1 0 32936 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1957_
timestamp 1688980957
transform 1 0 34224 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1958_
timestamp 1688980957
transform -1 0 32660 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1959_
timestamp 1688980957
transform 1 0 30728 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1960_
timestamp 1688980957
transform 1 0 30728 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1961_
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1962_
timestamp 1688980957
transform -1 0 31556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _1963_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30728 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1964_
timestamp 1688980957
transform 1 0 30360 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1965_
timestamp 1688980957
transform 1 0 30084 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1966_
timestamp 1688980957
transform -1 0 31924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1967_
timestamp 1688980957
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1968_
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1969_
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1970_
timestamp 1688980957
transform 1 0 31924 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1971_
timestamp 1688980957
transform 1 0 31188 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1972_
timestamp 1688980957
transform 1 0 30084 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1973_
timestamp 1688980957
transform -1 0 29992 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1974_
timestamp 1688980957
transform 1 0 29624 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1975_
timestamp 1688980957
transform 1 0 30452 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1976_
timestamp 1688980957
transform -1 0 30452 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1977_
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1978_
timestamp 1688980957
transform -1 0 30728 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1979_
timestamp 1688980957
transform -1 0 30452 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1980_
timestamp 1688980957
transform -1 0 30084 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1981_
timestamp 1688980957
transform -1 0 31372 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1982_
timestamp 1688980957
transform 1 0 30452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1983_
timestamp 1688980957
transform 1 0 28980 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1984_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30268 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1985_
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1986_
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1987_
timestamp 1688980957
transform 1 0 36616 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1988_
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1989_
timestamp 1688980957
transform -1 0 40480 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1990_
timestamp 1688980957
transform -1 0 39744 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1991_
timestamp 1688980957
transform 1 0 38824 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1992_
timestamp 1688980957
transform 1 0 38088 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1993_
timestamp 1688980957
transform -1 0 37076 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1994_
timestamp 1688980957
transform -1 0 25760 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1995_
timestamp 1688980957
transform -1 0 25300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1996_
timestamp 1688980957
transform -1 0 24380 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1997_
timestamp 1688980957
transform -1 0 23920 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1998_
timestamp 1688980957
transform -1 0 22540 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1999_
timestamp 1688980957
transform -1 0 23000 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2000_
timestamp 1688980957
transform -1 0 21436 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2001_
timestamp 1688980957
transform -1 0 20700 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2002_
timestamp 1688980957
transform 1 0 19504 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2003_
timestamp 1688980957
transform -1 0 18768 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2004_
timestamp 1688980957
transform 1 0 15824 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2005_
timestamp 1688980957
transform 1 0 10948 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2006_
timestamp 1688980957
transform 1 0 11500 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2007_
timestamp 1688980957
transform -1 0 10120 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2008_
timestamp 1688980957
transform -1 0 8924 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2009_
timestamp 1688980957
transform -1 0 8740 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2010_
timestamp 1688980957
transform -1 0 8372 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2011_
timestamp 1688980957
transform 1 0 18584 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2012_
timestamp 1688980957
transform -1 0 7636 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2013_
timestamp 1688980957
transform -1 0 4876 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2014_
timestamp 1688980957
transform -1 0 5704 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2015_
timestamp 1688980957
transform -1 0 4508 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2016_
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2017_
timestamp 1688980957
transform 1 0 4508 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2018_
timestamp 1688980957
transform 1 0 3864 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2019_
timestamp 1688980957
transform 1 0 4324 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2020_
timestamp 1688980957
transform 1 0 6072 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2021_
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2022_
timestamp 1688980957
transform 1 0 7360 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2023_
timestamp 1688980957
transform -1 0 8832 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2024_
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2025_
timestamp 1688980957
transform 1 0 11592 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2026_
timestamp 1688980957
transform 1 0 13432 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2027_
timestamp 1688980957
transform -1 0 14812 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2028_
timestamp 1688980957
transform -1 0 16008 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2029_
timestamp 1688980957
transform 1 0 15548 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2030_
timestamp 1688980957
transform 1 0 18124 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2031_
timestamp 1688980957
transform -1 0 19964 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2032_
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2033_
timestamp 1688980957
transform 1 0 24656 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2034_
timestamp 1688980957
transform -1 0 24288 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2035_
timestamp 1688980957
transform 1 0 26588 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2036_
timestamp 1688980957
transform -1 0 27508 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2037_
timestamp 1688980957
transform 1 0 26772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2038_
timestamp 1688980957
transform -1 0 28704 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1688980957
transform -1 0 27600 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2040_
timestamp 1688980957
transform 1 0 25852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1688980957
transform -1 0 27324 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2042_
timestamp 1688980957
transform -1 0 26864 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2043_
timestamp 1688980957
transform 1 0 27600 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2044_
timestamp 1688980957
transform -1 0 28152 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2045_
timestamp 1688980957
transform 1 0 26680 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 1688980957
transform -1 0 26496 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2047_
timestamp 1688980957
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2048_
timestamp 1688980957
transform 1 0 36064 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2049_
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2050_
timestamp 1688980957
transform 1 0 19872 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2051_
timestamp 1688980957
transform -1 0 42688 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2052_
timestamp 1688980957
transform -1 0 42780 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2053_
timestamp 1688980957
transform 1 0 42596 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2054_
timestamp 1688980957
transform -1 0 42780 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2055_
timestamp 1688980957
transform -1 0 43424 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2056_
timestamp 1688980957
transform 1 0 43424 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 1688980957
transform 1 0 40848 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2058_
timestamp 1688980957
transform -1 0 40388 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2059_
timestamp 1688980957
transform 1 0 39836 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2060_
timestamp 1688980957
transform -1 0 39744 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2061_
timestamp 1688980957
transform 1 0 38456 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2062_
timestamp 1688980957
transform 1 0 38180 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2063_
timestamp 1688980957
transform 1 0 37536 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2064_
timestamp 1688980957
transform -1 0 37536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2065_
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2066_
timestamp 1688980957
transform 1 0 36064 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2067_
timestamp 1688980957
transform 1 0 36156 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2068_
timestamp 1688980957
transform -1 0 38824 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2069_
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2070_
timestamp 1688980957
transform 1 0 37812 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2071_
timestamp 1688980957
transform 1 0 36616 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2072_
timestamp 1688980957
transform 1 0 41400 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2073_
timestamp 1688980957
transform -1 0 42228 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2074_
timestamp 1688980957
transform 1 0 41676 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2075_
timestamp 1688980957
transform 1 0 41032 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2076_
timestamp 1688980957
transform -1 0 39836 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2077_
timestamp 1688980957
transform 1 0 38180 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2078_
timestamp 1688980957
transform 1 0 37076 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2079_
timestamp 1688980957
transform -1 0 22264 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2080_
timestamp 1688980957
transform -1 0 21344 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2081_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 1688980957
transform -1 0 17480 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2084_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2085_
timestamp 1688980957
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2086_
timestamp 1688980957
transform 1 0 18032 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2087_
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2088_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2089_
timestamp 1688980957
transform 1 0 15732 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2090_
timestamp 1688980957
transform -1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2091_
timestamp 1688980957
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2092_
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2093_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2094_
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2095_
timestamp 1688980957
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2096_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2097_
timestamp 1688980957
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2098_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2099_
timestamp 1688980957
transform -1 0 12972 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2100_
timestamp 1688980957
transform 1 0 12788 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2101_
timestamp 1688980957
transform 1 0 15088 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2102_
timestamp 1688980957
transform -1 0 15088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2103_
timestamp 1688980957
transform 1 0 12236 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2104_
timestamp 1688980957
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2105_
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2106_
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2107_
timestamp 1688980957
transform 1 0 13340 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2108_
timestamp 1688980957
transform -1 0 12880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2109_
timestamp 1688980957
transform 1 0 21344 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2110_
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2111_
timestamp 1688980957
transform 1 0 22448 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2112_
timestamp 1688980957
transform 1 0 22080 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2113_
timestamp 1688980957
transform 1 0 24748 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2114_
timestamp 1688980957
transform -1 0 24748 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2115_
timestamp 1688980957
transform 1 0 25944 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2116_
timestamp 1688980957
transform 1 0 26312 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2117_
timestamp 1688980957
transform 1 0 22632 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2118_
timestamp 1688980957
transform -1 0 22632 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2119_
timestamp 1688980957
transform -1 0 24564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2120_
timestamp 1688980957
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2121_
timestamp 1688980957
transform 1 0 13524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2122_
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2123_
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2124_
timestamp 1688980957
transform -1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2125_
timestamp 1688980957
transform -1 0 13984 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2126_
timestamp 1688980957
transform 1 0 13156 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2127_
timestamp 1688980957
transform -1 0 14720 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2128_
timestamp 1688980957
transform -1 0 12144 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2129_
timestamp 1688980957
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2130_
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2131_
timestamp 1688980957
transform -1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2132_
timestamp 1688980957
transform 1 0 15088 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2133_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2134_
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2135_
timestamp 1688980957
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2136_
timestamp 1688980957
transform -1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2137_
timestamp 1688980957
transform -1 0 11960 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2138_
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2139_
timestamp 1688980957
transform 1 0 17664 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2140_
timestamp 1688980957
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2141_
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2142_
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2143_
timestamp 1688980957
transform -1 0 18124 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2144_
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2145_
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2146_
timestamp 1688980957
transform -1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2147_
timestamp 1688980957
transform -1 0 12052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2148_
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2149_
timestamp 1688980957
transform -1 0 12236 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2150_
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2151_
timestamp 1688980957
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2152_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2153_
timestamp 1688980957
transform 1 0 15088 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2154_
timestamp 1688980957
transform 1 0 12420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2155_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2156_
timestamp 1688980957
transform -1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2157_
timestamp 1688980957
transform -1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2158_
timestamp 1688980957
transform -1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2159_
timestamp 1688980957
transform -1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2160_
timestamp 1688980957
transform -1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2161_
timestamp 1688980957
transform -1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2162_
timestamp 1688980957
transform -1 0 19504 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2163_
timestamp 1688980957
transform -1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2164_
timestamp 1688980957
transform 1 0 19504 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _2165_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _2166_
timestamp 1688980957
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2167_
timestamp 1688980957
transform 1 0 32292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2168_
timestamp 1688980957
transform 1 0 31556 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2169_
timestamp 1688980957
transform 1 0 30820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2170_
timestamp 1688980957
transform -1 0 30360 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _2171_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30912 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__and2b_1  _2172_
timestamp 1688980957
transform 1 0 31924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2173_
timestamp 1688980957
transform 1 0 31280 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2174_
timestamp 1688980957
transform 1 0 29348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2175_
timestamp 1688980957
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2176_
timestamp 1688980957
transform 1 0 31096 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2177_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_2  _2178_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2179_
timestamp 1688980957
transform 1 0 31464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2180_
timestamp 1688980957
transform 1 0 31188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2181_
timestamp 1688980957
transform 1 0 32752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2182_
timestamp 1688980957
transform -1 0 31280 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2183_
timestamp 1688980957
transform -1 0 32568 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2184_
timestamp 1688980957
transform -1 0 30268 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2185_
timestamp 1688980957
transform -1 0 32108 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2186_
timestamp 1688980957
transform -1 0 32016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _2187_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30452 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_2  _2188_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _2189_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2190_
timestamp 1688980957
transform -1 0 29992 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2191_
timestamp 1688980957
transform -1 0 31280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2192_
timestamp 1688980957
transform -1 0 30360 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2193_
timestamp 1688980957
transform -1 0 30268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2194_
timestamp 1688980957
transform -1 0 32016 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31556 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2196_
timestamp 1688980957
transform -1 0 30728 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2197_
timestamp 1688980957
transform -1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2198_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2199_
timestamp 1688980957
transform 1 0 31280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2200_
timestamp 1688980957
transform -1 0 31004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2201_
timestamp 1688980957
transform -1 0 28796 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _2202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2203_
timestamp 1688980957
transform -1 0 29164 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2204_
timestamp 1688980957
transform -1 0 28428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2205_
timestamp 1688980957
transform -1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2206_
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _2207_
timestamp 1688980957
transform -1 0 28888 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2208_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2209_
timestamp 1688980957
transform -1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2210_
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2211_
timestamp 1688980957
transform 1 0 25576 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _2212_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2213_
timestamp 1688980957
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2214_
timestamp 1688980957
transform -1 0 30728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2215_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2216_
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2217_
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2218_
timestamp 1688980957
transform -1 0 31372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2219_
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2220_
timestamp 1688980957
transform 1 0 25576 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2221_
timestamp 1688980957
transform -1 0 29348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2222_
timestamp 1688980957
transform -1 0 32384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2223_
timestamp 1688980957
transform 1 0 31464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2224_
timestamp 1688980957
transform -1 0 29532 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _2225_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28520 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2226_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2227_
timestamp 1688980957
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2228_
timestamp 1688980957
transform -1 0 22724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2229_
timestamp 1688980957
transform 1 0 22632 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2230_
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2231_
timestamp 1688980957
transform -1 0 20700 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2232_
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2233_
timestamp 1688980957
transform -1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2234_
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _2235_
timestamp 1688980957
transform 1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2236_
timestamp 1688980957
transform -1 0 15088 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2237_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2238_
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2239_
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2240_
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2241_
timestamp 1688980957
transform -1 0 17664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2242_
timestamp 1688980957
transform 1 0 16928 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _2243_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2244_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2245_
timestamp 1688980957
transform -1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2246_
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2247_
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2248_
timestamp 1688980957
transform -1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2249_
timestamp 1688980957
transform -1 0 14536 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2250_
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2251_
timestamp 1688980957
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2252_
timestamp 1688980957
transform -1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2253_
timestamp 1688980957
transform 1 0 15916 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a31o_1  _2254_
timestamp 1688980957
transform 1 0 30452 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2255_
timestamp 1688980957
transform -1 0 29992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2256_
timestamp 1688980957
transform 1 0 26680 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2257_
timestamp 1688980957
transform 1 0 26312 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2258_
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2259_
timestamp 1688980957
transform 1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _2260_
timestamp 1688980957
transform -1 0 27600 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _2261_
timestamp 1688980957
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2262_
timestamp 1688980957
transform -1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2263_
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2264_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2265_
timestamp 1688980957
transform -1 0 21620 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2266_
timestamp 1688980957
transform -1 0 28612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2267_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2268_
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2269_
timestamp 1688980957
transform 1 0 25576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2270_
timestamp 1688980957
transform 1 0 24288 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2271_
timestamp 1688980957
transform -1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2272_
timestamp 1688980957
transform 1 0 16008 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2273_
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2274_
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2275_
timestamp 1688980957
transform 1 0 15456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2276_
timestamp 1688980957
transform -1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2277_
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2278_
timestamp 1688980957
transform -1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2279_
timestamp 1688980957
transform -1 0 14444 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2280_
timestamp 1688980957
transform 1 0 14904 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _2281_
timestamp 1688980957
transform -1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2282_
timestamp 1688980957
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2283_
timestamp 1688980957
transform -1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2284_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2285_
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2286_
timestamp 1688980957
transform -1 0 32292 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2287_
timestamp 1688980957
transform -1 0 29072 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2288_
timestamp 1688980957
transform 1 0 27508 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2289_
timestamp 1688980957
transform 1 0 25208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2290_
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2291_
timestamp 1688980957
transform 1 0 24656 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2292_
timestamp 1688980957
transform 1 0 23368 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2293_
timestamp 1688980957
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2294_
timestamp 1688980957
transform -1 0 16100 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2295_
timestamp 1688980957
transform 1 0 14536 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2296_
timestamp 1688980957
transform -1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _2297_
timestamp 1688980957
transform 1 0 16192 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2298_
timestamp 1688980957
transform 1 0 16100 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _2299_
timestamp 1688980957
transform -1 0 19136 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2300_
timestamp 1688980957
transform -1 0 17940 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _2301_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _2302_
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2303_
timestamp 1688980957
transform -1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2304_
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2305_
timestamp 1688980957
transform -1 0 20976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2306_
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _2307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2308_
timestamp 1688980957
transform -1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2309_
timestamp 1688980957
transform -1 0 19872 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2310_
timestamp 1688980957
transform -1 0 20792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2311_
timestamp 1688980957
transform -1 0 20976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2312_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2313_
timestamp 1688980957
transform -1 0 14536 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2314_
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2315_
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _2316_
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2317_
timestamp 1688980957
transform 1 0 20792 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2318_
timestamp 1688980957
transform -1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2319_
timestamp 1688980957
transform 1 0 28980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2320_
timestamp 1688980957
transform 1 0 28612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2321_
timestamp 1688980957
transform -1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2322_
timestamp 1688980957
transform 1 0 27048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2323_
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2324_
timestamp 1688980957
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2325_
timestamp 1688980957
transform -1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2326_
timestamp 1688980957
transform 1 0 21252 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2327_
timestamp 1688980957
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2328_
timestamp 1688980957
transform -1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2329_
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2330_
timestamp 1688980957
transform 1 0 15364 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2331_
timestamp 1688980957
transform 1 0 17940 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2332_
timestamp 1688980957
transform 1 0 16192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2333_
timestamp 1688980957
transform -1 0 17112 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2334_
timestamp 1688980957
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2335_
timestamp 1688980957
transform -1 0 17572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2336_
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2337_
timestamp 1688980957
transform -1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2338_
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2339_
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2340_
timestamp 1688980957
transform -1 0 17480 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2341_
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2342_
timestamp 1688980957
transform 1 0 26956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2343_
timestamp 1688980957
transform 1 0 24472 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2344_
timestamp 1688980957
transform 1 0 22448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2345_
timestamp 1688980957
transform -1 0 23000 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2346_
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2347_
timestamp 1688980957
transform -1 0 22356 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2348_
timestamp 1688980957
transform 1 0 31096 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2349_
timestamp 1688980957
transform 1 0 30084 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2350_
timestamp 1688980957
transform -1 0 29900 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2351_
timestamp 1688980957
transform 1 0 28060 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2352_
timestamp 1688980957
transform -1 0 27232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2353_
timestamp 1688980957
transform 1 0 26772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2354_
timestamp 1688980957
transform -1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2355_
timestamp 1688980957
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2356_
timestamp 1688980957
transform -1 0 13984 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2357_
timestamp 1688980957
transform 1 0 13524 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2358_
timestamp 1688980957
transform -1 0 19136 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2359_
timestamp 1688980957
transform -1 0 18492 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2360_
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _2361_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18584 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2362_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2363_
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _2364_
timestamp 1688980957
transform 1 0 16744 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2365_
timestamp 1688980957
transform -1 0 18032 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2366_
timestamp 1688980957
transform -1 0 18860 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _2367_
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2368_
timestamp 1688980957
transform -1 0 19872 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2369_
timestamp 1688980957
transform 1 0 12144 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _2370_
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2371_
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _2372_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2373_
timestamp 1688980957
transform -1 0 11408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2374_
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2375_
timestamp 1688980957
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2376_
timestamp 1688980957
transform -1 0 12972 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__a311o_1  _2377_
timestamp 1688980957
transform 1 0 30728 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2378_
timestamp 1688980957
transform -1 0 29348 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2379_
timestamp 1688980957
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2380_
timestamp 1688980957
transform 1 0 24748 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2381_
timestamp 1688980957
transform 1 0 23460 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2382_
timestamp 1688980957
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2383_
timestamp 1688980957
transform -1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2384_
timestamp 1688980957
transform 1 0 21988 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2385_
timestamp 1688980957
transform -1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2386_
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2387_
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2388_
timestamp 1688980957
transform -1 0 13248 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2389_
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2390_
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2391_
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2392_
timestamp 1688980957
transform -1 0 12236 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2393_
timestamp 1688980957
transform 1 0 12420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2394_
timestamp 1688980957
transform -1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2395_
timestamp 1688980957
transform -1 0 11960 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _2396_
timestamp 1688980957
transform -1 0 13340 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _2397_
timestamp 1688980957
transform -1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2398_
timestamp 1688980957
transform 1 0 28336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 1688980957
transform 1 0 27232 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2400_
timestamp 1688980957
transform 1 0 26128 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2401_
timestamp 1688980957
transform 1 0 22632 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2402_
timestamp 1688980957
transform -1 0 22632 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2404_
timestamp 1688980957
transform -1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2405_
timestamp 1688980957
transform 1 0 17848 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2406_
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2407_
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2408_
timestamp 1688980957
transform -1 0 19136 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2409_
timestamp 1688980957
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2410_
timestamp 1688980957
transform -1 0 18216 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2411_
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2412_
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2413_
timestamp 1688980957
transform -1 0 15916 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2414_
timestamp 1688980957
transform -1 0 16284 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2415_
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _2416_
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2417_
timestamp 1688980957
transform -1 0 20424 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2419_
timestamp 1688980957
transform -1 0 27232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2420_
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2421_
timestamp 1688980957
transform 1 0 22632 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _2422_
timestamp 1688980957
transform -1 0 20884 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2423_
timestamp 1688980957
transform 1 0 19872 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2424_
timestamp 1688980957
transform -1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2425_
timestamp 1688980957
transform 1 0 24748 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2426_
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2427_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2428_
timestamp 1688980957
transform 1 0 11960 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2429_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2430_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2431_
timestamp 1688980957
transform -1 0 11408 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2432_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2433_
timestamp 1688980957
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2434_
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2435_
timestamp 1688980957
transform -1 0 12052 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2436_
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2437_
timestamp 1688980957
transform 1 0 21896 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2438_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2439_
timestamp 1688980957
transform -1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2440_
timestamp 1688980957
transform -1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2441_
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2442_
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2443_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2444_
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2445_
timestamp 1688980957
transform -1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2446_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__or3_1  _2447_
timestamp 1688980957
transform -1 0 26864 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2448_
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2449_
timestamp 1688980957
transform -1 0 23920 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2450_
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2451_
timestamp 1688980957
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _2452_
timestamp 1688980957
transform 1 0 20516 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2453_
timestamp 1688980957
transform 1 0 19872 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2454_
timestamp 1688980957
transform -1 0 19504 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2455_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _2456_
timestamp 1688980957
transform 1 0 17204 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2457_
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2458_
timestamp 1688980957
transform 1 0 19504 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2459_
timestamp 1688980957
transform -1 0 20516 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2460_
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2461_
timestamp 1688980957
transform -1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2462_
timestamp 1688980957
transform -1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2463_
timestamp 1688980957
transform 1 0 23184 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2464_
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2465_
timestamp 1688980957
transform 1 0 19872 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2466_
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2467_
timestamp 1688980957
transform -1 0 19780 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2468_
timestamp 1688980957
transform 1 0 22724 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2469_
timestamp 1688980957
transform -1 0 20884 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _2470_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2471_
timestamp 1688980957
transform -1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2472_
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2473_
timestamp 1688980957
transform -1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2474_
timestamp 1688980957
transform -1 0 21160 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2475_
timestamp 1688980957
transform -1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2476_
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2477_
timestamp 1688980957
transform -1 0 21712 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2478_
timestamp 1688980957
transform -1 0 17664 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2479_
timestamp 1688980957
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2480_
timestamp 1688980957
transform -1 0 20608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2481_
timestamp 1688980957
transform -1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _2482_
timestamp 1688980957
transform -1 0 20056 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2483_
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2484_
timestamp 1688980957
transform -1 0 24288 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2485_
timestamp 1688980957
transform -1 0 24288 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2486_
timestamp 1688980957
transform 1 0 23644 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2487_
timestamp 1688980957
transform 1 0 19596 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2488_
timestamp 1688980957
transform -1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2489_
timestamp 1688980957
transform -1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2490_
timestamp 1688980957
transform -1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2491_
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2492_
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2493_
timestamp 1688980957
transform -1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2494_
timestamp 1688980957
transform -1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2495_
timestamp 1688980957
transform -1 0 20608 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2496_
timestamp 1688980957
transform -1 0 21620 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2497_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2498_
timestamp 1688980957
transform 1 0 24564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2499_
timestamp 1688980957
transform -1 0 25392 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2500_
timestamp 1688980957
transform 1 0 25392 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _2501_
timestamp 1688980957
transform -1 0 23552 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2502_
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2503_
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 22356 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2505_
timestamp 1688980957
transform -1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 1688980957
transform 1 0 16744 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2507_
timestamp 1688980957
transform 1 0 16100 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 1688980957
transform 1 0 17940 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2509_
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2511_
timestamp 1688980957
transform 1 0 17204 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2512_
timestamp 1688980957
transform -1 0 15824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2513_
timestamp 1688980957
transform 1 0 15272 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2514_
timestamp 1688980957
transform 1 0 14996 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2515_
timestamp 1688980957
transform 1 0 15640 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2516_
timestamp 1688980957
transform 1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2518_
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2519_
timestamp 1688980957
transform 1 0 13984 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2520_
timestamp 1688980957
transform -1 0 12144 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2521_
timestamp 1688980957
transform 1 0 10488 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2522_
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2524_
timestamp 1688980957
transform 1 0 10212 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2525_
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2526_
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2527_
timestamp 1688980957
transform 1 0 9384 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2528_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2529_
timestamp 1688980957
transform 1 0 10304 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2530_
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2532_
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2533_
timestamp 1688980957
transform 1 0 23276 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2534_
timestamp 1688980957
transform 1 0 19688 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2535_
timestamp 1688980957
transform -1 0 19136 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2536_
timestamp 1688980957
transform 1 0 20608 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2537_
timestamp 1688980957
transform 1 0 20148 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 1688980957
transform -1 0 22908 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 1688980957
transform 1 0 24656 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2541_
timestamp 1688980957
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 1688980957
transform 1 0 23644 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2543_
timestamp 1688980957
transform 1 0 21988 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2544_
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2545_
timestamp 1688980957
transform -1 0 23920 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2546_
timestamp 1688980957
transform 1 0 21988 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2547_
timestamp 1688980957
transform -1 0 21712 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2548_
timestamp 1688980957
transform 1 0 20056 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2549_
timestamp 1688980957
transform -1 0 19504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2550_
timestamp 1688980957
transform 1 0 17204 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2551_
timestamp 1688980957
transform 1 0 17756 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2552_
timestamp 1688980957
transform 1 0 17664 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2553_
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2554_
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2555_
timestamp 1688980957
transform -1 0 13432 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2556_
timestamp 1688980957
transform 1 0 14168 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 1688980957
transform 1 0 8188 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2558_
timestamp 1688980957
transform -1 0 7360 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2559_
timestamp 1688980957
transform 1 0 7544 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2560_
timestamp 1688980957
transform 1 0 7360 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 1688980957
transform 1 0 2668 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2562_
timestamp 1688980957
transform 1 0 2116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2563_
timestamp 1688980957
transform 1 0 2024 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2564_
timestamp 1688980957
transform 1 0 1748 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2565_
timestamp 1688980957
transform -1 0 5612 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2566_
timestamp 1688980957
transform 1 0 5612 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 1688980957
transform 1 0 2576 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 1688980957
transform 1 0 2116 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2569_
timestamp 1688980957
transform 1 0 5336 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2570_
timestamp 1688980957
transform 1 0 5060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2571_
timestamp 1688980957
transform 1 0 20240 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2572_
timestamp 1688980957
transform 1 0 9752 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2573_
timestamp 1688980957
transform 1 0 8556 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2574_
timestamp 1688980957
transform -1 0 11408 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2575_
timestamp 1688980957
transform 1 0 12420 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2576_
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2577_
timestamp 1688980957
transform 1 0 13616 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2579_
timestamp 1688980957
transform 1 0 15732 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2580_
timestamp 1688980957
transform 1 0 19228 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2581_
timestamp 1688980957
transform -1 0 18308 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2582_
timestamp 1688980957
transform -1 0 22264 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2583_
timestamp 1688980957
transform 1 0 23000 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2584_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2585_
timestamp 1688980957
transform -1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2586_
timestamp 1688980957
transform 1 0 19504 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2587_
timestamp 1688980957
transform -1 0 19504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2588_
timestamp 1688980957
transform -1 0 18768 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2589_
timestamp 1688980957
transform 1 0 18584 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2590_
timestamp 1688980957
transform 1 0 15548 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2591_
timestamp 1688980957
transform -1 0 15364 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2592_
timestamp 1688980957
transform -1 0 13524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2593_
timestamp 1688980957
transform 1 0 11776 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2594_
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2595_
timestamp 1688980957
transform 1 0 8648 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2596_
timestamp 1688980957
transform 1 0 7544 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2597_
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2598_
timestamp 1688980957
transform 1 0 7176 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2599_
timestamp 1688980957
transform 1 0 3864 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2600_
timestamp 1688980957
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2601_
timestamp 1688980957
transform -1 0 3680 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2602_
timestamp 1688980957
transform 1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2603_
timestamp 1688980957
transform 1 0 3956 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2604_
timestamp 1688980957
transform -1 0 3956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2605_
timestamp 1688980957
transform 1 0 3864 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2606_
timestamp 1688980957
transform -1 0 3036 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2607_
timestamp 1688980957
transform -1 0 7176 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2608_
timestamp 1688980957
transform 1 0 6900 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2609_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2610_
timestamp 1688980957
transform 1 0 8280 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2611_
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2612_
timestamp 1688980957
transform 1 0 10488 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2613_
timestamp 1688980957
transform 1 0 13064 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2614_
timestamp 1688980957
transform 1 0 13156 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2615_
timestamp 1688980957
transform 1 0 15364 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2616_
timestamp 1688980957
transform -1 0 15272 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2617_
timestamp 1688980957
transform -1 0 19136 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2618_
timestamp 1688980957
transform 1 0 18584 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2619_
timestamp 1688980957
transform 1 0 24288 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2620_
timestamp 1688980957
transform -1 0 24288 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2621_
timestamp 1688980957
transform 1 0 21620 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2622_
timestamp 1688980957
transform 1 0 21252 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2623_
timestamp 1688980957
transform 1 0 19872 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2624_
timestamp 1688980957
transform 1 0 19596 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2625_
timestamp 1688980957
transform 1 0 17848 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2626_
timestamp 1688980957
transform 1 0 17848 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2627_
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2628_
timestamp 1688980957
transform -1 0 16560 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2629_
timestamp 1688980957
transform -1 0 15456 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2630_
timestamp 1688980957
transform -1 0 13524 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2631_
timestamp 1688980957
transform -1 0 13984 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2632_
timestamp 1688980957
transform 1 0 9568 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2633_
timestamp 1688980957
transform -1 0 9476 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2634_
timestamp 1688980957
transform 1 0 8740 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2635_
timestamp 1688980957
transform -1 0 8832 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2636_
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2637_
timestamp 1688980957
transform 1 0 3312 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2638_
timestamp 1688980957
transform 1 0 2392 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2639_
timestamp 1688980957
transform 1 0 1932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2640_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2641_
timestamp 1688980957
transform 1 0 5888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2642_
timestamp 1688980957
transform 1 0 2392 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2643_
timestamp 1688980957
transform 1 0 1932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2644_
timestamp 1688980957
transform 1 0 5428 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2645_
timestamp 1688980957
transform 1 0 5152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2646_
timestamp 1688980957
transform 1 0 9108 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2647_
timestamp 1688980957
transform -1 0 9108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2648_
timestamp 1688980957
transform 1 0 11592 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2649_
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2650_
timestamp 1688980957
transform -1 0 14904 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2651_
timestamp 1688980957
transform 1 0 14904 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2652_
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2653_
timestamp 1688980957
transform -1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2654_
timestamp 1688980957
transform 1 0 18308 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2655_
timestamp 1688980957
transform 1 0 18216 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2656_
timestamp 1688980957
transform 1 0 17296 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2657_
timestamp 1688980957
transform 1 0 17204 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2658_
timestamp 1688980957
transform -1 0 18768 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _2659_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2660_
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2661_
timestamp 1688980957
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2662_
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2663_
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2664_
timestamp 1688980957
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2665_
timestamp 1688980957
transform 1 0 12604 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2666_
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2667_
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2668_
timestamp 1688980957
transform 1 0 11960 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2669_
timestamp 1688980957
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2670_
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2671_
timestamp 1688980957
transform -1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2672_
timestamp 1688980957
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2673_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2674_
timestamp 1688980957
transform -1 0 20976 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2675_
timestamp 1688980957
transform -1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2676_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2677_
timestamp 1688980957
transform -1 0 29992 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2678_
timestamp 1688980957
transform 1 0 26220 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2679_
timestamp 1688980957
transform 1 0 24380 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2680_
timestamp 1688980957
transform 1 0 21804 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2681_
timestamp 1688980957
transform 1 0 21344 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 1688980957
transform 1 0 21252 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 21160 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 38180 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2685_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2686_
timestamp 1688980957
transform 1 0 24932 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2690_
timestamp 1688980957
transform 1 0 25944 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2691_
timestamp 1688980957
transform 1 0 23828 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform 1 0 24932 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform -1 0 24196 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2696_
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2697_
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2698_
timestamp 1688980957
transform 1 0 26680 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 1688980957
transform 1 0 26956 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 26312 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2703_
timestamp 1688980957
transform 1 0 27876 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2704_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2705_
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2706_
timestamp 1688980957
transform -1 0 3496 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 1688980957
transform 1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2708_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2710_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2711_
timestamp 1688980957
transform -1 0 8280 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2712_
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2714_
timestamp 1688980957
transform -1 0 10764 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2715_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2716_
timestamp 1688980957
transform -1 0 8280 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2717_
timestamp 1688980957
transform 1 0 7636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2718_
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2719_
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2720_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _2721_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2722_
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2723_
timestamp 1688980957
transform 1 0 30452 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 1688980957
transform 1 0 32384 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 1688980957
transform 1 0 32936 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 1688980957
transform 1 0 32752 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 1688980957
transform 1 0 35328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 1688980957
transform 1 0 35420 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 1688980957
transform -1 0 39376 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 1688980957
transform -1 0 40480 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 1688980957
transform 1 0 39284 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 1688980957
transform 1 0 40296 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 1688980957
transform 1 0 43056 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 1688980957
transform 1 0 43056 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2736_
timestamp 1688980957
transform -1 0 43516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2737_
timestamp 1688980957
transform -1 0 43700 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2738_
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2739_
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2740_
timestamp 1688980957
transform -1 0 39100 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2741_
timestamp 1688980957
transform 1 0 34776 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2742_
timestamp 1688980957
transform 1 0 37260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2743_
timestamp 1688980957
transform 1 0 36340 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2744_
timestamp 1688980957
transform -1 0 40204 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2745_
timestamp 1688980957
transform -1 0 41676 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2746_
timestamp 1688980957
transform 1 0 36800 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2747_
timestamp 1688980957
transform 1 0 37536 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2748_
timestamp 1688980957
transform -1 0 34960 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2749_
timestamp 1688980957
transform -1 0 34132 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2750_
timestamp 1688980957
transform -1 0 35420 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2751_
timestamp 1688980957
transform -1 0 34132 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2752_
timestamp 1688980957
transform -1 0 36800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2753_
timestamp 1688980957
transform 1 0 28520 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2754_
timestamp 1688980957
transform -1 0 32016 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2755_
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2756_
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 1688980957
transform -1 0 37812 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 1688980957
transform 1 0 29348 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2759_
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2760_
timestamp 1688980957
transform -1 0 30636 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2761_
timestamp 1688980957
transform 1 0 11592 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2762_
timestamp 1688980957
transform 1 0 27600 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2763_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2764_
timestamp 1688980957
transform 1 0 9200 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2765_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2766_
timestamp 1688980957
transform -1 0 37904 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2767_
timestamp 1688980957
transform 1 0 32844 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2768_
timestamp 1688980957
transform -1 0 40756 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2769_
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2770_
timestamp 1688980957
transform 1 0 26496 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2771_
timestamp 1688980957
transform 1 0 29532 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2772_
timestamp 1688980957
transform 1 0 27600 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2773_
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2774_
timestamp 1688980957
transform 1 0 34960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2775_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2776_
timestamp 1688980957
transform 1 0 32292 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 1688980957
transform 1 0 25944 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 1688980957
transform -1 0 44160 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2785_
timestamp 1688980957
transform 1 0 37812 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2786_
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2787_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2788_
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2789_
timestamp 1688980957
transform 1 0 35972 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2790_
timestamp 1688980957
transform 1 0 35512 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2791_
timestamp 1688980957
transform -1 0 37904 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2792_
timestamp 1688980957
transform -1 0 34592 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 1688980957
transform -1 0 32752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 1688980957
transform -1 0 34500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 1688980957
transform 1 0 30544 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2796_
timestamp 1688980957
transform -1 0 36616 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2797_
timestamp 1688980957
transform -1 0 38548 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2798_
timestamp 1688980957
transform 1 0 35328 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 1688980957
transform -1 0 32660 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 1688980957
transform 1 0 34132 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 1688980957
transform 1 0 29992 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 1688980957
transform -1 0 35604 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 1688980957
transform 1 0 30728 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 1688980957
transform -1 0 36524 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 1688980957
transform -1 0 38088 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 1688980957
transform -1 0 37720 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 1688980957
transform 1 0 33948 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2808_
timestamp 1688980957
transform -1 0 33948 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 1688980957
transform 1 0 30268 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2810_
timestamp 1688980957
transform 1 0 28796 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 1688980957
transform 1 0 28152 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2812_
timestamp 1688980957
transform 1 0 27416 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2813_
timestamp 1688980957
transform 1 0 35512 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2814_
timestamp 1688980957
transform 1 0 37260 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2815_
timestamp 1688980957
transform 1 0 39928 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2816_
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2817_
timestamp 1688980957
transform 1 0 38824 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2818_
timestamp 1688980957
transform -1 0 40112 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2819_
timestamp 1688980957
transform -1 0 39560 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2820_
timestamp 1688980957
transform -1 0 37260 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2821_
timestamp 1688980957
transform 1 0 25300 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2822_
timestamp 1688980957
transform 1 0 22448 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2823_
timestamp 1688980957
transform -1 0 22356 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2824_
timestamp 1688980957
transform -1 0 20608 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2825_
timestamp 1688980957
transform -1 0 18308 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2826_
timestamp 1688980957
transform -1 0 11132 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2827_
timestamp 1688980957
transform 1 0 6440 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2828_
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2829_
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2830_
timestamp 1688980957
transform 1 0 1564 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2831_
timestamp 1688980957
transform 1 0 1840 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2832_
timestamp 1688980957
transform -1 0 6164 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2833_
timestamp 1688980957
transform -1 0 7452 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2834_
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2835_
timestamp 1688980957
transform -1 0 12696 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2836_
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2837_
timestamp 1688980957
transform -1 0 18124 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2838_
timestamp 1688980957
transform 1 0 19136 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2839_
timestamp 1688980957
transform -1 0 28244 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2840_
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2841_
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2842_
timestamp 1688980957
transform 1 0 24380 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2843_
timestamp 1688980957
transform 1 0 26496 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2844_
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2845_
timestamp 1688980957
transform 1 0 35604 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2846_
timestamp 1688980957
transform 1 0 42780 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2847_
timestamp 1688980957
transform 1 0 42780 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2848_
timestamp 1688980957
transform 1 0 42688 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2849_
timestamp 1688980957
transform 1 0 40388 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2850_
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2851_
timestamp 1688980957
transform 1 0 37720 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2852_
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2853_
timestamp 1688980957
transform -1 0 37076 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2854_
timestamp 1688980957
transform 1 0 40664 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2855_
timestamp 1688980957
transform 1 0 42412 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2856_
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2857_
timestamp 1688980957
transform 1 0 39928 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2858_
timestamp 1688980957
transform 1 0 38824 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2859_
timestamp 1688980957
transform 1 0 37628 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2860_
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2861_
timestamp 1688980957
transform -1 0 32292 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2862_
timestamp 1688980957
transform 1 0 27140 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2863_
timestamp 1688980957
transform -1 0 44620 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2864_
timestamp 1688980957
transform 1 0 42964 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2865_
timestamp 1688980957
transform -1 0 44712 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2866_
timestamp 1688980957
transform 1 0 41032 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2867_
timestamp 1688980957
transform 1 0 40204 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2868_
timestamp 1688980957
transform 1 0 38732 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2869_
timestamp 1688980957
transform 1 0 37352 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2870_
timestamp 1688980957
transform 1 0 37444 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _2871_
timestamp 1688980957
transform 1 0 17848 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2872_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2873_
timestamp 1688980957
transform 1 0 16652 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2874_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2875_
timestamp 1688980957
transform 1 0 14260 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2876_
timestamp 1688980957
transform 1 0 12052 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2877_
timestamp 1688980957
transform -1 0 11408 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2878_
timestamp 1688980957
transform -1 0 9476 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2879_
timestamp 1688980957
transform -1 0 5612 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2880_
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2881_
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2882_
timestamp 1688980957
transform 1 0 6348 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2883_
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2884_
timestamp 1688980957
transform 1 0 8924 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2885_
timestamp 1688980957
transform 1 0 10672 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2886_
timestamp 1688980957
transform 1 0 11960 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2887_
timestamp 1688980957
transform 1 0 13892 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2888_
timestamp 1688980957
transform -1 0 16008 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2889_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18124 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2890_
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2891_
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2892_
timestamp 1688980957
transform 1 0 15272 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2893_
timestamp 1688980957
transform 1 0 15640 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2894_
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2895_
timestamp 1688980957
transform 1 0 12144 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2896_
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2897_
timestamp 1688980957
transform -1 0 12788 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2898_
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2899_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2900_
timestamp 1688980957
transform 1 0 10304 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2901_
timestamp 1688980957
transform -1 0 13340 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2902_
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2903_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2904_
timestamp 1688980957
transform 1 0 24472 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2905_
timestamp 1688980957
transform 1 0 24656 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2906_
timestamp 1688980957
transform 1 0 22816 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2907_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2908_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2909_
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2910_
timestamp 1688980957
transform 1 0 20976 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2911_
timestamp 1688980957
transform 1 0 20516 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2912_
timestamp 1688980957
transform 1 0 22356 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2913_
timestamp 1688980957
transform -1 0 19136 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2914_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2915_
timestamp 1688980957
transform 1 0 22448 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2916_
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2917_
timestamp 1688980957
transform 1 0 20976 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2918_
timestamp 1688980957
transform 1 0 19504 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2919_
timestamp 1688980957
transform 1 0 19780 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2920_
timestamp 1688980957
transform 1 0 21528 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2921_
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2922_
timestamp 1688980957
transform 1 0 24380 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2923_
timestamp 1688980957
transform 1 0 24932 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2924_
timestamp 1688980957
transform 1 0 22080 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2925_
timestamp 1688980957
transform 1 0 15272 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2926_
timestamp 1688980957
transform 1 0 17296 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2927_
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2928_
timestamp 1688980957
transform 1 0 14628 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2929_
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2930_
timestamp 1688980957
transform 1 0 12788 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2931_
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2932_
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2933_
timestamp 1688980957
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2934_
timestamp 1688980957
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2935_
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2936_
timestamp 1688980957
transform 1 0 9384 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2937_
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2938_
timestamp 1688980957
transform 1 0 19228 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2939_
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2940_
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2941_
timestamp 1688980957
transform -1 0 26220 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2942_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2943_
timestamp 1688980957
transform 1 0 23920 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2944_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2945_
timestamp 1688980957
transform 1 0 19504 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2946_
timestamp 1688980957
transform 1 0 17388 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2947_
timestamp 1688980957
transform 1 0 15640 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2948_
timestamp 1688980957
transform 1 0 12420 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2949_
timestamp 1688980957
transform 1 0 7360 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2950_
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2951_
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2952_
timestamp 1688980957
transform 1 0 1472 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2953_
timestamp 1688980957
transform 1 0 4416 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2954_
timestamp 1688980957
transform 1 0 1564 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2955_
timestamp 1688980957
transform 1 0 4600 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2956_
timestamp 1688980957
transform 1 0 8280 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2957_
timestamp 1688980957
transform -1 0 12052 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2958_
timestamp 1688980957
transform 1 0 13248 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2959_
timestamp 1688980957
transform 1 0 15088 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2960_
timestamp 1688980957
transform 1 0 18308 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2961_
timestamp 1688980957
transform 1 0 21988 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2962_
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2963_
timestamp 1688980957
transform 1 0 19504 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2964_
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2965_
timestamp 1688980957
transform 1 0 15364 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2966_
timestamp 1688980957
transform 1 0 10948 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2967_
timestamp 1688980957
transform 1 0 7176 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2968_
timestamp 1688980957
transform 1 0 6716 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2969_
timestamp 1688980957
transform 1 0 3036 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2970_
timestamp 1688980957
transform -1 0 3312 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2971_
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2972_
timestamp 1688980957
transform 1 0 3036 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2973_
timestamp 1688980957
transform -1 0 6532 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2974_
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2975_
timestamp 1688980957
transform 1 0 10120 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2976_
timestamp 1688980957
transform 1 0 12236 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2977_
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2978_
timestamp 1688980957
transform 1 0 17664 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2979_
timestamp 1688980957
transform -1 0 26220 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2980_
timestamp 1688980957
transform 1 0 20700 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2981_
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2982_
timestamp 1688980957
transform 1 0 17388 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2983_
timestamp 1688980957
transform -1 0 17848 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2984_
timestamp 1688980957
transform 1 0 13524 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2985_
timestamp 1688980957
transform 1 0 9476 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2986_
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2987_
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2988_
timestamp 1688980957
transform 1 0 1472 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2989_
timestamp 1688980957
transform 1 0 5152 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2990_
timestamp 1688980957
transform 1 0 1472 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2991_
timestamp 1688980957
transform 1 0 4692 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2992_
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2993_
timestamp 1688980957
transform 1 0 11040 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2994_
timestamp 1688980957
transform -1 0 14812 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2995_
timestamp 1688980957
transform -1 0 17296 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2996_
timestamp 1688980957
transform 1 0 17296 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2997_
timestamp 1688980957
transform -1 0 18124 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2998_
timestamp 1688980957
transform -1 0 16192 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2999_
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _3000_
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3001_
timestamp 1688980957
transform 1 0 18216 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _3002_
timestamp 1688980957
transform -1 0 21712 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _3003_
timestamp 1688980957
transform 1 0 41860 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25852 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform 1 0 34132 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform -1 0 33028 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1688980957
transform 1 0 12144 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1688980957
transform -1 0 19780 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1688980957
transform -1 0 14812 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1688980957
transform 1 0 3864 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1688980957
transform -1 0 5612 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1688980957
transform 1 0 9016 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1688980957
transform -1 0 20792 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1688980957
transform 1 0 19688 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1688980957
transform 1 0 15456 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1688980957
transform 1 0 20976 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1688980957
transform 1 0 24932 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1688980957
transform -1 0 29348 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1688980957
transform 1 0 27140 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1688980957
transform -1 0 28060 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1688980957
transform -1 0 33948 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1688980957
transform 1 0 40572 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1688980957
transform 1 0 42044 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1688980957
transform -1 0 39008 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1688980957
transform -1 0 28796 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1688980957
transform -1 0 33948 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1688980957
transform 1 0 37904 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1688980957
transform 1 0 43056 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_clk
timestamp 1688980957
transform 1 0 39836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1688980957
transform 1 0 42964 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1688980957
transform 1 0 35420 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1688980957
transform -1 0 31372 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1688980957
transform -1 0 31372 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1688980957
transform 1 0 22448 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1688980957
transform -1 0 18676 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_37_clk
timestamp 1688980957
transform -1 0 8832 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_38_clk
timestamp 1688980957
transform -1 0 10212 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_39_clk
timestamp 1688980957
transform -1 0 10580 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1688980957
transform -1 0 6992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1688980957
transform -1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1688980957
transform -1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1688980957
transform -1 0 11040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1688980957
transform -1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1688980957
transform -1 0 24748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1688980957
transform -1 0 36156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1688980957
transform -1 0 35328 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1688980957
transform -1 0 26680 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 1688980957
transform -1 0 24564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1688980957
transform -1 0 38456 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1688980957
transform 1 0 37996 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1688980957
transform -1 0 10304 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1688980957
transform -1 0 13800 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1688980957
transform -1 0 6256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1688980957
transform -1 0 8004 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1688980957
transform 1 0 6992 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1688980957
transform -1 0 16008 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout44
timestamp 1688980957
transform -1 0 14904 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1688980957
transform -1 0 29348 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1688980957
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1688980957
transform 1 0 35604 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1688980957
transform 1 0 41676 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1688980957
transform 1 0 35052 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1688980957
transform -1 0 25668 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1688980957
transform -1 0 25300 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1688980957
transform 1 0 35328 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1688980957
transform 1 0 35788 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1688980957
transform 1 0 25300 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1688980957
transform 1 0 7544 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_273
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_317
timestamp 1688980957
transform 1 0 30268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_329 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_344
timestamp 1688980957
transform 1 0 32752 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_356
timestamp 1688980957
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_461 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_468
timestamp 1688980957
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_98
timestamp 1688980957
transform 1 0 10120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_129
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_141
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_265
timestamp 1688980957
transform 1 0 25484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_272
timestamp 1688980957
transform 1 0 26128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_327
timestamp 1688980957
transform 1 0 31188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_331
timestamp 1688980957
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1688980957
transform 1 0 32476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_345
timestamp 1688980957
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_371
timestamp 1688980957
transform 1 0 35236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_416
timestamp 1688980957
transform 1 0 39376 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_424
timestamp 1688980957
transform 1 0 40112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_51
timestamp 1688980957
transform 1 0 5796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_57
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_100
timestamp 1688980957
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_124
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_132
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_192
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_296
timestamp 1688980957
transform 1 0 28336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_315
timestamp 1688980957
transform 1 0 30084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_380
timestamp 1688980957
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_384
timestamp 1688980957
transform 1 0 36432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_393
timestamp 1688980957
transform 1 0 37260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_397
timestamp 1688980957
transform 1 0 37628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_409
timestamp 1688980957
transform 1 0 38732 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_37
timestamp 1688980957
transform 1 0 4508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_45
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_85
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_121
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_134
timestamp 1688980957
transform 1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_182
timestamp 1688980957
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_213
timestamp 1688980957
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_265
timestamp 1688980957
transform 1 0 25484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_269
timestamp 1688980957
transform 1 0 25852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_287
timestamp 1688980957
transform 1 0 27508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_295
timestamp 1688980957
transform 1 0 28244 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_318
timestamp 1688980957
transform 1 0 30360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_330
timestamp 1688980957
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_345
timestamp 1688980957
transform 1 0 32844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_368
timestamp 1688980957
transform 1 0 34960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_406
timestamp 1688980957
transform 1 0 38456 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_437
timestamp 1688980957
transform 1 0 41308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_469
timestamp 1688980957
transform 1 0 44252 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_475
timestamp 1688980957
transform 1 0 44804 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1688980957
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_92
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_104
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_200
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_206
timestamp 1688980957
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_219
timestamp 1688980957
transform 1 0 21252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_329
timestamp 1688980957
transform 1 0 31372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_341
timestamp 1688980957
transform 1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_402
timestamp 1688980957
transform 1 0 38088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_409
timestamp 1688980957
transform 1 0 38732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_425
timestamp 1688980957
transform 1 0 40204 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_439
timestamp 1688980957
transform 1 0 41492 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_456
timestamp 1688980957
transform 1 0 43056 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_468
timestamp 1688980957
transform 1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_7
timestamp 1688980957
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_44
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp 1688980957
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_117
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_133
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_148
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_160
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_175
timestamp 1688980957
transform 1 0 17204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_183
timestamp 1688980957
transform 1 0 17940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_195
timestamp 1688980957
transform 1 0 19044 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_234
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_253
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_269
timestamp 1688980957
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1688980957
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_287
timestamp 1688980957
transform 1 0 27508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_299
timestamp 1688980957
transform 1 0 28612 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_307
timestamp 1688980957
transform 1 0 29348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_368
timestamp 1688980957
transform 1 0 34960 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_384
timestamp 1688980957
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_413
timestamp 1688980957
transform 1 0 39100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_435
timestamp 1688980957
transform 1 0 41124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_458
timestamp 1688980957
transform 1 0 43240 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_464
timestamp 1688980957
transform 1 0 43792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_118
timestamp 1688980957
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_130
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_134
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_152
timestamp 1688980957
transform 1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_169
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_184
timestamp 1688980957
transform 1 0 18032 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_213
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_220
timestamp 1688980957
transform 1 0 21344 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_232
timestamp 1688980957
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_244
timestamp 1688980957
transform 1 0 23552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_329
timestamp 1688980957
transform 1 0 31372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_343
timestamp 1688980957
transform 1 0 32660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_359
timestamp 1688980957
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_397
timestamp 1688980957
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_402
timestamp 1688980957
transform 1 0 38088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_414
timestamp 1688980957
transform 1 0 39192 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_453
timestamp 1688980957
transform 1 0 42780 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_107
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_141
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_148
timestamp 1688980957
transform 1 0 14720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_162
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_180
timestamp 1688980957
transform 1 0 17664 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_199
timestamp 1688980957
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_206
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_218
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_243
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_254
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_269
timestamp 1688980957
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1688980957
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_359
timestamp 1688980957
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_371
timestamp 1688980957
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_383
timestamp 1688980957
transform 1 0 36340 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_406
timestamp 1688980957
transform 1 0 38456 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_418
timestamp 1688980957
transform 1 0 39560 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_430
timestamp 1688980957
transform 1 0 40664 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_442
timestamp 1688980957
transform 1 0 41768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_463
timestamp 1688980957
transform 1 0 43700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_471
timestamp 1688980957
transform 1 0 44436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_49
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_154
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_163
timestamp 1688980957
transform 1 0 16100 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_174
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_237
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_250
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_273
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_282
timestamp 1688980957
transform 1 0 27048 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_287
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_299
timestamp 1688980957
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_332
timestamp 1688980957
transform 1 0 31648 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_338
timestamp 1688980957
transform 1 0 32200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_359
timestamp 1688980957
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_394
timestamp 1688980957
transform 1 0 37352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_455
timestamp 1688980957
transform 1 0 42964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_71
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_83
timestamp 1688980957
transform 1 0 8740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_95
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_127
timestamp 1688980957
transform 1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_139
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_150
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_157
timestamp 1688980957
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1688980957
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_229
timestamp 1688980957
transform 1 0 22172 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_244
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_256
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_270
timestamp 1688980957
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_302
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_314
timestamp 1688980957
transform 1 0 29992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_326
timestamp 1688980957
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_334
timestamp 1688980957
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_380
timestamp 1688980957
transform 1 0 36064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_423
timestamp 1688980957
transform 1 0 40020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_430
timestamp 1688980957
transform 1 0 40664 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_436
timestamp 1688980957
transform 1 0 41216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_453
timestamp 1688980957
transform 1 0 42780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_475
timestamp 1688980957
transform 1 0 44804 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_182
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_212
timestamp 1688980957
transform 1 0 20608 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_220
timestamp 1688980957
transform 1 0 21344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_226
timestamp 1688980957
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_314
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_329
timestamp 1688980957
transform 1 0 31372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_341
timestamp 1688980957
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_353
timestamp 1688980957
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 1688980957
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_399
timestamp 1688980957
transform 1 0 37812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_411
timestamp 1688980957
transform 1 0 38916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_416
timestamp 1688980957
transform 1 0 39376 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_441
timestamp 1688980957
transform 1 0 41676 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_463
timestamp 1688980957
transform 1 0 43700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_123
timestamp 1688980957
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_135
timestamp 1688980957
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_153
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_159
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_180
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_192
timestamp 1688980957
transform 1 0 18768 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_229
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_241
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_271
timestamp 1688980957
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_290
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_354
timestamp 1688980957
transform 1 0 33672 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_381
timestamp 1688980957
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_425
timestamp 1688980957
transform 1 0 40204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_433
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_442
timestamp 1688980957
transform 1 0 41768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_465
timestamp 1688980957
transform 1 0 43884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_113
timestamp 1688980957
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_127
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_157
timestamp 1688980957
transform 1 0 15548 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_185
timestamp 1688980957
transform 1 0 18124 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_210
timestamp 1688980957
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_222
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_230
timestamp 1688980957
transform 1 0 22264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_241
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_271
timestamp 1688980957
transform 1 0 26036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_283
timestamp 1688980957
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_288
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_292
timestamp 1688980957
transform 1 0 27968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_298
timestamp 1688980957
transform 1 0 28520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_305
timestamp 1688980957
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_325
timestamp 1688980957
transform 1 0 31004 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_340
timestamp 1688980957
transform 1 0 32384 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_360
timestamp 1688980957
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_393
timestamp 1688980957
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_399
timestamp 1688980957
transform 1 0 37812 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_405
timestamp 1688980957
transform 1 0 38364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_417
timestamp 1688980957
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_426
timestamp 1688980957
transform 1 0 40296 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_438
timestamp 1688980957
transform 1 0 41400 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_452
timestamp 1688980957
transform 1 0 42688 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_456
timestamp 1688980957
transform 1 0 43056 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_468
timestamp 1688980957
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_127
timestamp 1688980957
transform 1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_135
timestamp 1688980957
transform 1 0 13524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_151
timestamp 1688980957
transform 1 0 14996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_172
timestamp 1688980957
transform 1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_212
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_239
timestamp 1688980957
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_254
timestamp 1688980957
transform 1 0 24472 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_266
timestamp 1688980957
transform 1 0 25576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_276
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_290
timestamp 1688980957
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_302
timestamp 1688980957
transform 1 0 28888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_319
timestamp 1688980957
transform 1 0 30452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_345
timestamp 1688980957
transform 1 0 32844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_368
timestamp 1688980957
transform 1 0 34960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_383
timestamp 1688980957
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_403
timestamp 1688980957
transform 1 0 38180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_416
timestamp 1688980957
transform 1 0 39376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_427
timestamp 1688980957
transform 1 0 40388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_435
timestamp 1688980957
transform 1 0 41124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 1688980957
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_454
timestamp 1688980957
transform 1 0 42872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_466
timestamp 1688980957
transform 1 0 43976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_474
timestamp 1688980957
transform 1 0 44712 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_105
timestamp 1688980957
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_151
timestamp 1688980957
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_163
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_171
timestamp 1688980957
transform 1 0 16836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_183
timestamp 1688980957
transform 1 0 17940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_217
timestamp 1688980957
transform 1 0 21068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_235
timestamp 1688980957
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_247
timestamp 1688980957
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_263
timestamp 1688980957
transform 1 0 25300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_288
timestamp 1688980957
transform 1 0 27600 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_296
timestamp 1688980957
transform 1 0 28336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_327
timestamp 1688980957
transform 1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_336
timestamp 1688980957
transform 1 0 32016 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_348
timestamp 1688980957
transform 1 0 33120 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_356
timestamp 1688980957
transform 1 0 33856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_461
timestamp 1688980957
transform 1 0 43516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_473
timestamp 1688980957
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_120
timestamp 1688980957
transform 1 0 12144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_129
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1688980957
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_153
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_179
timestamp 1688980957
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_191
timestamp 1688980957
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_206
timestamp 1688980957
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_238
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_265
timestamp 1688980957
transform 1 0 25484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_275
timestamp 1688980957
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_288
timestamp 1688980957
transform 1 0 27600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_328
timestamp 1688980957
transform 1 0 31280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_342
timestamp 1688980957
transform 1 0 32568 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_350
timestamp 1688980957
transform 1 0 33304 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_401
timestamp 1688980957
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_425
timestamp 1688980957
transform 1 0 40204 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_436
timestamp 1688980957
transform 1 0 41216 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_473
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_190
timestamp 1688980957
transform 1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_204
timestamp 1688980957
transform 1 0 19872 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_216
timestamp 1688980957
transform 1 0 20976 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_228
timestamp 1688980957
transform 1 0 22080 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_236
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1688980957
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_257
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_266
timestamp 1688980957
transform 1 0 25576 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_278
timestamp 1688980957
transform 1 0 26680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_290
timestamp 1688980957
transform 1 0 27784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1688980957
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_340
timestamp 1688980957
transform 1 0 32384 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_352
timestamp 1688980957
transform 1 0 33488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_379
timestamp 1688980957
transform 1 0 35972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_414
timestamp 1688980957
transform 1 0 39192 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 1688980957
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 1688980957
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 1688980957
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_133
timestamp 1688980957
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_140
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_214
timestamp 1688980957
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1688980957
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_275
timestamp 1688980957
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_291
timestamp 1688980957
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_295
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_300
timestamp 1688980957
transform 1 0 28704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_306
timestamp 1688980957
transform 1 0 29256 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_312
timestamp 1688980957
transform 1 0 29808 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_318
timestamp 1688980957
transform 1 0 30360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_322
timestamp 1688980957
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_332
timestamp 1688980957
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_342
timestamp 1688980957
transform 1 0 32568 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_354
timestamp 1688980957
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_372
timestamp 1688980957
transform 1 0 35328 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_384
timestamp 1688980957
transform 1 0 36432 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_401
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_413
timestamp 1688980957
transform 1 0 39100 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_425
timestamp 1688980957
transform 1 0 40204 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_437
timestamp 1688980957
transform 1 0 41308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_445
timestamp 1688980957
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_473
timestamp 1688980957
transform 1 0 44620 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_129
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_156
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_173
timestamp 1688980957
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_180
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 1688980957
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_215
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_224
timestamp 1688980957
transform 1 0 21712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_243
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_295
timestamp 1688980957
transform 1 0 28244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_299
timestamp 1688980957
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_314
timestamp 1688980957
transform 1 0 29992 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_339
timestamp 1688980957
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_351
timestamp 1688980957
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_371
timestamp 1688980957
transform 1 0 35236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_379
timestamp 1688980957
transform 1 0 35972 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_400
timestamp 1688980957
transform 1 0 37904 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_412
timestamp 1688980957
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_68
timestamp 1688980957
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_75
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_87
timestamp 1688980957
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_95
timestamp 1688980957
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_107
timestamp 1688980957
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_134
timestamp 1688980957
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_146
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_157
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_174
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_189
timestamp 1688980957
transform 1 0 18492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_197
timestamp 1688980957
transform 1 0 19228 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_229
timestamp 1688980957
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_234
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_256
timestamp 1688980957
transform 1 0 24656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_262
timestamp 1688980957
transform 1 0 25208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_272
timestamp 1688980957
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_285
timestamp 1688980957
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_290
timestamp 1688980957
transform 1 0 27784 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_302
timestamp 1688980957
transform 1 0 28888 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_313
timestamp 1688980957
transform 1 0 29900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_321
timestamp 1688980957
transform 1 0 30636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_334
timestamp 1688980957
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_347
timestamp 1688980957
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_359
timestamp 1688980957
transform 1 0 34132 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_371
timestamp 1688980957
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_383
timestamp 1688980957
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_431
timestamp 1688980957
transform 1 0 40756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_443
timestamp 1688980957
transform 1 0 41860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1688980957
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_457
timestamp 1688980957
transform 1 0 43148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_462
timestamp 1688980957
transform 1 0 43608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_471
timestamp 1688980957
transform 1 0 44436 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_475
timestamp 1688980957
transform 1 0 44804 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_59
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_105
timestamp 1688980957
transform 1 0 10764 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_111
timestamp 1688980957
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_118
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_124
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_225
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_230
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_264
timestamp 1688980957
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_268
timestamp 1688980957
transform 1 0 25760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_273
timestamp 1688980957
transform 1 0 26220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_327
timestamp 1688980957
transform 1 0 31188 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_341
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_353
timestamp 1688980957
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_371
timestamp 1688980957
transform 1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_383
timestamp 1688980957
transform 1 0 36340 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_398
timestamp 1688980957
transform 1 0 37720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_410
timestamp 1688980957
transform 1 0 38824 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_418
timestamp 1688980957
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_437
timestamp 1688980957
transform 1 0 41308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_445
timestamp 1688980957
transform 1 0 42044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_468
timestamp 1688980957
transform 1 0 44160 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_130
timestamp 1688980957
transform 1 0 13064 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_156
timestamp 1688980957
transform 1 0 15456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_189
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_196
timestamp 1688980957
transform 1 0 19136 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_208
timestamp 1688980957
transform 1 0 20240 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1688980957
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_263
timestamp 1688980957
transform 1 0 25300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_299
timestamp 1688980957
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_306
timestamp 1688980957
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_318
timestamp 1688980957
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_365
timestamp 1688980957
transform 1 0 34684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_388
timestamp 1688980957
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_419
timestamp 1688980957
transform 1 0 39652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 1688980957
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 1688980957
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_473
timestamp 1688980957
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_106
timestamp 1688980957
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_122
timestamp 1688980957
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_161
timestamp 1688980957
transform 1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_170
timestamp 1688980957
transform 1 0 16744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_187
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_215
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_227
timestamp 1688980957
transform 1 0 21988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_239
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_270
timestamp 1688980957
transform 1 0 25944 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_284
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_296
timestamp 1688980957
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_324
timestamp 1688980957
transform 1 0 30912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_332
timestamp 1688980957
transform 1 0 31648 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_341
timestamp 1688980957
transform 1 0 32476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_353
timestamp 1688980957
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_361
timestamp 1688980957
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_385
timestamp 1688980957
transform 1 0 36524 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_397
timestamp 1688980957
transform 1 0 37628 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_409
timestamp 1688980957
transform 1 0 38732 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_417
timestamp 1688980957
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1688980957
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 1688980957
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_77
timestamp 1688980957
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_121
timestamp 1688980957
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_127
timestamp 1688980957
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_132
timestamp 1688980957
transform 1 0 13248 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_138
timestamp 1688980957
transform 1 0 13800 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_184
timestamp 1688980957
transform 1 0 18032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_196
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_243
timestamp 1688980957
transform 1 0 23460 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_255
timestamp 1688980957
transform 1 0 24564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_263
timestamp 1688980957
transform 1 0 25300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_275
timestamp 1688980957
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_290
timestamp 1688980957
transform 1 0 27784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_302
timestamp 1688980957
transform 1 0 28888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_306
timestamp 1688980957
transform 1 0 29256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_333
timestamp 1688980957
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_374
timestamp 1688980957
transform 1 0 35512 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_383
timestamp 1688980957
transform 1 0 36340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_401
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_413
timestamp 1688980957
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_425
timestamp 1688980957
transform 1 0 40204 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_437
timestamp 1688980957
transform 1 0 41308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_445
timestamp 1688980957
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_461
timestamp 1688980957
transform 1 0 43516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_470
timestamp 1688980957
transform 1 0 44344 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_105
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_111
timestamp 1688980957
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_148
timestamp 1688980957
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_152
timestamp 1688980957
transform 1 0 15088 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_159
timestamp 1688980957
transform 1 0 15732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_167
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_173
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_185
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_208
timestamp 1688980957
transform 1 0 20240 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_244
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_269
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_285
timestamp 1688980957
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_297
timestamp 1688980957
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_305
timestamp 1688980957
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_339
timestamp 1688980957
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_351
timestamp 1688980957
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_399
timestamp 1688980957
transform 1 0 37812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_405
timestamp 1688980957
transform 1 0 38364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_414
timestamp 1688980957
transform 1 0 39192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_441
timestamp 1688980957
transform 1 0 41676 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_463
timestamp 1688980957
transform 1 0 43700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 1688980957
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_65
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_79
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_87
timestamp 1688980957
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_155
timestamp 1688980957
transform 1 0 15364 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_180
timestamp 1688980957
transform 1 0 17664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_192
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_198
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_203
timestamp 1688980957
transform 1 0 19780 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_215
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_236
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_244
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_268
timestamp 1688980957
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_287
timestamp 1688980957
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_309
timestamp 1688980957
transform 1 0 29532 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_323
timestamp 1688980957
transform 1 0 30820 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_382
timestamp 1688980957
transform 1 0 36248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_390
timestamp 1688980957
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_407
timestamp 1688980957
transform 1 0 38548 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_419
timestamp 1688980957
transform 1 0 39652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_431
timestamp 1688980957
transform 1 0 40756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_443
timestamp 1688980957
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1688980957
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_457
timestamp 1688980957
transform 1 0 43148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_467
timestamp 1688980957
transform 1 0 44068 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_475
timestamp 1688980957
transform 1 0 44804 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_61
timestamp 1688980957
transform 1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_95
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_107
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_119
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_131
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_168
timestamp 1688980957
transform 1 0 16560 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_263
timestamp 1688980957
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_275
timestamp 1688980957
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_287
timestamp 1688980957
transform 1 0 27508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_329
timestamp 1688980957
transform 1 0 31372 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_337
timestamp 1688980957
transform 1 0 32108 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_349
timestamp 1688980957
transform 1 0 33212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_361
timestamp 1688980957
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_416
timestamp 1688980957
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1688980957
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1688980957
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 1688980957
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_469
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_65
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_70
timestamp 1688980957
transform 1 0 7544 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_82
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_94
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1688980957
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_192
timestamp 1688980957
transform 1 0 18768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_206
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_211
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_233
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_245
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_257
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1688980957
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_301
timestamp 1688980957
transform 1 0 28796 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_327
timestamp 1688980957
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_374
timestamp 1688980957
transform 1 0 35512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_386
timestamp 1688980957
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_404
timestamp 1688980957
transform 1 0 38272 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_416
timestamp 1688980957
transform 1 0 39376 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_428
timestamp 1688980957
transform 1 0 40480 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_440
timestamp 1688980957
transform 1 0 41584 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 1688980957
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_473
timestamp 1688980957
transform 1 0 44620 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_66
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_78
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_134
timestamp 1688980957
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_161
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_166
timestamp 1688980957
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_178
timestamp 1688980957
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_190
timestamp 1688980957
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_269
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_291
timestamp 1688980957
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_295
timestamp 1688980957
transform 1 0 28244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_304
timestamp 1688980957
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_397
timestamp 1688980957
transform 1 0 37628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_409
timestamp 1688980957
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_417
timestamp 1688980957
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 1688980957
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 1688980957
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_98
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_104
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_123
timestamp 1688980957
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_135
timestamp 1688980957
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_147
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_151
timestamp 1688980957
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_158
timestamp 1688980957
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_267
timestamp 1688980957
transform 1 0 25668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_271
timestamp 1688980957
transform 1 0 26036 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_275
timestamp 1688980957
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_345
timestamp 1688980957
transform 1 0 32844 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_377
timestamp 1688980957
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_381
timestamp 1688980957
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_389
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_416
timestamp 1688980957
transform 1 0 39376 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_428
timestamp 1688980957
transform 1 0 40480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_440
timestamp 1688980957
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_473
timestamp 1688980957
transform 1 0 44620 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1688980957
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1688980957
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_100
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_112
timestamp 1688980957
transform 1 0 11408 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_124
timestamp 1688980957
transform 1 0 12512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1688980957
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_144
timestamp 1688980957
transform 1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_155
timestamp 1688980957
transform 1 0 15364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_174
timestamp 1688980957
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_205
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_236
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_262
timestamp 1688980957
transform 1 0 25208 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_270
timestamp 1688980957
transform 1 0 25944 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_281
timestamp 1688980957
transform 1 0 26956 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_322
timestamp 1688980957
transform 1 0 30728 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_330
timestamp 1688980957
transform 1 0 31464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_340
timestamp 1688980957
transform 1 0 32384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_353
timestamp 1688980957
transform 1 0 33580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_378
timestamp 1688980957
transform 1 0 35880 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_406
timestamp 1688980957
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_418
timestamp 1688980957
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 1688980957
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 1688980957
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1688980957
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_159
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_186
timestamp 1688980957
transform 1 0 18216 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_203
timestamp 1688980957
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_211
timestamp 1688980957
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_241
timestamp 1688980957
transform 1 0 23276 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_267
timestamp 1688980957
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_324
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_357
timestamp 1688980957
transform 1 0 33948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_379
timestamp 1688980957
transform 1 0 35972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_398
timestamp 1688980957
transform 1 0 37720 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_410
timestamp 1688980957
transform 1 0 38824 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_422
timestamp 1688980957
transform 1 0 39928 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_434
timestamp 1688980957
transform 1 0 41032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_446
timestamp 1688980957
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 1688980957
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_473
timestamp 1688980957
transform 1 0 44620 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_114
timestamp 1688980957
transform 1 0 11592 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1688980957
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_182
timestamp 1688980957
transform 1 0 17848 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_190
timestamp 1688980957
transform 1 0 18584 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_206
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_218
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_230
timestamp 1688980957
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_273
timestamp 1688980957
transform 1 0 26220 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_278
timestamp 1688980957
transform 1 0 26680 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_290
timestamp 1688980957
transform 1 0 27784 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_298
timestamp 1688980957
transform 1 0 28520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_316
timestamp 1688980957
transform 1 0 30176 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_324
timestamp 1688980957
transform 1 0 30912 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_344
timestamp 1688980957
transform 1 0 32752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_352
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_360
timestamp 1688980957
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_380
timestamp 1688980957
transform 1 0 36064 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_396
timestamp 1688980957
transform 1 0 37536 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_408
timestamp 1688980957
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_415
timestamp 1688980957
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1688980957
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1688980957
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 1688980957
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 1688980957
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 1688980957
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_100
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_212
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1688980957
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_325
timestamp 1688980957
transform 1 0 31004 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_346
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_358
timestamp 1688980957
transform 1 0 34040 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_370
timestamp 1688980957
transform 1 0 35144 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_378
timestamp 1688980957
transform 1 0 35880 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_382
timestamp 1688980957
transform 1 0 36248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_390
timestamp 1688980957
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_399
timestamp 1688980957
transform 1 0 37812 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_423
timestamp 1688980957
transform 1 0 40020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_435
timestamp 1688980957
transform 1 0 41124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1688980957
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_473
timestamp 1688980957
transform 1 0 44620 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_111
timestamp 1688980957
transform 1 0 11316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_149
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_161
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_173
timestamp 1688980957
transform 1 0 17020 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 1688980957
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_232
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_340
timestamp 1688980957
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_352
timestamp 1688980957
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_373
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_401
timestamp 1688980957
transform 1 0 37996 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_417
timestamp 1688980957
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_457
timestamp 1688980957
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 1688980957
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_156
timestamp 1688980957
transform 1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_162
timestamp 1688980957
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_178
timestamp 1688980957
transform 1 0 17480 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_192
timestamp 1688980957
transform 1 0 18768 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_241
timestamp 1688980957
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_270
timestamp 1688980957
transform 1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_275
timestamp 1688980957
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_290
timestamp 1688980957
transform 1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_313
timestamp 1688980957
transform 1 0 29900 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_325
timestamp 1688980957
transform 1 0 31004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_369
timestamp 1688980957
transform 1 0 35052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_401
timestamp 1688980957
transform 1 0 37996 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_418
timestamp 1688980957
transform 1 0 39560 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_430
timestamp 1688980957
transform 1 0 40664 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_442
timestamp 1688980957
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 1688980957
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_473
timestamp 1688980957
transform 1 0 44620 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_136
timestamp 1688980957
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_170
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_180
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_184
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_241
timestamp 1688980957
transform 1 0 23276 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_247
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_262
timestamp 1688980957
transform 1 0 25208 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_268
timestamp 1688980957
transform 1 0 25760 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 1688980957
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_316
timestamp 1688980957
transform 1 0 30176 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_328
timestamp 1688980957
transform 1 0 31280 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_340
timestamp 1688980957
transform 1 0 32384 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_352
timestamp 1688980957
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_368
timestamp 1688980957
transform 1 0 34960 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_378
timestamp 1688980957
transform 1 0 35880 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_429
timestamp 1688980957
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_441
timestamp 1688980957
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_453
timestamp 1688980957
transform 1 0 42780 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_465
timestamp 1688980957
transform 1 0 43884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_473
timestamp 1688980957
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_95
timestamp 1688980957
transform 1 0 9844 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_107
timestamp 1688980957
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_129
timestamp 1688980957
transform 1 0 12972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_141
timestamp 1688980957
transform 1 0 14076 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_146
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_150
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_177
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_206
timestamp 1688980957
transform 1 0 20056 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_213
timestamp 1688980957
transform 1 0 20700 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 1688980957
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_247
timestamp 1688980957
transform 1 0 23828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_270
timestamp 1688980957
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_278
timestamp 1688980957
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_313
timestamp 1688980957
transform 1 0 29900 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_321
timestamp 1688980957
transform 1 0 30636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_333
timestamp 1688980957
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_360
timestamp 1688980957
transform 1 0 34224 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_368
timestamp 1688980957
transform 1 0 34960 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_417
timestamp 1688980957
transform 1 0 39468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_421
timestamp 1688980957
transform 1 0 39836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_429
timestamp 1688980957
transform 1 0 40572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_433
timestamp 1688980957
transform 1 0 40940 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_442
timestamp 1688980957
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_473
timestamp 1688980957
transform 1 0 44620 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_88
timestamp 1688980957
transform 1 0 9200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_168
timestamp 1688980957
transform 1 0 16560 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_202
timestamp 1688980957
transform 1 0 19688 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_241
timestamp 1688980957
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1688980957
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_280
timestamp 1688980957
transform 1 0 26864 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_286
timestamp 1688980957
transform 1 0 27416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_295
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_303
timestamp 1688980957
transform 1 0 28980 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_314
timestamp 1688980957
transform 1 0 29992 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_330
timestamp 1688980957
transform 1 0 31464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_334
timestamp 1688980957
transform 1 0 31832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_386
timestamp 1688980957
transform 1 0 36616 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_398
timestamp 1688980957
transform 1 0 37720 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 1688980957
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_460
timestamp 1688980957
transform 1 0 43424 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_472
timestamp 1688980957
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_138
timestamp 1688980957
transform 1 0 13800 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_150
timestamp 1688980957
transform 1 0 14904 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_182
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_219
timestamp 1688980957
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_231
timestamp 1688980957
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_269
timestamp 1688980957
transform 1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_278
timestamp 1688980957
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_309
timestamp 1688980957
transform 1 0 29532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_321
timestamp 1688980957
transform 1 0 30636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_333
timestamp 1688980957
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_344
timestamp 1688980957
transform 1 0 32752 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_356
timestamp 1688980957
transform 1 0 33856 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_368
timestamp 1688980957
transform 1 0 34960 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_386
timestamp 1688980957
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_407
timestamp 1688980957
transform 1 0 38548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_89
timestamp 1688980957
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_108
timestamp 1688980957
transform 1 0 11040 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_129
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_147
timestamp 1688980957
transform 1 0 14628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_161
timestamp 1688980957
transform 1 0 15916 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_185
timestamp 1688980957
transform 1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_205
timestamp 1688980957
transform 1 0 19964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_229
timestamp 1688980957
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_241
timestamp 1688980957
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_257
timestamp 1688980957
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_275
timestamp 1688980957
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_287
timestamp 1688980957
transform 1 0 27508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_297
timestamp 1688980957
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_313
timestamp 1688980957
transform 1 0 29900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_325
timestamp 1688980957
transform 1 0 31004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_337
timestamp 1688980957
transform 1 0 32108 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_350
timestamp 1688980957
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_373
timestamp 1688980957
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_414
timestamp 1688980957
transform 1 0 39192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_474
timestamp 1688980957
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_109
timestamp 1688980957
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_121
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_179
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_192
timestamp 1688980957
transform 1 0 18768 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_213
timestamp 1688980957
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_243
timestamp 1688980957
transform 1 0 23460 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_255
timestamp 1688980957
transform 1 0 24564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_301
timestamp 1688980957
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_309
timestamp 1688980957
transform 1 0 29532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_321
timestamp 1688980957
transform 1 0 30636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_333
timestamp 1688980957
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_354
timestamp 1688980957
transform 1 0 33672 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_370
timestamp 1688980957
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_382
timestamp 1688980957
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_390
timestamp 1688980957
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_399
timestamp 1688980957
transform 1 0 37812 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_416
timestamp 1688980957
transform 1 0 39376 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_432
timestamp 1688980957
transform 1 0 40848 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_440
timestamp 1688980957
transform 1 0 41584 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_444
timestamp 1688980957
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_94
timestamp 1688980957
transform 1 0 9752 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_98
timestamp 1688980957
transform 1 0 10120 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_116
timestamp 1688980957
transform 1 0 11776 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_128
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_150
timestamp 1688980957
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_216
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_228
timestamp 1688980957
transform 1 0 22080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_287
timestamp 1688980957
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_299
timestamp 1688980957
transform 1 0 28612 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_314
timestamp 1688980957
transform 1 0 29992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_326
timestamp 1688980957
transform 1 0 31096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_353
timestamp 1688980957
transform 1 0 33580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_361
timestamp 1688980957
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_386
timestamp 1688980957
transform 1 0 36616 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_405
timestamp 1688980957
transform 1 0 38364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_417
timestamp 1688980957
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_441
timestamp 1688980957
transform 1 0 41676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_456
timestamp 1688980957
transform 1 0 43056 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_460
timestamp 1688980957
transform 1 0 43424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_464
timestamp 1688980957
transform 1 0 43792 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_89
timestamp 1688980957
transform 1 0 9292 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_142
timestamp 1688980957
transform 1 0 14168 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_154
timestamp 1688980957
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_178
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_188
timestamp 1688980957
transform 1 0 18400 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_196
timestamp 1688980957
transform 1 0 19136 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_219
timestamp 1688980957
transform 1 0 21252 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_234
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_247
timestamp 1688980957
transform 1 0 23828 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_260
timestamp 1688980957
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_272
timestamp 1688980957
transform 1 0 26128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_276
timestamp 1688980957
transform 1 0 26496 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_302
timestamp 1688980957
transform 1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_311
timestamp 1688980957
transform 1 0 29716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_323
timestamp 1688980957
transform 1 0 30820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_327
timestamp 1688980957
transform 1 0 31188 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_359
timestamp 1688980957
transform 1 0 34132 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_371
timestamp 1688980957
transform 1 0 35236 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_383
timestamp 1688980957
transform 1 0 36340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_407
timestamp 1688980957
transform 1 0 38548 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_426
timestamp 1688980957
transform 1 0 40296 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_432
timestamp 1688980957
transform 1 0 40848 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_438
timestamp 1688980957
transform 1 0 41400 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_446
timestamp 1688980957
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_456
timestamp 1688980957
transform 1 0 43056 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_474
timestamp 1688980957
transform 1 0 44712 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_122
timestamp 1688980957
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_134
timestamp 1688980957
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_160
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_167
timestamp 1688980957
transform 1 0 16468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_246
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_273
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_285
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_297
timestamp 1688980957
transform 1 0 28428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_316
timestamp 1688980957
transform 1 0 30176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_370
timestamp 1688980957
transform 1 0 35144 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_78
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_87
timestamp 1688980957
transform 1 0 9108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_99
timestamp 1688980957
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_121
timestamp 1688980957
transform 1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_152
timestamp 1688980957
transform 1 0 15088 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_164
timestamp 1688980957
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_186
timestamp 1688980957
transform 1 0 18216 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_198
timestamp 1688980957
transform 1 0 19320 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_210
timestamp 1688980957
transform 1 0 20424 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_240
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_269
timestamp 1688980957
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_277
timestamp 1688980957
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_290
timestamp 1688980957
transform 1 0 27784 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_296
timestamp 1688980957
transform 1 0 28336 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_323
timestamp 1688980957
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_357
timestamp 1688980957
transform 1 0 33948 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_372
timestamp 1688980957
transform 1 0 35328 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_468
timestamp 1688980957
transform 1 0 44160 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_61
timestamp 1688980957
transform 1 0 6716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_91
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_100
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_112
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_118
timestamp 1688980957
transform 1 0 11960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_164
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_176
timestamp 1688980957
transform 1 0 17296 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_188
timestamp 1688980957
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_203
timestamp 1688980957
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_210
timestamp 1688980957
transform 1 0 20424 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_222
timestamp 1688980957
transform 1 0 21528 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_250
timestamp 1688980957
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_262
timestamp 1688980957
transform 1 0 25208 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_274
timestamp 1688980957
transform 1 0 26312 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_299
timestamp 1688980957
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_407
timestamp 1688980957
transform 1 0 38548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_417
timestamp 1688980957
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_432
timestamp 1688980957
transform 1 0 40848 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_444
timestamp 1688980957
transform 1 0 41952 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_456
timestamp 1688980957
transform 1 0 43056 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_468
timestamp 1688980957
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_6
timestamp 1688980957
transform 1 0 1656 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_18
timestamp 1688980957
transform 1 0 2760 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_26
timestamp 1688980957
transform 1 0 3496 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_65
timestamp 1688980957
transform 1 0 7084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_121
timestamp 1688980957
transform 1 0 12236 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_138
timestamp 1688980957
transform 1 0 13800 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_154
timestamp 1688980957
transform 1 0 15272 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_166
timestamp 1688980957
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_203
timestamp 1688980957
transform 1 0 19780 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_221
timestamp 1688980957
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_233
timestamp 1688980957
transform 1 0 22540 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_248
timestamp 1688980957
transform 1 0 23920 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_254
timestamp 1688980957
transform 1 0 24472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_275
timestamp 1688980957
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_365
timestamp 1688980957
transform 1 0 34684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_389
timestamp 1688980957
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_405
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_409
timestamp 1688980957
transform 1 0 38732 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_413
timestamp 1688980957
transform 1 0 39100 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_422
timestamp 1688980957
transform 1 0 39928 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_434
timestamp 1688980957
transform 1 0 41032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_446
timestamp 1688980957
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_471
timestamp 1688980957
transform 1 0 44436 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_475
timestamp 1688980957
transform 1 0 44804 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_62
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_103
timestamp 1688980957
transform 1 0 10580 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_112
timestamp 1688980957
transform 1 0 11408 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_124
timestamp 1688980957
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_173
timestamp 1688980957
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_229
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_241
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_275
timestamp 1688980957
transform 1 0 26404 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_287
timestamp 1688980957
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_299
timestamp 1688980957
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1688980957
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_375
timestamp 1688980957
transform 1 0 35604 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_382
timestamp 1688980957
transform 1 0 36248 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_394
timestamp 1688980957
transform 1 0 37352 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_406
timestamp 1688980957
transform 1 0 38456 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 1688980957
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 1688980957
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_47
timestamp 1688980957
transform 1 0 5428 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1688980957
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_60
timestamp 1688980957
transform 1 0 6624 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_72
timestamp 1688980957
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_84
timestamp 1688980957
transform 1 0 8832 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_96
timestamp 1688980957
transform 1 0 9936 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_118
timestamp 1688980957
transform 1 0 11960 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_128
timestamp 1688980957
transform 1 0 12880 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_140
timestamp 1688980957
transform 1 0 13984 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_209
timestamp 1688980957
transform 1 0 20332 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_213
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_241
timestamp 1688980957
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_301
timestamp 1688980957
transform 1 0 28796 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_309
timestamp 1688980957
transform 1 0 29532 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_321
timestamp 1688980957
transform 1 0 30636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_333
timestamp 1688980957
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_340
timestamp 1688980957
transform 1 0 32384 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_352
timestamp 1688980957
transform 1 0 33488 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_364
timestamp 1688980957
transform 1 0 34592 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_382
timestamp 1688980957
transform 1 0 36248 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_390
timestamp 1688980957
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_428
timestamp 1688980957
transform 1 0 40480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_449
timestamp 1688980957
transform 1 0 42412 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_100
timestamp 1688980957
transform 1 0 10304 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_108
timestamp 1688980957
transform 1 0 11040 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_112
timestamp 1688980957
transform 1 0 11408 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_124
timestamp 1688980957
transform 1 0 12512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_136
timestamp 1688980957
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_144
timestamp 1688980957
transform 1 0 14352 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_152
timestamp 1688980957
transform 1 0 15088 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_160
timestamp 1688980957
transform 1 0 15824 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_172
timestamp 1688980957
transform 1 0 16928 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_184
timestamp 1688980957
transform 1 0 18032 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_201
timestamp 1688980957
transform 1 0 19596 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_211
timestamp 1688980957
transform 1 0 20516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_223
timestamp 1688980957
transform 1 0 21620 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_227
timestamp 1688980957
transform 1 0 21988 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_239
timestamp 1688980957
transform 1 0 23092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_261
timestamp 1688980957
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_273
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_292
timestamp 1688980957
transform 1 0 27968 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_300
timestamp 1688980957
transform 1 0 28704 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_323
timestamp 1688980957
transform 1 0 30820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_331
timestamp 1688980957
transform 1 0 31556 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_341
timestamp 1688980957
transform 1 0 32476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_347
timestamp 1688980957
transform 1 0 33028 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_356
timestamp 1688980957
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_371
timestamp 1688980957
transform 1 0 35236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_418
timestamp 1688980957
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_446
timestamp 1688980957
transform 1 0 42136 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_456
timestamp 1688980957
transform 1 0 43056 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_460
timestamp 1688980957
transform 1 0 43424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_465
timestamp 1688980957
transform 1 0 43884 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_473
timestamp 1688980957
transform 1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_54
timestamp 1688980957
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_89
timestamp 1688980957
transform 1 0 9292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_101
timestamp 1688980957
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_109
timestamp 1688980957
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_121
timestamp 1688980957
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_128
timestamp 1688980957
transform 1 0 12880 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_140
timestamp 1688980957
transform 1 0 13984 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_152
timestamp 1688980957
transform 1 0 15088 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_160
timestamp 1688980957
transform 1 0 15824 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_173
timestamp 1688980957
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_185
timestamp 1688980957
transform 1 0 18124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_218
timestamp 1688980957
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_253
timestamp 1688980957
transform 1 0 24380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_265
timestamp 1688980957
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_301
timestamp 1688980957
transform 1 0 28796 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_307
timestamp 1688980957
transform 1 0 29348 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_314
timestamp 1688980957
transform 1 0 29992 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_326
timestamp 1688980957
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_334
timestamp 1688980957
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_358
timestamp 1688980957
transform 1 0 34040 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_370
timestamp 1688980957
transform 1 0 35144 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_382
timestamp 1688980957
transform 1 0 36248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_390
timestamp 1688980957
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_423
timestamp 1688980957
transform 1 0 40020 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_429
timestamp 1688980957
transform 1 0 40572 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_434
timestamp 1688980957
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_446
timestamp 1688980957
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_449
timestamp 1688980957
transform 1 0 42412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_455
timestamp 1688980957
transform 1 0 42964 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_463
timestamp 1688980957
transform 1 0 43700 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_475
timestamp 1688980957
transform 1 0 44804 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_45
timestamp 1688980957
transform 1 0 5244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_57
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_69
timestamp 1688980957
transform 1 0 7452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_81
timestamp 1688980957
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_88
timestamp 1688980957
transform 1 0 9200 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_101
timestamp 1688980957
transform 1 0 10396 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_105
timestamp 1688980957
transform 1 0 10764 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_150
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_158
timestamp 1688980957
transform 1 0 15640 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_190
timestamp 1688980957
transform 1 0 18584 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_215
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_280
timestamp 1688980957
transform 1 0 26864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_286
timestamp 1688980957
transform 1 0 27416 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_298
timestamp 1688980957
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_306
timestamp 1688980957
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_316
timestamp 1688980957
transform 1 0 30176 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_328
timestamp 1688980957
transform 1 0 31280 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_340
timestamp 1688980957
transform 1 0 32384 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_346
timestamp 1688980957
transform 1 0 32936 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_354
timestamp 1688980957
transform 1 0 33672 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_358
timestamp 1688980957
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_373
timestamp 1688980957
transform 1 0 35420 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_398
timestamp 1688980957
transform 1 0 37720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_410
timestamp 1688980957
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_418
timestamp 1688980957
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_421
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_430
timestamp 1688980957
transform 1 0 40664 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_442
timestamp 1688980957
transform 1 0 41768 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_450
timestamp 1688980957
transform 1 0 42504 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_460
timestamp 1688980957
transform 1 0 43424 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_472
timestamp 1688980957
transform 1 0 44528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_12
timestamp 1688980957
transform 1 0 2208 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_35
timestamp 1688980957
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_47
timestamp 1688980957
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_89
timestamp 1688980957
transform 1 0 9292 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_106
timestamp 1688980957
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_119
timestamp 1688980957
transform 1 0 12052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_128
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_160
timestamp 1688980957
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_188
timestamp 1688980957
transform 1 0 18400 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_220
timestamp 1688980957
transform 1 0 21344 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_292
timestamp 1688980957
transform 1 0 27968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_304
timestamp 1688980957
transform 1 0 29072 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_313
timestamp 1688980957
transform 1 0 29900 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_325
timestamp 1688980957
transform 1 0 31004 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_333
timestamp 1688980957
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_347
timestamp 1688980957
transform 1 0 33028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_351
timestamp 1688980957
transform 1 0 33396 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_379
timestamp 1688980957
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_397
timestamp 1688980957
transform 1 0 37628 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_418
timestamp 1688980957
transform 1 0 39560 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_430
timestamp 1688980957
transform 1 0 40664 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_442
timestamp 1688980957
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_449
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_467
timestamp 1688980957
transform 1 0 44068 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_475
timestamp 1688980957
transform 1 0 44804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_11
timestamp 1688980957
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_23
timestamp 1688980957
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_75
timestamp 1688980957
transform 1 0 8004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_106
timestamp 1688980957
transform 1 0 10856 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_118
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_126
timestamp 1688980957
transform 1 0 12696 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_136
timestamp 1688980957
transform 1 0 13616 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_146
timestamp 1688980957
transform 1 0 14536 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_158
timestamp 1688980957
transform 1 0 15640 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_170
timestamp 1688980957
transform 1 0 16744 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_183
timestamp 1688980957
transform 1 0 17940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_205
timestamp 1688980957
transform 1 0 19964 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_210
timestamp 1688980957
transform 1 0 20424 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_230
timestamp 1688980957
transform 1 0 22264 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_316
timestamp 1688980957
transform 1 0 30176 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_328
timestamp 1688980957
transform 1 0 31280 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_336
timestamp 1688980957
transform 1 0 32016 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_342
timestamp 1688980957
transform 1 0 32568 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_354
timestamp 1688980957
transform 1 0 33672 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_362
timestamp 1688980957
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_373
timestamp 1688980957
transform 1 0 35420 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_401
timestamp 1688980957
transform 1 0 37996 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_415
timestamp 1688980957
transform 1 0 39284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_429
timestamp 1688980957
transform 1 0 40572 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_441
timestamp 1688980957
transform 1 0 41676 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_449
timestamp 1688980957
transform 1 0 42412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_474
timestamp 1688980957
transform 1 0 44712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_20
timestamp 1688980957
transform 1 0 2944 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_50
timestamp 1688980957
transform 1 0 5704 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_78
timestamp 1688980957
transform 1 0 8280 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_90
timestamp 1688980957
transform 1 0 9384 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_96
timestamp 1688980957
transform 1 0 9936 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_108
timestamp 1688980957
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_119
timestamp 1688980957
transform 1 0 12052 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_127
timestamp 1688980957
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_131
timestamp 1688980957
transform 1 0 13156 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_140
timestamp 1688980957
transform 1 0 13984 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_152
timestamp 1688980957
transform 1 0 15088 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_179
timestamp 1688980957
transform 1 0 17572 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_192
timestamp 1688980957
transform 1 0 18768 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_204
timestamp 1688980957
transform 1 0 19872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_210
timestamp 1688980957
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1688980957
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_233
timestamp 1688980957
transform 1 0 22540 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_258
timestamp 1688980957
transform 1 0 24840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_266
timestamp 1688980957
transform 1 0 25576 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_277
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_290
timestamp 1688980957
transform 1 0 27784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_302
timestamp 1688980957
transform 1 0 28888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_312
timestamp 1688980957
transform 1 0 29808 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_320
timestamp 1688980957
transform 1 0 30544 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_326
timestamp 1688980957
transform 1 0 31096 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_330
timestamp 1688980957
transform 1 0 31464 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_342
timestamp 1688980957
transform 1 0 32568 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_350
timestamp 1688980957
transform 1 0 33304 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_362
timestamp 1688980957
transform 1 0 34408 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_374
timestamp 1688980957
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_386
timestamp 1688980957
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_423
timestamp 1688980957
transform 1 0 40020 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1688980957
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_461
timestamp 1688980957
transform 1 0 43516 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_467
timestamp 1688980957
transform 1 0 44068 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_475
timestamp 1688980957
transform 1 0 44804 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_55
timestamp 1688980957
transform 1 0 6164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_93
timestamp 1688980957
transform 1 0 9660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_113
timestamp 1688980957
transform 1 0 11500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_119
timestamp 1688980957
transform 1 0 12052 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_125
timestamp 1688980957
transform 1 0 12604 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_183
timestamp 1688980957
transform 1 0 17940 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_192
timestamp 1688980957
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_303
timestamp 1688980957
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_335
timestamp 1688980957
transform 1 0 31924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_353
timestamp 1688980957
transform 1 0 33580 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_362
timestamp 1688980957
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_398
timestamp 1688980957
transform 1 0 37720 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_409
timestamp 1688980957
transform 1 0 38732 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1688980957
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 1688980957
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 1688980957
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 1688980957
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_7
timestamp 1688980957
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_52
timestamp 1688980957
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_68
timestamp 1688980957
transform 1 0 7360 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_79
timestamp 1688980957
transform 1 0 8372 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_92
timestamp 1688980957
transform 1 0 9568 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_121
timestamp 1688980957
transform 1 0 12236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_133
timestamp 1688980957
transform 1 0 13340 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_139
timestamp 1688980957
transform 1 0 13892 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_158
timestamp 1688980957
transform 1 0 15640 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_177
timestamp 1688980957
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_185
timestamp 1688980957
transform 1 0 18124 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_194
timestamp 1688980957
transform 1 0 18952 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_208
timestamp 1688980957
transform 1 0 20240 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_216
timestamp 1688980957
transform 1 0 20976 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_222
timestamp 1688980957
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_245
timestamp 1688980957
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_287
timestamp 1688980957
transform 1 0 27508 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_312
timestamp 1688980957
transform 1 0 29808 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_334
timestamp 1688980957
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_345
timestamp 1688980957
transform 1 0 32844 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_381
timestamp 1688980957
transform 1 0 36156 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_413
timestamp 1688980957
transform 1 0 39100 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_438
timestamp 1688980957
transform 1 0 41400 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1688980957
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_449
timestamp 1688980957
transform 1 0 42412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_463
timestamp 1688980957
transform 1 0 43700 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_471
timestamp 1688980957
transform 1 0 44436 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_475
timestamp 1688980957
transform 1 0 44804 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_25
timestamp 1688980957
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_45
timestamp 1688980957
transform 1 0 5244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_49
timestamp 1688980957
transform 1 0 5612 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_58
timestamp 1688980957
transform 1 0 6440 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_64
timestamp 1688980957
transform 1 0 6992 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_108
timestamp 1688980957
transform 1 0 11040 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_115
timestamp 1688980957
transform 1 0 11684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_119
timestamp 1688980957
transform 1 0 12052 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_138
timestamp 1688980957
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_145
timestamp 1688980957
transform 1 0 14444 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_154
timestamp 1688980957
transform 1 0 15272 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_188
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_232
timestamp 1688980957
transform 1 0 22448 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_244
timestamp 1688980957
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_258
timestamp 1688980957
transform 1 0 24840 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_270
timestamp 1688980957
transform 1 0 25944 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_282
timestamp 1688980957
transform 1 0 27048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_286
timestamp 1688980957
transform 1 0 27416 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_354
timestamp 1688980957
transform 1 0 33672 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_360
timestamp 1688980957
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_375
timestamp 1688980957
transform 1 0 35604 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_393
timestamp 1688980957
transform 1 0 37260 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_417
timestamp 1688980957
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_441
timestamp 1688980957
transform 1 0 41676 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_472
timestamp 1688980957
transform 1 0 44528 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_14
timestamp 1688980957
transform 1 0 2392 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_26
timestamp 1688980957
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_38
timestamp 1688980957
transform 1 0 4600 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_48
timestamp 1688980957
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_65
timestamp 1688980957
transform 1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_71
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_79
timestamp 1688980957
transform 1 0 8372 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_92
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_100
timestamp 1688980957
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_142
timestamp 1688980957
transform 1 0 14168 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_154
timestamp 1688980957
transform 1 0 15272 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_166
timestamp 1688980957
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_184
timestamp 1688980957
transform 1 0 18032 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_196
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_200
timestamp 1688980957
transform 1 0 19504 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_247
timestamp 1688980957
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_251
timestamp 1688980957
transform 1 0 24196 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_291
timestamp 1688980957
transform 1 0 27876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_303
timestamp 1688980957
transform 1 0 28980 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_315
timestamp 1688980957
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_327
timestamp 1688980957
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_340
timestamp 1688980957
transform 1 0 32384 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_356
timestamp 1688980957
transform 1 0 33856 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_368
timestamp 1688980957
transform 1 0 34960 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_445
timestamp 1688980957
transform 1 0 42044 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_22
timestamp 1688980957
transform 1 0 3128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_59
timestamp 1688980957
transform 1 0 6532 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_91
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_103
timestamp 1688980957
transform 1 0 10580 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_118
timestamp 1688980957
transform 1 0 11960 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_130
timestamp 1688980957
transform 1 0 13064 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_138
timestamp 1688980957
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_181
timestamp 1688980957
transform 1 0 17756 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_191
timestamp 1688980957
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_203
timestamp 1688980957
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_212
timestamp 1688980957
transform 1 0 20608 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_224
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_244
timestamp 1688980957
transform 1 0 23552 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_248
timestamp 1688980957
transform 1 0 23920 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_273
timestamp 1688980957
transform 1 0 26220 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_295
timestamp 1688980957
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_318
timestamp 1688980957
transform 1 0 30360 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_330
timestamp 1688980957
transform 1 0 31464 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_342
timestamp 1688980957
transform 1 0 32568 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_351
timestamp 1688980957
transform 1 0 33396 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_358
timestamp 1688980957
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_371
timestamp 1688980957
transform 1 0 35236 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_393
timestamp 1688980957
transform 1 0 37260 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_410
timestamp 1688980957
transform 1 0 38824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_418
timestamp 1688980957
transform 1 0 39560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_429
timestamp 1688980957
transform 1 0 40572 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_458
timestamp 1688980957
transform 1 0 43240 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_470
timestamp 1688980957
transform 1 0 44344 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_45
timestamp 1688980957
transform 1 0 5244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_76
timestamp 1688980957
transform 1 0 8096 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_84
timestamp 1688980957
transform 1 0 8832 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_116
timestamp 1688980957
transform 1 0 11776 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_128
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_136
timestamp 1688980957
transform 1 0 13616 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_150
timestamp 1688980957
transform 1 0 14904 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_162
timestamp 1688980957
transform 1 0 16008 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_197
timestamp 1688980957
transform 1 0 19228 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_233
timestamp 1688980957
transform 1 0 22540 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_264
timestamp 1688980957
transform 1 0 25392 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_276
timestamp 1688980957
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_328
timestamp 1688980957
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_348
timestamp 1688980957
transform 1 0 33120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_362
timestamp 1688980957
transform 1 0 34408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_371
timestamp 1688980957
transform 1 0 35236 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_378
timestamp 1688980957
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_390
timestamp 1688980957
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_401
timestamp 1688980957
transform 1 0 37996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_413
timestamp 1688980957
transform 1 0 39100 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_425
timestamp 1688980957
transform 1 0 40204 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1688980957
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1688980957
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_473
timestamp 1688980957
transform 1 0 44620 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_32
timestamp 1688980957
transform 1 0 4048 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_47
timestamp 1688980957
transform 1 0 5428 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_55
timestamp 1688980957
transform 1 0 6164 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_76
timestamp 1688980957
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_96
timestamp 1688980957
transform 1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_100
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_128
timestamp 1688980957
transform 1 0 12880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_132
timestamp 1688980957
transform 1 0 13248 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_185
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_216
timestamp 1688980957
transform 1 0 20976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_220
timestamp 1688980957
transform 1 0 21344 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_241
timestamp 1688980957
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_249
timestamp 1688980957
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_270
timestamp 1688980957
transform 1 0 25944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_278
timestamp 1688980957
transform 1 0 26680 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_317
timestamp 1688980957
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_358
timestamp 1688980957
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_385
timestamp 1688980957
transform 1 0 36524 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_397
timestamp 1688980957
transform 1 0 37628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_418
timestamp 1688980957
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_442
timestamp 1688980957
transform 1 0 41768 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_454
timestamp 1688980957
transform 1 0 42872 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_466
timestamp 1688980957
transform 1 0 43976 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_474
timestamp 1688980957
transform 1 0 44712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_32
timestamp 1688980957
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_44
timestamp 1688980957
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_77
timestamp 1688980957
transform 1 0 8188 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_89
timestamp 1688980957
transform 1 0 9292 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_101
timestamp 1688980957
transform 1 0 10396 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_121
timestamp 1688980957
transform 1 0 12236 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_133
timestamp 1688980957
transform 1 0 13340 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_145
timestamp 1688980957
transform 1 0 14444 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_157
timestamp 1688980957
transform 1 0 15548 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_165
timestamp 1688980957
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_178
timestamp 1688980957
transform 1 0 17480 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_190
timestamp 1688980957
transform 1 0 18584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_198
timestamp 1688980957
transform 1 0 19320 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_209
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_243
timestamp 1688980957
transform 1 0 23460 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_268
timestamp 1688980957
transform 1 0 25760 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_276
timestamp 1688980957
transform 1 0 26496 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_333
timestamp 1688980957
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_350
timestamp 1688980957
transform 1 0 33304 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_356
timestamp 1688980957
transform 1 0 33856 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_364
timestamp 1688980957
transform 1 0 34592 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_372
timestamp 1688980957
transform 1 0 35328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_380
timestamp 1688980957
transform 1 0 36064 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_388
timestamp 1688980957
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_424
timestamp 1688980957
transform 1 0 40112 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_469
timestamp 1688980957
transform 1 0 44252 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_475
timestamp 1688980957
transform 1 0 44804 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_6
timestamp 1688980957
transform 1 0 1656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_12
timestamp 1688980957
transform 1 0 2208 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_23
timestamp 1688980957
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_39
timestamp 1688980957
transform 1 0 4692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_66
timestamp 1688980957
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_73
timestamp 1688980957
transform 1 0 7820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_126
timestamp 1688980957
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_138
timestamp 1688980957
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_152
timestamp 1688980957
transform 1 0 15088 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_164
timestamp 1688980957
transform 1 0 16192 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_176
timestamp 1688980957
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_192
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_216
timestamp 1688980957
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_220
timestamp 1688980957
transform 1 0 21344 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_261
timestamp 1688980957
transform 1 0 25116 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_303
timestamp 1688980957
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_315
timestamp 1688980957
transform 1 0 30084 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_327
timestamp 1688980957
transform 1 0 31188 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_339
timestamp 1688980957
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_343
timestamp 1688980957
transform 1 0 32660 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_350
timestamp 1688980957
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_362
timestamp 1688980957
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_373
timestamp 1688980957
transform 1 0 35420 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_394
timestamp 1688980957
transform 1 0 37352 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_417
timestamp 1688980957
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 1688980957
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 1688980957
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_14
timestamp 1688980957
transform 1 0 2392 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_37
timestamp 1688980957
transform 1 0 4508 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_54
timestamp 1688980957
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_91
timestamp 1688980957
transform 1 0 9476 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_101
timestamp 1688980957
transform 1 0 10396 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_109
timestamp 1688980957
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_117
timestamp 1688980957
transform 1 0 11868 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_159
timestamp 1688980957
transform 1 0 15732 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_164
timestamp 1688980957
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_201
timestamp 1688980957
transform 1 0 19596 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_222
timestamp 1688980957
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_253
timestamp 1688980957
transform 1 0 24380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_269
timestamp 1688980957
transform 1 0 25852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_277
timestamp 1688980957
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_322
timestamp 1688980957
transform 1 0 30728 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_334
timestamp 1688980957
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_341
timestamp 1688980957
transform 1 0 32476 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_346
timestamp 1688980957
transform 1 0 32936 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_358
timestamp 1688980957
transform 1 0 34040 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_370
timestamp 1688980957
transform 1 0 35144 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_382
timestamp 1688980957
transform 1 0 36248 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_390
timestamp 1688980957
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_401
timestamp 1688980957
transform 1 0 37996 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_428
timestamp 1688980957
transform 1 0 40480 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 1688980957
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_473
timestamp 1688980957
transform 1 0 44620 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_21
timestamp 1688980957
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_59
timestamp 1688980957
transform 1 0 6532 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_111
timestamp 1688980957
transform 1 0 11316 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_123
timestamp 1688980957
transform 1 0 12420 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_135
timestamp 1688980957
transform 1 0 13524 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_157
timestamp 1688980957
transform 1 0 15548 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_174
timestamp 1688980957
transform 1 0 17112 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_193
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_205
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_229
timestamp 1688980957
transform 1 0 22172 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_267
timestamp 1688980957
transform 1 0 25668 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_275
timestamp 1688980957
transform 1 0 26404 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_287
timestamp 1688980957
transform 1 0 27508 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_299
timestamp 1688980957
transform 1 0 28612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_329
timestamp 1688980957
transform 1 0 31372 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_341
timestamp 1688980957
transform 1 0 32476 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_359
timestamp 1688980957
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_376
timestamp 1688980957
transform 1 0 35696 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_447
timestamp 1688980957
transform 1 0 42228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_459
timestamp 1688980957
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_471
timestamp 1688980957
transform 1 0 44436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 1688980957
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_41
timestamp 1688980957
transform 1 0 4876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_53
timestamp 1688980957
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_65
timestamp 1688980957
transform 1 0 7084 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_71
timestamp 1688980957
transform 1 0 7636 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_86
timestamp 1688980957
transform 1 0 9016 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_98
timestamp 1688980957
transform 1 0 10120 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_110
timestamp 1688980957
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_145
timestamp 1688980957
transform 1 0 14444 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_166
timestamp 1688980957
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_178
timestamp 1688980957
transform 1 0 17480 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_221
timestamp 1688980957
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_246
timestamp 1688980957
transform 1 0 23736 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_297
timestamp 1688980957
transform 1 0 28428 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_322
timestamp 1688980957
transform 1 0 30728 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_328
timestamp 1688980957
transform 1 0 31280 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_334
timestamp 1688980957
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_363
timestamp 1688980957
transform 1 0 34500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_377
timestamp 1688980957
transform 1 0 35788 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_388
timestamp 1688980957
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_421
timestamp 1688980957
transform 1 0 39836 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_442
timestamp 1688980957
transform 1 0 41768 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 1688980957
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_473
timestamp 1688980957
transform 1 0 44620 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_23
timestamp 1688980957
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_49
timestamp 1688980957
transform 1 0 5612 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_61
timestamp 1688980957
transform 1 0 6716 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_79
timestamp 1688980957
transform 1 0 8372 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_98
timestamp 1688980957
transform 1 0 10120 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_149
timestamp 1688980957
transform 1 0 14812 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_171
timestamp 1688980957
transform 1 0 16836 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_182
timestamp 1688980957
transform 1 0 17848 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_194
timestamp 1688980957
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_237
timestamp 1688980957
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_249
timestamp 1688980957
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_296
timestamp 1688980957
transform 1 0 28336 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_318
timestamp 1688980957
transform 1 0 30360 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_339
timestamp 1688980957
transform 1 0 32292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_351
timestamp 1688980957
transform 1 0 33396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_373
timestamp 1688980957
transform 1 0 35420 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_402
timestamp 1688980957
transform 1 0 38088 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_410
timestamp 1688980957
transform 1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_449
timestamp 1688980957
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_461
timestamp 1688980957
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_473
timestamp 1688980957
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_85
timestamp 1688980957
transform 1 0 8924 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_109
timestamp 1688980957
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_117
timestamp 1688980957
transform 1 0 11868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_155
timestamp 1688980957
transform 1 0 15364 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_159
timestamp 1688980957
transform 1 0 15732 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_180
timestamp 1688980957
transform 1 0 17664 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_186
timestamp 1688980957
transform 1 0 18216 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_212
timestamp 1688980957
transform 1 0 20608 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1688980957
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_233
timestamp 1688980957
transform 1 0 22540 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_254
timestamp 1688980957
transform 1 0 24472 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_266
timestamp 1688980957
transform 1 0 25576 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_274
timestamp 1688980957
transform 1 0 26312 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_294
timestamp 1688980957
transform 1 0 28152 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_306
timestamp 1688980957
transform 1 0 29256 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_318
timestamp 1688980957
transform 1 0 30360 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_330
timestamp 1688980957
transform 1 0 31464 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_349
timestamp 1688980957
transform 1 0 33212 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_363
timestamp 1688980957
transform 1 0 34500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_372
timestamp 1688980957
transform 1 0 35328 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_384
timestamp 1688980957
transform 1 0 36432 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_409
timestamp 1688980957
transform 1 0 38732 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_430
timestamp 1688980957
transform 1 0 40664 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_442
timestamp 1688980957
transform 1 0 41768 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 1688980957
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_473
timestamp 1688980957
transform 1 0 44620 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_25
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_48
timestamp 1688980957
transform 1 0 5520 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_105
timestamp 1688980957
transform 1 0 10764 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_112
timestamp 1688980957
transform 1 0 11408 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_129
timestamp 1688980957
transform 1 0 12972 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_205
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_215
timestamp 1688980957
transform 1 0 20884 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_227
timestamp 1688980957
transform 1 0 21988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_239
timestamp 1688980957
transform 1 0 23092 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1688980957
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_277
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_281
timestamp 1688980957
transform 1 0 26956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_288
timestamp 1688980957
transform 1 0 27600 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_300
timestamp 1688980957
transform 1 0 28704 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_398
timestamp 1688980957
transform 1 0 37720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_410
timestamp 1688980957
transform 1 0 38824 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_418
timestamp 1688980957
transform 1 0 39560 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1688980957
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 1688980957
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 1688980957
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 1688980957
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_50
timestamp 1688980957
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_77
timestamp 1688980957
transform 1 0 8188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_85
timestamp 1688980957
transform 1 0 8924 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_95
timestamp 1688980957
transform 1 0 9844 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_101
timestamp 1688980957
transform 1 0 10396 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_122
timestamp 1688980957
transform 1 0 12328 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_128
timestamp 1688980957
transform 1 0 12880 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_135
timestamp 1688980957
transform 1 0 13524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_154
timestamp 1688980957
transform 1 0 15272 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_164
timestamp 1688980957
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_189
timestamp 1688980957
transform 1 0 18492 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_196
timestamp 1688980957
transform 1 0 19136 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_220
timestamp 1688980957
transform 1 0 21344 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_239
timestamp 1688980957
transform 1 0 23092 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_306
timestamp 1688980957
transform 1 0 29256 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_314
timestamp 1688980957
transform 1 0 29992 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_334
timestamp 1688980957
transform 1 0 31832 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_343
timestamp 1688980957
transform 1 0 32660 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_351
timestamp 1688980957
transform 1 0 33396 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_365
timestamp 1688980957
transform 1 0 34684 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_377
timestamp 1688980957
transform 1 0 35788 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_389
timestamp 1688980957
transform 1 0 36892 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1688980957
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 1688980957
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_473
timestamp 1688980957
transform 1 0 44620 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_7
timestamp 1688980957
transform 1 0 1748 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_34
timestamp 1688980957
transform 1 0 4232 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_43
timestamp 1688980957
transform 1 0 5060 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_59
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_67
timestamp 1688980957
transform 1 0 7268 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_73
timestamp 1688980957
transform 1 0 7820 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_81
timestamp 1688980957
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_94
timestamp 1688980957
transform 1 0 9752 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_122
timestamp 1688980957
transform 1 0 12328 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_185
timestamp 1688980957
transform 1 0 18124 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_213
timestamp 1688980957
transform 1 0 20700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_217
timestamp 1688980957
transform 1 0 21068 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_243
timestamp 1688980957
transform 1 0 23460 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1688980957
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_260
timestamp 1688980957
transform 1 0 25024 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_272
timestamp 1688980957
transform 1 0 26128 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_278
timestamp 1688980957
transform 1 0 26680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_287
timestamp 1688980957
transform 1 0 27508 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_298
timestamp 1688980957
transform 1 0 28520 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_306
timestamp 1688980957
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_317
timestamp 1688980957
transform 1 0 30268 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_348
timestamp 1688980957
transform 1 0 33120 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_368
timestamp 1688980957
transform 1 0 34960 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_372
timestamp 1688980957
transform 1 0 35328 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_379
timestamp 1688980957
transform 1 0 35972 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_391
timestamp 1688980957
transform 1 0 37076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_403
timestamp 1688980957
transform 1 0 38180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_415
timestamp 1688980957
transform 1 0 39284 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1688980957
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 1688980957
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 1688980957
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 1688980957
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_65
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_110
timestamp 1688980957
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_162
timestamp 1688980957
transform 1 0 16008 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_177
timestamp 1688980957
transform 1 0 17388 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_216
timestamp 1688980957
transform 1 0 20976 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_255
timestamp 1688980957
transform 1 0 24564 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_265
timestamp 1688980957
transform 1 0 25484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1688980957
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_340
timestamp 1688980957
transform 1 0 32384 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_348
timestamp 1688980957
transform 1 0 33120 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_369
timestamp 1688980957
transform 1 0 35052 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_381
timestamp 1688980957
transform 1 0 36156 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_389
timestamp 1688980957
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1688980957
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 1688980957
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 1688980957
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 1688980957
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 1688980957
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_473
timestamp 1688980957
transform 1 0 44620 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_35
timestamp 1688980957
transform 1 0 4324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_39
timestamp 1688980957
transform 1 0 4692 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_48
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_75
timestamp 1688980957
transform 1 0 8004 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_193
timestamp 1688980957
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_206
timestamp 1688980957
transform 1 0 20056 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_218
timestamp 1688980957
transform 1 0 21160 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_239
timestamp 1688980957
transform 1 0 23092 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_248
timestamp 1688980957
transform 1 0 23920 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_293
timestamp 1688980957
transform 1 0 28060 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_305
timestamp 1688980957
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_309
timestamp 1688980957
transform 1 0 29532 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_325
timestamp 1688980957
transform 1 0 31004 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_337
timestamp 1688980957
transform 1 0 32108 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_343
timestamp 1688980957
transform 1 0 32660 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_360
timestamp 1688980957
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_373
timestamp 1688980957
transform 1 0 35420 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_385
timestamp 1688980957
transform 1 0 36524 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_397
timestamp 1688980957
transform 1 0 37628 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_409
timestamp 1688980957
transform 1 0 38732 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_417
timestamp 1688980957
transform 1 0 39468 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 1688980957
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 1688980957
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 1688980957
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 1688980957
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 1688980957
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 1688980957
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_61
timestamp 1688980957
transform 1 0 6716 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_84
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_90
timestamp 1688980957
transform 1 0 9384 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_99
timestamp 1688980957
transform 1 0 10212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_134
timestamp 1688980957
transform 1 0 13432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_146
timestamp 1688980957
transform 1 0 14536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_158
timestamp 1688980957
transform 1 0 15640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_166
timestamp 1688980957
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_177
timestamp 1688980957
transform 1 0 17388 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_189
timestamp 1688980957
transform 1 0 18492 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_193
timestamp 1688980957
transform 1 0 18860 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_214
timestamp 1688980957
transform 1 0 20792 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_222
timestamp 1688980957
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1688980957
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1688980957
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1688980957
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_281
timestamp 1688980957
transform 1 0 26956 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_287
timestamp 1688980957
transform 1 0 27508 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_299
timestamp 1688980957
transform 1 0 28612 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_311
timestamp 1688980957
transform 1 0 29716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_323
timestamp 1688980957
transform 1 0 30820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1688980957
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_381
timestamp 1688980957
transform 1 0 36156 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_389
timestamp 1688980957
transform 1 0 36892 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1688980957
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1688980957
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1688980957
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 1688980957
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 1688980957
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 1688980957
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1688980957
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 1688980957
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_473
timestamp 1688980957
transform 1 0 44620 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_61
timestamp 1688980957
transform 1 0 6716 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_70
timestamp 1688980957
transform 1 0 7544 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_82
timestamp 1688980957
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_93
timestamp 1688980957
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_119
timestamp 1688980957
transform 1 0 12052 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_131
timestamp 1688980957
transform 1 0 13156 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_156
timestamp 1688980957
transform 1 0 15456 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_162
timestamp 1688980957
transform 1 0 16008 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_174
timestamp 1688980957
transform 1 0 17112 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_186
timestamp 1688980957
transform 1 0 18216 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_206
timestamp 1688980957
transform 1 0 20056 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_218
timestamp 1688980957
transform 1 0 21160 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_226
timestamp 1688980957
transform 1 0 21896 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_232
timestamp 1688980957
transform 1 0 22448 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_248
timestamp 1688980957
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_261
timestamp 1688980957
transform 1 0 25116 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_265
timestamp 1688980957
transform 1 0 25484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_269
timestamp 1688980957
transform 1 0 25852 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_290
timestamp 1688980957
transform 1 0 27784 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_302
timestamp 1688980957
transform 1 0 28888 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_309
timestamp 1688980957
transform 1 0 29532 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1688980957
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1688980957
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1688980957
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1688980957
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1688980957
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1688980957
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1688980957
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1688980957
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1688980957
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1688980957
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1688980957
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 1688980957
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 1688980957
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 1688980957
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_77
timestamp 1688980957
transform 1 0 8188 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_149
timestamp 1688980957
transform 1 0 14812 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_178
timestamp 1688980957
transform 1 0 17480 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_211
timestamp 1688980957
transform 1 0 20516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1688980957
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_245
timestamp 1688980957
transform 1 0 23644 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_249
timestamp 1688980957
transform 1 0 24012 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_272
timestamp 1688980957
transform 1 0 26128 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_301
timestamp 1688980957
transform 1 0 28796 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_313
timestamp 1688980957
transform 1 0 29900 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_325
timestamp 1688980957
transform 1 0 31004 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_333
timestamp 1688980957
transform 1 0 31740 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1688980957
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1688980957
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1688980957
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1688980957
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1688980957
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1688980957
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1688980957
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1688980957
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1688980957
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1688980957
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 1688980957
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 1688980957
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1688980957
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_461
timestamp 1688980957
transform 1 0 43516 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_469
timestamp 1688980957
transform 1 0 44252 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_105
timestamp 1688980957
transform 1 0 10764 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_153
timestamp 1688980957
transform 1 0 15180 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1688980957
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_209
timestamp 1688980957
transform 1 0 20332 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_217
timestamp 1688980957
transform 1 0 21068 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1688980957
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1688980957
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1688980957
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1688980957
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 1688980957
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 1688980957
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1688980957
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1688980957
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1688980957
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1688980957
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1688980957
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1688980957
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1688980957
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1688980957
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1688980957
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1688980957
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 1688980957
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 1688980957
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1688980957
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1688980957
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_104
timestamp 1688980957
transform 1 0 10672 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_116
timestamp 1688980957
transform 1 0 11776 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_128
timestamp 1688980957
transform 1 0 12880 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_165
timestamp 1688980957
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_189
timestamp 1688980957
transform 1 0 18492 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_201
timestamp 1688980957
transform 1 0 19596 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_213
timestamp 1688980957
transform 1 0 20700 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_221
timestamp 1688980957
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_225
timestamp 1688980957
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_235
timestamp 1688980957
transform 1 0 22724 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_245
timestamp 1688980957
transform 1 0 23644 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_252
timestamp 1688980957
transform 1 0 24288 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_256
timestamp 1688980957
transform 1 0 24656 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_267
timestamp 1688980957
transform 1 0 25668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1688980957
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_322
timestamp 1688980957
transform 1 0 30728 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_334
timestamp 1688980957
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1688980957
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1688980957
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1688980957
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1688980957
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1688980957
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1688980957
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1688980957
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1688980957
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1688980957
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 1688980957
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 1688980957
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 1688980957
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1688980957
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 1688980957
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_473
timestamp 1688980957
transform 1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_13
timestamp 1688980957
transform 1 0 2300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_25
timestamp 1688980957
transform 1 0 3404 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_57
timestamp 1688980957
transform 1 0 6348 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_63
timestamp 1688980957
transform 1 0 6900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_75
timestamp 1688980957
transform 1 0 8004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1688980957
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_109
timestamp 1688980957
transform 1 0 11132 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_113
timestamp 1688980957
transform 1 0 11500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_125
timestamp 1688980957
transform 1 0 12604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_137
timestamp 1688980957
transform 1 0 13708 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_141
timestamp 1688980957
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1688980957
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_165
timestamp 1688980957
transform 1 0 16284 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_169
timestamp 1688980957
transform 1 0 16652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_181
timestamp 1688980957
transform 1 0 17756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_193
timestamp 1688980957
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1688980957
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1688980957
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_221
timestamp 1688980957
transform 1 0 21436 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_232
timestamp 1688980957
transform 1 0 22448 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_244
timestamp 1688980957
transform 1 0 23552 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1688980957
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1688980957
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1688980957
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_277
timestamp 1688980957
transform 1 0 26588 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_281
timestamp 1688980957
transform 1 0 26956 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_285
timestamp 1688980957
transform 1 0 27324 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_289
timestamp 1688980957
transform 1 0 27692 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_293
timestamp 1688980957
transform 1 0 28060 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_297
timestamp 1688980957
transform 1 0 28428 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_305
timestamp 1688980957
transform 1 0 29164 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1688980957
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1688980957
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_333
timestamp 1688980957
transform 1 0 31740 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_337
timestamp 1688980957
transform 1 0 32108 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_345
timestamp 1688980957
transform 1 0 32844 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_349
timestamp 1688980957
transform 1 0 33212 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_361
timestamp 1688980957
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1688980957
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1688980957
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_389
timestamp 1688980957
transform 1 0 36892 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_393
timestamp 1688980957
transform 1 0 37260 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_405
timestamp 1688980957
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_417
timestamp 1688980957
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 1688980957
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_433
timestamp 1688980957
transform 1 0 40940 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_441
timestamp 1688980957
transform 1 0 41676 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_449
timestamp 1688980957
transform 1 0 42412 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_461
timestamp 1688980957
transform 1 0 43516 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_473
timestamp 1688980957
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 35604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 10948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 29072 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 43148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 11684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 31556 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 4508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 41308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 21896 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 1840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 27784 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 37996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 8556 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold35
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 43976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 19596 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 20148 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 35604 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 37996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 40388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 40480 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 16928 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 19044 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold45
timestamp 1688980957
transform -1 0 28428 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 13432 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 15548 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 14812 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 43240 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 41676 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 8188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 17388 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 16100 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 28796 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 27692 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 30728 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 39376 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 9660 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 7636 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 5336 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 4784 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 20884 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 41032 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 5428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 4784 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 32844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 5704 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 6808 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 36432 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 35880 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 23184 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 23460 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 31004 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 5520 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 3588 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 25116 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 23736 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 40572 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 38824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 29532 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 23644 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 21988 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 41400 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 24840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 3772 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 39376 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 38548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 12696 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 12972 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 10212 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 8096 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 36156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 25116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold102
timestamp 1688980957
transform -1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 34040 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 20700 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 19320 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 33120 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 27692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 43884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 42136 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform 1 0 32660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 43148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 43884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 36892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 31372 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 38732 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 37444 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 33580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 33948 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 36892 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 37260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 37996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 36248 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform 1 0 23184 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 32660 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 35420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 40572 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 38916 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 33580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 14904 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 41768 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 21620 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 20608 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 38180 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 33028 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 19136 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 35420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 26312 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform -1 0 42320 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 39468 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform -1 0 35420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 35696 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 44620 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 37076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform -1 0 23736 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 8832 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 9384 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 18216 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 3404 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 42228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 27692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 39008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 39836 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 40020 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform -1 0 14168 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 38456 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform 1 0 21896 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 44712 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 43884 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform -1 0 26220 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform -1 0 9660 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 34224 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 23000 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 40296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 4140 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 3220 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 20516 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform 1 0 9936 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 10028 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform -1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 41768 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 25944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 15456 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform -1 0 18216 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform -1 0 17848 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 18860 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 5704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 12604 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 24380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform -1 0 17848 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 42412 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform -1 0 19136 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 9844 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform -1 0 36800 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 15364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 4048 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 35236 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 37996 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 19964 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 28520 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform 1 0 27140 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 26128 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 43056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform -1 0 25116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform -1 0 23092 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 3128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 22540 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform -1 0 13616 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 30452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 13800 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold221
timestamp 1688980957
transform -1 0 18216 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform -1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 19872 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 18768 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform -1 0 35420 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 7728 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform -1 0 32108 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform 1 0 37536 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 39008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 21252 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 35144 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 42228 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 16560 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 19964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform 1 0 25208 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 37996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform 1 0 19228 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 36432 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform 1 0 33488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform 1 0 23092 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 26404 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform -1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 23644 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 9844 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 39284 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 5060 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 23736 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 36616 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 26404 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform -1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform -1 0 22264 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 21528 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform 1 0 26404 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform -1 0 42044 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform -1 0 23368 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform -1 0 44896 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform -1 0 42320 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 24196 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 44620 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 14904 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 44896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 33212 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 26772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1688980957
transform 1 0 6532 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1688980957
transform 1 0 44528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45172 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45172 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45172 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45172 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45172 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45172 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45172 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 45172 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 45172 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 45172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 45172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 45172 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 45172 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 45172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 45172 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 45172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 45172 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 45172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 45172 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 45172 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 45172 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 45172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 45172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 45172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 45172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 45172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 45172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 45172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 45172 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 45172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 45172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 45172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 45172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 45172 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 45172 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 45172 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 45172 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 45172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 45172 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 45172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 45172 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 45172 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 45172 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 45172 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 45172 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 45172 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 45172 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 45172 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 45172 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 45172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 45172 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 45172 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 45172 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 45172 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 45172 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 45172 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 45172 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 45172 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 45172 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 45172 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 45172 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 45172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 45172 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 45172 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 45172 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 45172 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 45172 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 45172 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 45172 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 45172 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 45172 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 45172 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 45172 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 45172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1688980957
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1688980957
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1688980957
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1688980957
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1688980957
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1688980957
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1688980957
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1688980957
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1688980957
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1688980957
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1688980957
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1688980957
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1688980957
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1688980957
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1688980957
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1688980957
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1688980957
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1688980957
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1688980957
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1688980957
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1688980957
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1688980957
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1688980957
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1688980957
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1688980957
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1688980957
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1688980957
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1688980957
transform 1 0 6256 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1688980957
transform 1 0 11408 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1688980957
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1688980957
transform 1 0 16560 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1688980957
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1688980957
transform 1 0 21712 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1688980957
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1688980957
transform 1 0 26864 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1688980957
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1688980957
transform 1 0 32016 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1688980957
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1688980957
transform 1 0 37168 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1688980957
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1688980957
transform 1 0 42320 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  wire21
timestamp 1688980957
transform 1 0 23736 0 1 32640
box -38 -48 590 592
<< labels >>
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 45537 44208 46337 44328 0 FreeSans 480 0 0 0 cs
port 1 nsew signal input
flabel metal2 s 41878 47681 41934 48481 0 FreeSans 224 90 0 0 gpio[0]
port 2 nsew signal input
flabel metal2 s 23846 47681 23902 48481 0 FreeSans 224 90 0 0 gpio[10]
port 3 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpio[11]
port 4 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpio[12]
port 5 nsew signal input
flabel metal3 s 45537 6808 46337 6928 0 FreeSans 480 0 0 0 gpio[13]
port 6 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 gpio[14]
port 7 nsew signal input
flabel metal3 s 45537 34688 46337 34808 0 FreeSans 480 0 0 0 gpio[15]
port 8 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio[16]
port 9 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio[1]
port 10 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 gpio[2]
port 11 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio[3]
port 12 nsew signal input
flabel metal2 s 14830 47681 14886 48481 0 FreeSans 224 90 0 0 gpio[4]
port 13 nsew signal input
flabel metal3 s 45537 25168 46337 25288 0 FreeSans 480 0 0 0 gpio[5]
port 14 nsew signal input
flabel metal3 s 0 46248 800 46368 0 FreeSans 480 0 0 0 gpio[6]
port 15 nsew signal input
flabel metal2 s 32862 47681 32918 48481 0 FreeSans 224 90 0 0 gpio[7]
port 16 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 gpio[8]
port 17 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 gpio[9]
port 18 nsew signal input
flabel metal2 s 6458 47681 6514 48481 0 FreeSans 224 90 0 0 nrst
port 19 nsew signal input
flabel metal3 s 45537 16328 46337 16448 0 FreeSans 480 0 0 0 pwm
port 20 nsew signal tristate
flabel metal4 s 4208 2128 4528 46288 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 34928 2128 35248 46288 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 19568 2128 19888 46288 0 FreeSans 1920 90 0 0 vssd1
port 22 nsew ground bidirectional
rlabel metal1 23138 46240 23138 46240 0 vccd1
rlabel metal1 23138 45696 23138 45696 0 vssd1
rlabel metal1 25254 22984 25254 22984 0 _0000_
rlabel metal1 23644 21862 23644 21862 0 _0001_
rlabel metal1 24518 20570 24518 20570 0 _0002_
rlabel metal2 26174 21794 26174 21794 0 _0003_
rlabel metal1 26312 17714 26312 17714 0 _0004_
rlabel metal1 23782 18190 23782 18190 0 _0005_
rlabel metal1 23966 19278 23966 19278 0 _0006_
rlabel metal1 27232 19414 27232 19414 0 _0007_
rlabel metal1 25070 24854 25070 24854 0 _0008_
rlabel metal1 23828 25330 23828 25330 0 _0009_
rlabel metal1 27048 25942 27048 25942 0 _0010_
rlabel metal1 24472 26418 24472 26418 0 _0011_
rlabel metal1 26808 27642 26808 27642 0 _0012_
rlabel metal1 27048 29206 27048 29206 0 _0013_
rlabel metal1 27324 30294 27324 30294 0 _0014_
rlabel metal1 27186 31858 27186 31858 0 _0015_
rlabel metal1 26450 32810 26450 32810 0 _0016_
rlabel metal1 28014 33422 28014 33422 0 _0017_
rlabel metal1 24472 3434 24472 3434 0 _0018_
rlabel metal1 22724 4658 22724 4658 0 _0019_
rlabel metal1 25520 5882 25520 5882 0 _0020_
rlabel metal1 27416 23290 27416 23290 0 _0021_
rlabel metal1 32614 22542 32614 22542 0 _0022_
rlabel via1 36287 22202 36287 22202 0 _0023_
rlabel metal1 35650 23834 35650 23834 0 _0024_
rlabel metal1 37444 18666 37444 18666 0 _0025_
rlabel metal1 33994 17714 33994 17714 0 _0026_
rlabel metal2 32430 18156 32430 18156 0 _0027_
rlabel metal1 33948 23154 33948 23154 0 _0028_
rlabel metal1 31096 26010 31096 26010 0 _0029_
rlabel metal1 34270 25364 34270 25364 0 _0030_
rlabel metal1 36202 27098 36202 27098 0 _0031_
rlabel metal1 35558 29274 35558 29274 0 _0032_
rlabel metal1 32890 28458 32890 28458 0 _0033_
rlabel metal1 34270 31382 34270 31382 0 _0034_
rlabel metal1 31004 33082 31004 33082 0 _0035_
rlabel metal1 34592 33082 34592 33082 0 _0036_
rlabel metal1 31832 36210 31832 36210 0 _0037_
rlabel metal1 35374 36210 35374 36210 0 _0038_
rlabel metal1 36202 39508 36202 39508 0 _0039_
rlabel metal1 35834 40596 35834 40596 0 _0040_
rlabel metal1 34132 42330 34132 42330 0 _0041_
rlabel metal1 32936 42874 32936 42874 0 _0042_
rlabel metal1 30912 41786 30912 41786 0 _0043_
rlabel metal1 29348 41786 29348 41786 0 _0044_
rlabel metal1 28474 37944 28474 37944 0 _0045_
rlabel metal1 28375 36346 28375 36346 0 _0046_
rlabel metal1 35972 36890 35972 36890 0 _0047_
rlabel metal1 37398 38250 37398 38250 0 _0048_
rlabel metal2 40066 38828 40066 38828 0 _0049_
rlabel metal1 39974 37978 39974 37978 0 _0050_
rlabel metal2 39146 39236 39146 39236 0 _0051_
rlabel metal1 39744 36822 39744 36822 0 _0052_
rlabel metal1 39008 36210 39008 36210 0 _0053_
rlabel metal1 36156 34578 36156 34578 0 _0054_
rlabel metal1 24886 36890 24886 36890 0 _0055_
rlabel metal1 23414 37978 23414 37978 0 _0056_
rlabel metal1 21482 38862 21482 38862 0 _0057_
rlabel metal2 20194 39780 20194 39780 0 _0058_
rlabel metal1 17112 40154 17112 40154 0 _0059_
rlabel metal1 12834 40596 12834 40596 0 _0060_
rlabel metal1 8188 40154 8188 40154 0 _0061_
rlabel metal1 7636 39406 7636 39406 0 _0062_
rlabel metal1 4416 39066 4416 39066 0 _0063_
rlabel metal2 3542 40426 3542 40426 0 _0064_
rlabel metal1 3726 41004 3726 41004 0 _0065_
rlabel metal1 4968 41786 4968 41786 0 _0066_
rlabel metal1 6992 42330 6992 42330 0 _0067_
rlabel metal2 8142 42908 8142 42908 0 _0068_
rlabel metal2 12834 42228 12834 42228 0 _0069_
rlabel metal1 14398 40970 14398 40970 0 _0070_
rlabel metal2 16698 43044 16698 43044 0 _0071_
rlabel metal1 19320 41786 19320 41786 0 _0072_
rlabel metal1 27002 34578 27002 34578 0 _0073_
rlabel metal1 24702 42568 24702 42568 0 _0074_
rlabel metal1 27048 41786 27048 41786 0 _0075_
rlabel metal1 25300 40698 25300 40698 0 _0076_
rlabel metal2 26818 39916 26818 39916 0 _0077_
rlabel metal1 24797 39066 24797 39066 0 _0078_
rlabel metal1 35880 31926 35880 31926 0 _0079_
rlabel metal1 43102 34680 43102 34680 0 _0080_
rlabel metal1 42918 31858 42918 31858 0 _0081_
rlabel metal1 43240 33626 43240 33626 0 _0082_
rlabel metal1 40526 32470 40526 32470 0 _0083_
rlabel metal1 39928 32946 39928 32946 0 _0084_
rlabel metal1 38134 31654 38134 31654 0 _0085_
rlabel metal1 37536 29206 37536 29206 0 _0086_
rlabel metal1 36340 33966 36340 33966 0 _0087_
rlabel metal1 41492 34714 41492 34714 0 _0088_
rlabel metal1 42320 37774 42320 37774 0 _0089_
rlabel metal1 41952 36210 41952 36210 0 _0090_
rlabel metal1 41032 36686 41032 36686 0 _0091_
rlabel metal1 41262 33388 41262 33388 0 _0092_
rlabel metal1 38456 34714 38456 34714 0 _0093_
rlabel metal2 37122 33796 37122 33796 0 _0094_
rlabel metal2 17618 23970 17618 23970 0 _0095_
rlabel metal2 17894 22882 17894 22882 0 _0096_
rlabel metal2 17802 20706 17802 20706 0 _0097_
rlabel metal2 15778 21794 15778 21794 0 _0098_
rlabel via1 15957 18734 15957 18734 0 _0099_
rlabel metal2 14122 19142 14122 19142 0 _0100_
rlabel metal2 12466 19618 12466 19618 0 _0101_
rlabel metal2 10718 19618 10718 19618 0 _0102_
rlabel metal1 12665 23018 12665 23018 0 _0103_
rlabel metal1 15088 24378 15088 24378 0 _0104_
rlabel metal1 11863 22678 11863 22678 0 _0105_
rlabel metal2 10902 25058 10902 25058 0 _0106_
rlabel metal1 12926 25466 12926 25466 0 _0107_
rlabel via1 20281 28050 20281 28050 0 _0108_
rlabel via1 22116 29206 22116 29206 0 _0109_
rlabel metal1 24748 31654 24748 31654 0 _0110_
rlabel metal2 26358 31178 26358 31178 0 _0111_
rlabel metal2 22586 31144 22586 31144 0 _0112_
rlabel metal2 19090 21794 19090 21794 0 _0113_
rlabel metal1 22024 21522 22024 21522 0 _0114_
rlabel metal1 18671 19414 18671 19414 0 _0115_
rlabel metal1 21098 20842 21098 20842 0 _0116_
rlabel metal2 20654 18530 20654 18530 0 _0117_
rlabel metal1 22576 18258 22576 18258 0 _0118_
rlabel metal1 19412 18394 19412 18394 0 _0119_
rlabel metal1 21505 19482 21505 19482 0 _0120_
rlabel metal1 22816 22746 22816 22746 0 _0121_
rlabel metal1 19872 23290 19872 23290 0 _0122_
rlabel metal1 21098 23018 21098 23018 0 _0123_
rlabel metal1 19724 25262 19724 25262 0 _0124_
rlabel metal1 19913 25942 19913 25942 0 _0125_
rlabel metal2 21666 26146 21666 26146 0 _0126_
rlabel metal1 23736 28186 23736 28186 0 _0127_
rlabel metal1 24600 26962 24600 26962 0 _0128_
rlabel metal2 25438 28322 25438 28322 0 _0129_
rlabel metal1 21758 27472 21758 27472 0 _0130_
rlabel metal1 15863 25466 15863 25466 0 _0131_
rlabel metal1 17664 24922 17664 24922 0 _0132_
rlabel metal1 17158 26010 17158 26010 0 _0133_
rlabel metal1 14996 22746 14996 22746 0 _0134_
rlabel metal1 15456 19754 15456 19754 0 _0135_
rlabel metal1 13248 21862 13248 21862 0 _0136_
rlabel metal1 12190 20298 12190 20298 0 _0137_
rlabel metal1 9936 20570 9936 20570 0 _0138_
rlabel metal1 9936 23154 9936 23154 0 _0139_
rlabel metal1 13478 24718 13478 24718 0 _0140_
rlabel metal1 8648 22542 8648 22542 0 _0141_
rlabel metal1 9798 25466 9798 25466 0 _0142_
rlabel metal1 8004 25466 8004 25466 0 _0143_
rlabel metal1 19504 30294 19504 30294 0 _0144_
rlabel metal1 20148 31654 20148 31654 0 _0145_
rlabel metal1 23046 32470 23046 32470 0 _0146_
rlabel metal1 25898 33592 25898 33592 0 _0147_
rlabel metal2 22126 31518 22126 31518 0 _0148_
rlabel metal1 24042 35734 24042 35734 0 _0149_
rlabel metal1 21873 34714 21873 34714 0 _0150_
rlabel metal1 19626 36074 19626 36074 0 _0151_
rlabel metal2 17710 37638 17710 37638 0 _0152_
rlabel metal2 15962 38114 15962 38114 0 _0153_
rlabel metal2 14214 39202 14214 39202 0 _0154_
rlabel metal1 7482 38250 7482 38250 0 _0155_
rlabel via1 7401 33966 7401 33966 0 _0156_
rlabel metal2 2162 34850 2162 34850 0 _0157_
rlabel via1 1789 32470 1789 32470 0 _0158_
rlabel metal1 5193 32810 5193 32810 0 _0159_
rlabel metal2 2162 38114 2162 38114 0 _0160_
rlabel metal1 5014 37434 5014 37434 0 _0161_
rlabel via1 8597 44370 8597 44370 0 _0162_
rlabel metal1 12466 43724 12466 43724 0 _0163_
rlabel metal1 13616 45050 13616 45050 0 _0164_
rlabel metal1 15594 43962 15594 43962 0 _0165_
rlabel metal1 18430 44438 18430 44438 0 _0166_
rlabel metal2 23046 36550 23046 36550 0 _0167_
rlabel metal2 20838 37026 20838 37026 0 _0168_
rlabel metal1 19626 37162 19626 37162 0 _0169_
rlabel metal2 18630 38726 18630 38726 0 _0170_
rlabel metal1 15486 39338 15486 39338 0 _0171_
rlabel metal2 11546 39202 11546 39202 0 _0172_
rlabel metal1 7544 37434 7544 37434 0 _0173_
rlabel metal2 7222 32674 7222 32674 0 _0174_
rlabel metal1 3404 35258 3404 35258 0 _0175_
rlabel metal1 3189 33558 3189 33558 0 _0176_
rlabel metal2 3910 33762 3910 33762 0 _0177_
rlabel metal1 3256 37842 3256 37842 0 _0178_
rlabel metal1 6992 37434 6992 37434 0 _0179_
rlabel metal2 8326 41990 8326 41990 0 _0180_
rlabel metal1 10483 41514 10483 41514 0 _0181_
rlabel metal1 12875 42262 12875 42262 0 _0182_
rlabel metal1 16130 41514 16130 41514 0 _0183_
rlabel metal1 18349 42194 18349 42194 0 _0184_
rlabel metal1 25076 35258 25076 35258 0 _0185_
rlabel metal1 21160 32810 21160 32810 0 _0186_
rlabel metal1 19596 33898 19596 33898 0 _0187_
rlabel metal1 17710 35768 17710 35768 0 _0188_
rlabel metal1 16744 35530 16744 35530 0 _0189_
rlabel metal1 13892 39950 13892 39950 0 _0190_
rlabel metal1 9614 38250 9614 38250 0 _0191_
rlabel metal1 9016 33898 9016 33898 0 _0192_
rlabel metal1 3082 30906 3082 30906 0 _0193_
rlabel metal1 1840 30770 1840 30770 0 _0194_
rlabel metal1 5704 31858 5704 31858 0 _0195_
rlabel metal1 1886 36822 1886 36822 0 _0196_
rlabel metal1 5060 34986 5060 34986 0 _0197_
rlabel metal1 9144 45050 9144 45050 0 _0198_
rlabel metal1 11447 45050 11447 45050 0 _0199_
rlabel metal2 14490 44642 14490 44642 0 _0200_
rlabel metal2 16238 45084 16238 45084 0 _0201_
rlabel metal1 17933 45050 17933 45050 0 _0202_
rlabel metal1 17020 2890 17020 2890 0 _0203_
rlabel metal1 14904 3366 14904 3366 0 _0204_
rlabel metal1 11822 4658 11822 4658 0 _0205_
rlabel metal1 10672 5338 10672 5338 0 _0206_
rlabel metal1 18676 4182 18676 4182 0 _0207_
rlabel metal1 21252 4794 21252 4794 0 _0208_
rlabel metal1 24978 22746 24978 22746 0 _0209_
rlabel metal1 24104 21862 24104 21862 0 _0210_
rlabel metal1 24196 20434 24196 20434 0 _0211_
rlabel metal1 26680 21522 26680 21522 0 _0212_
rlabel metal2 26174 18428 26174 18428 0 _0213_
rlabel metal1 23230 18836 23230 18836 0 _0214_
rlabel metal1 24012 18938 24012 18938 0 _0215_
rlabel metal1 26818 19278 26818 19278 0 _0216_
rlabel metal1 24794 24378 24794 24378 0 _0217_
rlabel metal1 36662 32232 36662 32232 0 _0218_
rlabel metal1 23506 24922 23506 24922 0 _0219_
rlabel metal1 26680 25466 26680 25466 0 _0220_
rlabel metal1 24150 26010 24150 26010 0 _0221_
rlabel metal1 26726 27098 26726 27098 0 _0222_
rlabel metal1 26680 28730 26680 28730 0 _0223_
rlabel metal2 27186 30260 27186 30260 0 _0224_
rlabel metal1 26956 31450 26956 31450 0 _0225_
rlabel metal1 26542 32538 26542 32538 0 _0226_
rlabel metal1 27968 33082 27968 33082 0 _0227_
rlabel metal1 23690 7378 23690 7378 0 _0228_
rlabel metal1 23506 10642 23506 10642 0 _0229_
rlabel metal1 23230 9554 23230 9554 0 _0230_
rlabel metal1 23506 4998 23506 4998 0 _0231_
rlabel metal1 23966 4590 23966 4590 0 _0232_
rlabel metal1 25898 5134 25898 5134 0 _0233_
rlabel metal1 33994 5882 33994 5882 0 _0234_
rlabel metal1 24840 5202 24840 5202 0 _0235_
rlabel metal1 23782 4726 23782 4726 0 _0236_
rlabel metal1 27278 6732 27278 6732 0 _0237_
rlabel metal1 26220 12818 26220 12818 0 _0238_
rlabel metal2 25530 5338 25530 5338 0 _0239_
rlabel metal1 24978 5168 24978 5168 0 _0240_
rlabel metal1 23966 3604 23966 3604 0 _0241_
rlabel metal1 24794 5576 24794 5576 0 _0242_
rlabel metal1 24380 6426 24380 6426 0 _0243_
rlabel metal1 24334 5746 24334 5746 0 _0244_
rlabel metal1 23506 5168 23506 5168 0 _0245_
rlabel metal1 23460 6766 23460 6766 0 _0246_
rlabel metal1 24242 6630 24242 6630 0 _0247_
rlabel metal1 18538 39984 18538 39984 0 _0248_
rlabel metal1 36616 38250 36616 38250 0 _0249_
rlabel metal1 28060 23086 28060 23086 0 _0250_
rlabel metal2 27738 23562 27738 23562 0 _0251_
rlabel metal1 34615 18666 34615 18666 0 _0252_
rlabel metal1 29210 24820 29210 24820 0 _0253_
rlabel metal2 29762 23018 29762 23018 0 _0254_
rlabel metal2 29118 22644 29118 22644 0 _0255_
rlabel metal1 30590 23052 30590 23052 0 _0256_
rlabel metal1 30314 23188 30314 23188 0 _0257_
rlabel metal1 30774 22746 30774 22746 0 _0258_
rlabel metal2 32154 23494 32154 23494 0 _0259_
rlabel metal1 35696 21590 35696 21590 0 _0260_
rlabel metal1 34500 21998 34500 21998 0 _0261_
rlabel metal1 29624 21522 29624 21522 0 _0262_
rlabel metal1 34132 21998 34132 21998 0 _0263_
rlabel metal1 35190 22032 35190 22032 0 _0264_
rlabel metal1 34730 21964 34730 21964 0 _0265_
rlabel metal1 35834 21386 35834 21386 0 _0266_
rlabel metal1 36202 22678 36202 22678 0 _0267_
rlabel metal2 36110 22134 36110 22134 0 _0268_
rlabel metal1 36340 23630 36340 23630 0 _0269_
rlabel metal1 29210 21454 29210 21454 0 _0270_
rlabel metal1 35282 21454 35282 21454 0 _0271_
rlabel metal1 36294 21556 36294 21556 0 _0272_
rlabel metal1 36064 20842 36064 20842 0 _0273_
rlabel metal1 36432 21658 36432 21658 0 _0274_
rlabel metal1 35834 23732 35834 23732 0 _0275_
rlabel metal1 36064 23698 36064 23698 0 _0276_
rlabel metal2 36432 19346 36432 19346 0 _0277_
rlabel metal2 35374 21828 35374 21828 0 _0278_
rlabel metal1 35926 20434 35926 20434 0 _0279_
rlabel metal2 36846 19788 36846 19788 0 _0280_
rlabel metal2 29026 20604 29026 20604 0 _0281_
rlabel metal1 30551 18734 30551 18734 0 _0282_
rlabel metal1 33580 19142 33580 19142 0 _0283_
rlabel metal1 36984 19346 36984 19346 0 _0284_
rlabel metal1 37030 19414 37030 19414 0 _0285_
rlabel metal1 36294 19278 36294 19278 0 _0286_
rlabel metal1 35696 19346 35696 19346 0 _0287_
rlabel metal2 35558 19652 35558 19652 0 _0288_
rlabel metal1 35282 19346 35282 19346 0 _0289_
rlabel metal2 28658 18598 28658 18598 0 _0290_
rlabel metal1 33396 19822 33396 19822 0 _0291_
rlabel metal1 34776 19482 34776 19482 0 _0292_
rlabel metal1 33994 18632 33994 18632 0 _0293_
rlabel metal1 33902 18768 33902 18768 0 _0294_
rlabel metal1 32614 19346 32614 19346 0 _0295_
rlabel metal1 29026 19176 29026 19176 0 _0296_
rlabel metal1 29946 19278 29946 19278 0 _0297_
rlabel metal1 31050 19278 31050 19278 0 _0298_
rlabel metal1 32016 19822 32016 19822 0 _0299_
rlabel metal1 31096 19482 31096 19482 0 _0300_
rlabel metal1 32936 18734 32936 18734 0 _0301_
rlabel metal1 35742 19754 35742 19754 0 _0302_
rlabel metal1 35420 19890 35420 19890 0 _0303_
rlabel metal2 34914 19618 34914 19618 0 _0304_
rlabel metal1 34592 19822 34592 19822 0 _0305_
rlabel metal1 32522 20468 32522 20468 0 _0306_
rlabel metal1 31970 18802 31970 18802 0 _0307_
rlabel viali 31878 18712 31878 18712 0 _0308_
rlabel metal2 31418 20128 31418 20128 0 _0309_
rlabel metal1 29532 19482 29532 19482 0 _0310_
rlabel metal1 31510 19788 31510 19788 0 _0311_
rlabel metal1 32568 19822 32568 19822 0 _0312_
rlabel metal2 32338 20094 32338 20094 0 _0313_
rlabel metal2 32430 20672 32430 20672 0 _0314_
rlabel metal1 32016 20570 32016 20570 0 _0315_
rlabel metal1 32522 24174 32522 24174 0 _0316_
rlabel metal2 32246 20230 32246 20230 0 _0317_
rlabel metal1 32660 20570 32660 20570 0 _0318_
rlabel metal2 33258 24242 33258 24242 0 _0319_
rlabel metal1 29762 32402 29762 32402 0 _0320_
rlabel metal1 29394 20026 29394 20026 0 _0321_
rlabel metal2 29762 24548 29762 24548 0 _0322_
rlabel metal1 31970 24786 31970 24786 0 _0323_
rlabel metal2 33350 25806 33350 25806 0 _0324_
rlabel metal1 32844 24786 32844 24786 0 _0325_
rlabel metal2 31970 25364 31970 25364 0 _0326_
rlabel metal1 33028 25330 33028 25330 0 _0327_
rlabel metal2 31602 25670 31602 25670 0 _0328_
rlabel metal1 29072 24922 29072 24922 0 _0329_
rlabel metal1 32338 25194 32338 25194 0 _0330_
rlabel metal1 33488 26418 33488 26418 0 _0331_
rlabel metal2 33442 25976 33442 25976 0 _0332_
rlabel metal1 33626 26248 33626 26248 0 _0333_
rlabel metal1 33764 24922 33764 24922 0 _0334_
rlabel metal1 33626 25262 33626 25262 0 _0335_
rlabel metal1 29440 25670 29440 25670 0 _0336_
rlabel metal2 29670 26452 29670 26452 0 _0337_
rlabel metal1 34684 26350 34684 26350 0 _0338_
rlabel metal2 35282 27268 35282 27268 0 _0339_
rlabel metal1 33718 25908 33718 25908 0 _0340_
rlabel metal2 33994 26044 33994 26044 0 _0341_
rlabel metal2 35374 26044 35374 26044 0 _0342_
rlabel metal1 35788 26554 35788 26554 0 _0343_
rlabel metal1 35466 26962 35466 26962 0 _0344_
rlabel metal2 28842 26724 28842 26724 0 _0345_
rlabel viali 30590 26961 30590 26961 0 _0346_
rlabel metal2 35282 27931 35282 27931 0 _0347_
rlabel metal1 35604 27846 35604 27846 0 _0348_
rlabel metal1 35282 28118 35282 28118 0 _0349_
rlabel metal1 36064 27846 36064 27846 0 _0350_
rlabel metal1 35374 28492 35374 28492 0 _0351_
rlabel metal1 34914 26384 34914 26384 0 _0352_
rlabel metal1 34638 27438 34638 27438 0 _0353_
rlabel metal1 34500 27574 34500 27574 0 _0354_
rlabel metal1 34960 28730 34960 28730 0 _0355_
rlabel metal1 34224 29546 34224 29546 0 _0356_
rlabel metal1 30590 29206 30590 29206 0 _0357_
rlabel metal1 30268 29070 30268 29070 0 _0358_
rlabel metal1 33258 29104 33258 29104 0 _0359_
rlabel metal1 33718 30226 33718 30226 0 _0360_
rlabel metal1 33534 29274 33534 29274 0 _0361_
rlabel metal1 33994 29478 33994 29478 0 _0362_
rlabel metal1 34776 27574 34776 27574 0 _0363_
rlabel metal1 34132 30022 34132 30022 0 _0364_
rlabel metal1 33718 28424 33718 28424 0 _0365_
rlabel metal1 33396 28526 33396 28526 0 _0366_
rlabel metal1 32154 29580 32154 29580 0 _0367_
rlabel metal1 29900 29682 29900 29682 0 _0368_
rlabel metal1 31786 29648 31786 29648 0 _0369_
rlabel metal1 32292 29750 32292 29750 0 _0370_
rlabel metal1 32660 29818 32660 29818 0 _0371_
rlabel metal1 32936 30090 32936 30090 0 _0372_
rlabel metal1 33534 30362 33534 30362 0 _0373_
rlabel metal2 33534 31110 33534 31110 0 _0374_
rlabel metal1 32982 31212 32982 31212 0 _0375_
rlabel metal2 30222 30294 30222 30294 0 _0376_
rlabel metal1 32706 31280 32706 31280 0 _0377_
rlabel metal1 32752 32946 32752 32946 0 _0378_
rlabel metal1 32706 31450 32706 31450 0 _0379_
rlabel metal1 33350 34000 33350 34000 0 _0380_
rlabel metal1 33626 30192 33626 30192 0 _0381_
rlabel metal1 33092 30226 33092 30226 0 _0382_
rlabel metal1 32568 32402 32568 32402 0 _0383_
rlabel metal2 31510 33694 31510 33694 0 _0384_
rlabel metal2 31418 32708 31418 32708 0 _0385_
rlabel metal1 29808 32334 29808 32334 0 _0386_
rlabel metal2 29854 31654 29854 31654 0 _0387_
rlabel metal1 30498 31994 30498 31994 0 _0388_
rlabel metal2 30958 32708 30958 32708 0 _0389_
rlabel metal1 32614 32844 32614 32844 0 _0390_
rlabel metal1 32798 32470 32798 32470 0 _0391_
rlabel metal1 33166 32402 33166 32402 0 _0392_
rlabel metal1 33074 32334 33074 32334 0 _0393_
rlabel metal1 33534 32538 33534 32538 0 _0394_
rlabel metal1 33948 34578 33948 34578 0 _0395_
rlabel metal1 29716 32538 29716 32538 0 _0396_
rlabel via2 33626 34595 33626 34595 0 _0397_
rlabel metal2 33166 36142 33166 36142 0 _0398_
rlabel metal1 33534 34714 33534 34714 0 _0399_
rlabel metal1 34086 35054 34086 35054 0 _0400_
rlabel viali 32982 32879 32982 32879 0 _0401_
rlabel metal1 33718 35054 33718 35054 0 _0402_
rlabel metal1 32706 35734 32706 35734 0 _0403_
rlabel metal1 32752 35802 32752 35802 0 _0404_
rlabel via1 27301 41514 27301 41514 0 _0405_
rlabel metal1 32890 36754 32890 36754 0 _0406_
rlabel metal1 30222 35054 30222 35054 0 _0407_
rlabel metal2 30314 35428 30314 35428 0 _0408_
rlabel metal1 32476 36686 32476 36686 0 _0409_
rlabel metal1 33488 35666 33488 35666 0 _0410_
rlabel metal1 33718 35258 33718 35258 0 _0411_
rlabel metal1 33948 35802 33948 35802 0 _0412_
rlabel metal1 35512 40494 35512 40494 0 _0413_
rlabel metal1 34362 39950 34362 39950 0 _0414_
rlabel metal1 35650 38284 35650 38284 0 _0415_
rlabel metal1 35466 38352 35466 38352 0 _0416_
rlabel metal1 33994 38794 33994 38794 0 _0417_
rlabel metal2 34086 37264 34086 37264 0 _0418_
rlabel metal1 33074 37842 33074 37842 0 _0419_
rlabel metal1 33254 37978 33254 37978 0 _0420_
rlabel metal1 34822 38862 34822 38862 0 _0421_
rlabel metal1 35374 38896 35374 38896 0 _0422_
rlabel metal1 33350 40052 33350 40052 0 _0423_
rlabel metal2 35466 39508 35466 39508 0 _0424_
rlabel metal2 35282 40324 35282 40324 0 _0425_
rlabel metal1 33258 38896 33258 38896 0 _0426_
rlabel metal1 30820 42670 30820 42670 0 _0427_
rlabel metal1 33166 38998 33166 38998 0 _0428_
rlabel metal1 33028 38930 33028 38930 0 _0429_
rlabel metal1 34086 41106 34086 41106 0 _0430_
rlabel metal1 34914 41616 34914 41616 0 _0431_
rlabel metal1 34408 41174 34408 41174 0 _0432_
rlabel metal1 34454 41548 34454 41548 0 _0433_
rlabel metal1 33948 41242 33948 41242 0 _0434_
rlabel metal1 33810 42228 33810 42228 0 _0435_
rlabel metal1 34684 42058 34684 42058 0 _0436_
rlabel metal1 33994 42602 33994 42602 0 _0437_
rlabel metal1 33442 41786 33442 41786 0 _0438_
rlabel metal1 31142 41650 31142 41650 0 _0439_
rlabel metal2 32430 40086 32430 40086 0 _0440_
rlabel metal1 32614 41140 32614 41140 0 _0441_
rlabel metal1 31050 41548 31050 41548 0 _0442_
rlabel metal2 31786 42432 31786 42432 0 _0443_
rlabel metal2 32154 41055 32154 41055 0 _0444_
rlabel metal1 31280 41582 31280 41582 0 _0445_
rlabel metal1 31694 41480 31694 41480 0 _0446_
rlabel metal1 30360 41582 30360 41582 0 _0447_
rlabel metal1 31142 42194 31142 42194 0 _0448_
rlabel via1 29859 41514 29859 41514 0 _0449_
rlabel metal1 29816 41592 29816 41592 0 _0450_
rlabel metal1 31970 41990 31970 41990 0 _0451_
rlabel via1 31878 41123 31878 41123 0 _0452_
rlabel metal1 30958 38930 30958 38930 0 _0453_
rlabel metal1 29946 39542 29946 39542 0 _0454_
rlabel metal1 29716 39066 29716 39066 0 _0455_
rlabel metal1 30222 38998 30222 38998 0 _0456_
rlabel metal1 29854 38352 29854 38352 0 _0457_
rlabel metal2 29762 38522 29762 38522 0 _0458_
rlabel metal1 29854 37196 29854 37196 0 _0459_
rlabel metal2 30038 37434 30038 37434 0 _0460_
rlabel metal1 30682 36822 30682 36822 0 _0461_
rlabel metal2 29302 36822 29302 36822 0 _0462_
rlabel metal1 29210 36788 29210 36788 0 _0463_
rlabel metal1 30958 36346 30958 36346 0 _0464_
rlabel metal1 35466 36822 35466 36822 0 _0465_
rlabel metal1 25300 36754 25300 36754 0 _0466_
rlabel metal1 23920 37842 23920 37842 0 _0467_
rlabel metal2 16146 40358 16146 40358 0 _0468_
rlabel metal1 21988 38930 21988 38930 0 _0469_
rlabel metal1 19550 38896 19550 38896 0 _0470_
rlabel metal1 15870 39984 15870 39984 0 _0471_
rlabel metal1 11454 40494 11454 40494 0 _0472_
rlabel metal1 9752 39610 9752 39610 0 _0473_
rlabel metal2 8326 39882 8326 39882 0 _0474_
rlabel metal1 19113 41582 19113 41582 0 _0475_
rlabel metal1 6026 38930 6026 38930 0 _0476_
rlabel metal1 4462 41072 4462 41072 0 _0477_
rlabel metal1 4370 41242 4370 41242 0 _0478_
rlabel metal1 4370 41616 4370 41616 0 _0479_
rlabel metal1 6440 41786 6440 41786 0 _0480_
rlabel metal1 8280 41718 8280 41718 0 _0481_
rlabel metal1 11408 41582 11408 41582 0 _0482_
rlabel metal1 14306 42738 14306 42738 0 _0483_
rlabel metal2 15594 42500 15594 42500 0 _0484_
rlabel metal1 19918 41684 19918 41684 0 _0485_
rlabel metal1 24380 42330 24380 42330 0 _0486_
rlabel metal1 27186 41616 27186 41616 0 _0487_
rlabel metal2 27002 42330 27002 42330 0 _0488_
rlabel metal1 28106 40052 28106 40052 0 _0489_
rlabel metal1 26818 40052 26818 40052 0 _0490_
rlabel metal1 26818 39950 26818 39950 0 _0491_
rlabel metal1 26496 39814 26496 39814 0 _0492_
rlabel metal1 27771 39066 27771 39066 0 _0493_
rlabel metal1 27784 38726 27784 38726 0 _0494_
rlabel metal1 25668 39066 25668 39066 0 _0495_
rlabel metal1 36064 31790 36064 31790 0 _0496_
rlabel metal1 42826 33422 42826 33422 0 _0497_
rlabel metal1 42596 34170 42596 34170 0 _0498_
rlabel metal1 42596 31450 42596 31450 0 _0499_
rlabel metal1 43516 33490 43516 33490 0 _0500_
rlabel metal1 40526 31994 40526 31994 0 _0501_
rlabel metal1 39514 32980 39514 32980 0 _0502_
rlabel metal1 38456 31790 38456 31790 0 _0503_
rlabel metal1 37444 30226 37444 30226 0 _0504_
rlabel metal1 35972 38318 35972 38318 0 _0505_
rlabel metal1 41860 36618 41860 36618 0 _0506_
rlabel metal1 37398 36652 37398 36652 0 _0507_
rlabel metal1 37490 36822 37490 36822 0 _0508_
rlabel metal1 37858 36822 37858 36822 0 _0509_
rlabel metal1 41446 36720 41446 36720 0 _0510_
rlabel metal1 21206 41072 21206 41072 0 _0511_
rlabel metal1 18400 41650 18400 41650 0 _0512_
rlabel metal1 15456 19278 15456 19278 0 _0513_
rlabel metal1 17618 23290 17618 23290 0 _0514_
rlabel metal1 18446 21998 18446 21998 0 _0515_
rlabel metal1 18216 20298 18216 20298 0 _0516_
rlabel metal1 16974 21318 16974 21318 0 _0517_
rlabel metal1 17572 19482 17572 19482 0 _0518_
rlabel metal2 15226 19142 15226 19142 0 _0519_
rlabel metal1 12604 19346 12604 19346 0 _0520_
rlabel metal1 11224 19346 11224 19346 0 _0521_
rlabel metal1 15824 24242 15824 24242 0 _0522_
rlabel metal1 12972 23086 12972 23086 0 _0523_
rlabel metal1 14996 24174 14996 24174 0 _0524_
rlabel metal1 12190 23834 12190 23834 0 _0525_
rlabel metal1 11822 26554 11822 26554 0 _0526_
rlabel metal1 13018 25262 13018 25262 0 _0527_
rlabel metal2 21390 28934 21390 28934 0 _0528_
rlabel metal1 22724 28730 22724 28730 0 _0529_
rlabel metal1 24656 31790 24656 31790 0 _0530_
rlabel metal2 25990 31892 25990 31892 0 _0531_
rlabel metal1 22540 31790 22540 31790 0 _0532_
rlabel metal1 22310 12750 22310 12750 0 _0533_
rlabel metal1 18998 17102 18998 17102 0 _0534_
rlabel metal1 14030 6086 14030 6086 0 _0535_
rlabel metal1 12098 8942 12098 8942 0 _0536_
rlabel metal1 12834 4046 12834 4046 0 _0537_
rlabel metal1 14950 7310 14950 7310 0 _0538_
rlabel metal1 13248 7174 13248 7174 0 _0539_
rlabel metal1 14628 10574 14628 10574 0 _0540_
rlabel metal1 14398 11832 14398 11832 0 _0541_
rlabel metal1 13570 10166 13570 10166 0 _0542_
rlabel metal1 14858 2924 14858 2924 0 _0543_
rlabel metal1 14076 9554 14076 9554 0 _0544_
rlabel metal1 15410 15538 15410 15538 0 _0545_
rlabel metal2 15502 7718 15502 7718 0 _0546_
rlabel metal1 11730 14960 11730 14960 0 _0547_
rlabel metal1 13524 7378 13524 7378 0 _0548_
rlabel metal2 13754 7786 13754 7786 0 _0549_
rlabel metal2 18170 15504 18170 15504 0 _0550_
rlabel metal1 16560 8942 16560 8942 0 _0551_
rlabel metal1 12788 9622 12788 9622 0 _0552_
rlabel metal1 17664 16762 17664 16762 0 _0553_
rlabel metal1 14582 13872 14582 13872 0 _0554_
rlabel metal1 20746 13872 20746 13872 0 _0555_
rlabel metal1 17250 3910 17250 3910 0 _0556_
rlabel metal1 17480 15062 17480 15062 0 _0557_
rlabel metal1 13432 9146 13432 9146 0 _0558_
rlabel metal1 18078 11016 18078 11016 0 _0559_
rlabel metal1 17158 16762 17158 16762 0 _0560_
rlabel metal1 12374 12716 12374 12716 0 _0561_
rlabel metal1 15134 4454 15134 4454 0 _0562_
rlabel metal1 11500 7446 11500 7446 0 _0563_
rlabel metal2 15778 7106 15778 7106 0 _0564_
rlabel metal1 16514 9894 16514 9894 0 _0565_
rlabel metal1 16836 9350 16836 9350 0 _0566_
rlabel metal2 15502 10914 15502 10914 0 _0567_
rlabel metal1 12190 6970 12190 6970 0 _0568_
rlabel metal2 19550 7888 19550 7888 0 _0569_
rlabel metal1 17526 16082 17526 16082 0 _0570_
rlabel metal1 17756 15946 17756 15946 0 _0571_
rlabel metal1 16008 9010 16008 9010 0 _0572_
rlabel via3 17227 15300 17227 15300 0 _0573_
rlabel metal1 17526 15878 17526 15878 0 _0574_
rlabel metal1 19458 9996 19458 9996 0 _0575_
rlabel metal2 17250 10880 17250 10880 0 _0576_
rlabel metal1 19642 7922 19642 7922 0 _0577_
rlabel metal2 11454 14144 11454 14144 0 _0578_
rlabel metal1 18906 16966 18906 16966 0 _0579_
rlabel metal1 32154 5780 32154 5780 0 _0580_
rlabel metal1 32200 15402 32200 15402 0 _0581_
rlabel metal1 31326 15504 31326 15504 0 _0582_
rlabel metal1 29854 14960 29854 14960 0 _0583_
rlabel metal1 30268 14382 30268 14382 0 _0584_
rlabel via1 30037 8466 30037 8466 0 _0585_
rlabel metal1 32108 13294 32108 13294 0 _0586_
rlabel metal1 30636 13158 30636 13158 0 _0587_
rlabel metal1 30682 15028 30682 15028 0 _0588_
rlabel metal1 31326 15028 31326 15028 0 _0589_
rlabel metal1 30958 14994 30958 14994 0 _0590_
rlabel metal1 30176 9418 30176 9418 0 _0591_
rlabel metal1 31970 9588 31970 9588 0 _0592_
rlabel metal1 32062 8976 32062 8976 0 _0593_
rlabel metal2 31602 8636 31602 8636 0 _0594_
rlabel metal1 32154 12852 32154 12852 0 _0595_
rlabel metal1 31280 12682 31280 12682 0 _0596_
rlabel metal2 29026 11968 29026 11968 0 _0597_
rlabel metal1 28842 8466 28842 8466 0 _0598_
rlabel metal1 30774 8364 30774 8364 0 _0599_
rlabel metal1 31234 9554 31234 9554 0 _0600_
rlabel metal1 29624 8942 29624 8942 0 _0601_
rlabel metal1 27370 9452 27370 9452 0 _0602_
rlabel metal1 29440 12206 29440 12206 0 _0603_
rlabel metal1 28382 11628 28382 11628 0 _0604_
rlabel metal1 30866 11730 30866 11730 0 _0605_
rlabel metal1 29900 11866 29900 11866 0 _0606_
rlabel metal1 28842 8942 28842 8942 0 _0607_
rlabel metal1 31234 10030 31234 10030 0 _0608_
rlabel metal2 28382 10574 28382 10574 0 _0609_
rlabel metal1 27462 9452 27462 9452 0 _0610_
rlabel metal1 27554 9554 27554 9554 0 _0611_
rlabel metal2 25990 10574 25990 10574 0 _0612_
rlabel metal1 30820 12750 30820 12750 0 _0613_
rlabel metal1 28934 9112 28934 9112 0 _0614_
rlabel metal1 27094 7922 27094 7922 0 _0615_
rlabel metal1 29302 10642 29302 10642 0 _0616_
rlabel metal1 28428 11118 28428 11118 0 _0617_
rlabel metal1 27830 11050 27830 11050 0 _0618_
rlabel metal1 30222 10234 30222 10234 0 _0619_
rlabel metal1 28566 10540 28566 10540 0 _0620_
rlabel metal1 27830 8602 27830 8602 0 _0621_
rlabel metal1 26220 14994 26220 14994 0 _0622_
rlabel metal2 25806 7616 25806 7616 0 _0623_
rlabel metal1 25852 9146 25852 9146 0 _0624_
rlabel metal1 23184 15878 23184 15878 0 _0625_
rlabel metal1 27002 14416 27002 14416 0 _0626_
rlabel metal1 30866 11118 30866 11118 0 _0627_
rlabel via2 31418 11101 31418 11101 0 _0628_
rlabel metal2 30774 10574 30774 10574 0 _0629_
rlabel metal2 32246 10778 32246 10778 0 _0630_
rlabel metal1 32338 8908 32338 8908 0 _0631_
rlabel metal1 31004 8466 31004 8466 0 _0632_
rlabel metal1 26082 10540 26082 10540 0 _0633_
rlabel metal1 25852 10778 25852 10778 0 _0634_
rlabel metal2 29210 10404 29210 10404 0 _0635_
rlabel metal1 31970 11084 31970 11084 0 _0636_
rlabel metal1 29578 10438 29578 10438 0 _0637_
rlabel metal1 27186 10710 27186 10710 0 _0638_
rlabel metal2 28106 9860 28106 9860 0 _0639_
rlabel metal1 26174 10710 26174 10710 0 _0640_
rlabel metal2 24886 12342 24886 12342 0 _0641_
rlabel metal1 22172 8466 22172 8466 0 _0642_
rlabel metal1 20562 15368 20562 15368 0 _0643_
rlabel metal2 19274 19346 19274 19346 0 _0644_
rlabel metal1 19918 21454 19918 21454 0 _0645_
rlabel metal1 19044 21522 19044 21522 0 _0646_
rlabel metal2 14582 10812 14582 10812 0 _0647_
rlabel metal1 13386 14042 13386 14042 0 _0648_
rlabel metal1 15594 11186 15594 11186 0 _0649_
rlabel metal1 19182 9520 19182 9520 0 _0650_
rlabel metal1 16698 5746 16698 5746 0 _0651_
rlabel via1 12558 12631 12558 12631 0 _0652_
rlabel metal1 17940 6766 17940 6766 0 _0653_
rlabel metal1 17480 10642 17480 10642 0 _0654_
rlabel metal1 16468 10778 16468 10778 0 _0655_
rlabel metal1 19044 6154 19044 6154 0 _0656_
rlabel metal1 20010 7854 20010 7854 0 _0657_
rlabel metal2 15870 16830 15870 16830 0 _0658_
rlabel metal2 13386 12619 13386 12619 0 _0659_
rlabel metal1 15640 12206 15640 12206 0 _0660_
rlabel metal1 16848 11186 16848 11186 0 _0661_
rlabel metal1 14076 9010 14076 9010 0 _0662_
rlabel metal1 16146 9690 16146 9690 0 _0663_
rlabel metal1 16514 10064 16514 10064 0 _0664_
rlabel metal2 16882 10676 16882 10676 0 _0665_
rlabel metal1 19366 11288 19366 11288 0 _0666_
rlabel metal1 30122 7718 30122 7718 0 _0667_
rlabel metal1 28382 7786 28382 7786 0 _0668_
rlabel metal1 26174 8466 26174 8466 0 _0669_
rlabel metal1 25714 8942 25714 8942 0 _0670_
rlabel metal1 23092 8942 23092 8942 0 _0671_
rlabel metal1 22678 9622 22678 9622 0 _0672_
rlabel metal1 24288 10234 24288 10234 0 _0673_
rlabel metal2 22126 7616 22126 7616 0 _0674_
rlabel metal2 22678 10948 22678 10948 0 _0675_
rlabel metal2 23276 12614 23276 12614 0 _0676_
rlabel metal1 21666 20570 21666 20570 0 _0677_
rlabel metal2 27922 8126 27922 8126 0 _0678_
rlabel metal1 27140 14994 27140 14994 0 _0679_
rlabel metal1 25438 15538 25438 15538 0 _0680_
rlabel metal1 25208 11594 25208 11594 0 _0681_
rlabel metal1 19826 17272 19826 17272 0 _0682_
rlabel metal2 15318 15606 15318 15606 0 _0683_
rlabel metal1 16008 16626 16008 16626 0 _0684_
rlabel metal1 19780 7514 19780 7514 0 _0685_
rlabel metal2 20378 7837 20378 7837 0 _0686_
rlabel metal1 15410 16218 15410 16218 0 _0687_
rlabel metal1 19366 17238 19366 17238 0 _0688_
rlabel metal1 15134 11832 15134 11832 0 _0689_
rlabel metal1 14812 12954 14812 12954 0 _0690_
rlabel metal1 15548 12818 15548 12818 0 _0691_
rlabel metal1 14766 12750 14766 12750 0 _0692_
rlabel metal1 17250 13362 17250 13362 0 _0693_
rlabel metal1 19596 16218 19596 16218 0 _0694_
rlabel metal2 20010 18496 20010 18496 0 _0695_
rlabel metal1 18906 19890 18906 19890 0 _0696_
rlabel metal1 29118 10030 29118 10030 0 _0697_
rlabel metal1 28336 10234 28336 10234 0 _0698_
rlabel metal1 25668 8602 25668 8602 0 _0699_
rlabel metal1 24518 8874 24518 8874 0 _0700_
rlabel metal1 25162 9044 25162 9044 0 _0701_
rlabel metal1 24288 8806 24288 8806 0 _0702_
rlabel metal1 22034 8500 22034 8500 0 _0703_
rlabel metal1 14168 6426 14168 6426 0 _0704_
rlabel metal1 19458 6732 19458 6732 0 _0705_
rlabel metal2 16238 6222 16238 6222 0 _0706_
rlabel metal2 15226 6596 15226 6596 0 _0707_
rlabel metal1 17894 5542 17894 5542 0 _0708_
rlabel metal1 19136 6290 19136 6290 0 _0709_
rlabel metal1 19688 6426 19688 6426 0 _0710_
rlabel metal1 20102 6834 20102 6834 0 _0711_
rlabel metal1 21298 6834 21298 6834 0 _0712_
rlabel metal2 21850 8228 21850 8228 0 _0713_
rlabel metal1 21666 19890 21666 19890 0 _0714_
rlabel metal1 20838 20570 20838 20570 0 _0715_
rlabel metal1 20884 15130 20884 15130 0 _0716_
rlabel metal1 19596 14926 19596 14926 0 _0717_
rlabel metal2 14766 14127 14766 14127 0 _0718_
rlabel metal1 20516 14994 20516 14994 0 _0719_
rlabel metal2 20746 15164 20746 15164 0 _0720_
rlabel metal1 21574 15436 21574 15436 0 _0721_
rlabel metal1 13064 13294 13064 13294 0 _0722_
rlabel metal1 14398 14042 14398 14042 0 _0723_
rlabel metal1 14030 14858 14030 14858 0 _0724_
rlabel metal1 13133 13974 13133 13974 0 _0725_
rlabel metal1 14490 14586 14490 14586 0 _0726_
rlabel metal2 20838 13056 20838 13056 0 _0727_
rlabel metal2 14582 15351 14582 15351 0 _0728_
rlabel metal1 28658 11696 28658 11696 0 _0729_
rlabel metal1 28612 11322 28612 11322 0 _0730_
rlabel metal1 27968 11798 27968 11798 0 _0731_
rlabel metal1 27140 14382 27140 14382 0 _0732_
rlabel metal1 23414 15028 23414 15028 0 _0733_
rlabel metal2 21942 15266 21942 15266 0 _0734_
rlabel metal2 21758 15708 21758 15708 0 _0735_
rlabel metal1 21252 15674 21252 15674 0 _0736_
rlabel metal1 20608 18258 20608 18258 0 _0737_
rlabel metal1 18124 5882 18124 5882 0 _0738_
rlabel metal1 16238 6426 16238 6426 0 _0739_
rlabel metal2 17986 7106 17986 7106 0 _0740_
rlabel metal1 16606 6834 16606 6834 0 _0741_
rlabel metal1 17158 6970 17158 6970 0 _0742_
rlabel metal1 17296 8806 17296 8806 0 _0743_
rlabel metal2 17986 8228 17986 8228 0 _0744_
rlabel metal1 17802 7820 17802 7820 0 _0745_
rlabel metal1 18446 7412 18446 7412 0 _0746_
rlabel metal1 17710 7344 17710 7344 0 _0747_
rlabel metal1 17250 7378 17250 7378 0 _0748_
rlabel metal2 17434 7888 17434 7888 0 _0749_
rlabel metal1 22954 8874 22954 8874 0 _0750_
rlabel metal2 25162 11526 25162 11526 0 _0751_
rlabel metal2 22770 10812 22770 10812 0 _0752_
rlabel metal1 22954 9044 22954 9044 0 _0753_
rlabel via3 22701 16660 22701 16660 0 _0754_
rlabel metal1 22172 17850 22172 17850 0 _0755_
rlabel metal1 30866 11866 30866 11866 0 _0756_
rlabel metal1 29900 12410 29900 12410 0 _0757_
rlabel metal1 28934 13294 28934 13294 0 _0758_
rlabel metal2 26542 13702 26542 13702 0 _0759_
rlabel metal1 27048 14586 27048 14586 0 _0760_
rlabel metal1 25806 15402 25806 15402 0 _0761_
rlabel metal1 25208 15674 25208 15674 0 _0762_
rlabel metal1 19642 18156 19642 18156 0 _0763_
rlabel metal1 13570 9996 13570 9996 0 _0764_
rlabel metal1 14858 10200 14858 10200 0 _0765_
rlabel metal1 18446 11696 18446 11696 0 _0766_
rlabel metal1 19366 11084 19366 11084 0 _0767_
rlabel metal1 19228 4590 19228 4590 0 _0768_
rlabel metal1 19136 11186 19136 11186 0 _0769_
rlabel metal1 18906 18122 18906 18122 0 _0770_
rlabel metal1 17756 14042 17756 14042 0 _0771_
rlabel metal1 17435 14926 17435 14926 0 _0772_
rlabel metal1 18262 15130 18262 15130 0 _0773_
rlabel metal2 18814 17476 18814 17476 0 _0774_
rlabel metal1 19550 18224 19550 18224 0 _0775_
rlabel metal1 12650 11866 12650 11866 0 _0776_
rlabel metal1 12581 10098 12581 10098 0 _0777_
rlabel metal1 11500 9350 11500 9350 0 _0778_
rlabel metal1 12742 9486 12742 9486 0 _0779_
rlabel metal1 11454 6766 11454 6766 0 _0780_
rlabel metal2 11914 8432 11914 8432 0 _0781_
rlabel metal1 12098 9690 12098 9690 0 _0782_
rlabel via2 11086 10251 11086 10251 0 _0783_
rlabel metal1 29164 12614 29164 12614 0 _0784_
rlabel metal1 28336 12750 28336 12750 0 _0785_
rlabel metal1 26726 12886 26726 12886 0 _0786_
rlabel metal1 24196 11866 24196 11866 0 _0787_
rlabel metal1 23782 9690 23782 9690 0 _0788_
rlabel metal1 22126 10540 22126 10540 0 _0789_
rlabel via3 22517 18020 22517 18020 0 _0790_
rlabel metal1 21758 18938 21758 18938 0 _0791_
rlabel metal1 12328 14994 12328 14994 0 _0792_
rlabel metal1 12926 15130 12926 15130 0 _0793_
rlabel viali 13205 14858 13205 14858 0 _0794_
rlabel metal1 13340 15538 13340 15538 0 _0795_
rlabel metal1 12006 14382 12006 14382 0 _0796_
rlabel metal1 12098 14994 12098 14994 0 _0797_
rlabel metal2 12190 15300 12190 15300 0 _0798_
rlabel metal1 11500 12818 11500 12818 0 _0799_
rlabel metal1 11730 13260 11730 13260 0 _0800_
rlabel metal1 12144 13498 12144 13498 0 _0801_
rlabel via2 11454 15419 11454 15419 0 _0802_
rlabel metal1 22540 15402 22540 15402 0 _0803_
rlabel metal1 27416 13362 27416 13362 0 _0804_
rlabel metal1 26680 14246 26680 14246 0 _0805_
rlabel metal1 24610 14790 24610 14790 0 _0806_
rlabel metal1 22632 15130 22632 15130 0 _0807_
rlabel metal1 22816 23086 22816 23086 0 _0808_
rlabel metal1 22586 22610 22586 22610 0 _0809_
rlabel metal1 18492 14246 18492 14246 0 _0810_
rlabel metal2 16514 15810 16514 15810 0 _0811_
rlabel metal1 18630 14348 18630 14348 0 _0812_
rlabel metal1 18952 13702 18952 13702 0 _0813_
rlabel viali 18077 12818 18077 12818 0 _0814_
rlabel metal1 18170 12954 18170 12954 0 _0815_
rlabel metal1 19780 14042 19780 14042 0 _0816_
rlabel metal2 15962 13532 15962 13532 0 _0817_
rlabel metal1 15410 14586 15410 14586 0 _0818_
rlabel metal1 20102 13940 20102 13940 0 _0819_
rlabel metal1 17434 14450 17434 14450 0 _0820_
rlabel metal1 19090 14484 19090 14484 0 _0821_
rlabel metal1 20470 14450 20470 14450 0 _0822_
rlabel metal2 23414 7752 23414 7752 0 _0823_
rlabel metal1 25990 13260 25990 13260 0 _0824_
rlabel metal1 24288 12954 24288 12954 0 _0825_
rlabel metal1 21298 14314 21298 14314 0 _0826_
rlabel metal2 20884 14586 20884 14586 0 _0827_
rlabel metal1 19688 23086 19688 23086 0 _0828_
rlabel metal1 25438 13906 25438 13906 0 _0829_
rlabel metal1 25024 15334 25024 15334 0 _0830_
rlabel metal1 24380 15674 24380 15674 0 _0831_
rlabel metal1 12052 8058 12052 8058 0 _0832_
rlabel metal1 11638 11866 11638 11866 0 _0833_
rlabel metal1 12236 12818 12236 12818 0 _0834_
rlabel metal1 11730 12682 11730 12682 0 _0835_
rlabel metal1 11592 12954 11592 12954 0 _0836_
rlabel metal1 12696 13498 12696 13498 0 _0837_
rlabel metal1 11960 14042 11960 14042 0 _0838_
rlabel metal2 12006 14739 12006 14739 0 _0839_
rlabel metal1 21068 15674 21068 15674 0 _0840_
rlabel metal1 22011 16150 22011 16150 0 _0841_
rlabel metal1 21298 22746 21298 22746 0 _0842_
rlabel metal2 14306 16796 14306 16796 0 _0843_
rlabel metal1 14950 11866 14950 11866 0 _0844_
rlabel metal1 14490 16218 14490 16218 0 _0845_
rlabel metal1 14490 15436 14490 15436 0 _0846_
rlabel metal1 14858 15674 14858 15674 0 _0847_
rlabel metal1 13888 11866 13888 11866 0 _0848_
rlabel metal1 16376 16762 16376 16762 0 _0849_
rlabel metal1 26312 13362 26312 13362 0 _0850_
rlabel metal1 25714 16082 25714 16082 0 _0851_
rlabel metal2 23414 16354 23414 16354 0 _0852_
rlabel metal1 20470 17068 20470 17068 0 _0853_
rlabel metal1 20424 17306 20424 17306 0 _0854_
rlabel metal2 20562 25568 20562 25568 0 _0855_
rlabel metal1 19642 24922 19642 24922 0 _0856_
rlabel metal1 17158 12342 17158 12342 0 _0857_
rlabel metal1 17687 12410 17687 12410 0 _0858_
rlabel metal1 20608 10098 20608 10098 0 _0859_
rlabel metal1 20286 11764 20286 11764 0 _0860_
rlabel metal1 20332 12682 20332 12682 0 _0861_
rlabel metal2 20654 11713 20654 11713 0 _0862_
rlabel metal1 19366 11696 19366 11696 0 _0863_
rlabel metal1 20010 11866 20010 11866 0 _0864_
rlabel metal1 23828 10778 23828 10778 0 _0865_
rlabel metal1 21229 12750 21229 12750 0 _0866_
rlabel metal1 20056 12954 20056 12954 0 _0867_
rlabel metal1 19504 25874 19504 25874 0 _0868_
rlabel metal1 22448 12954 22448 12954 0 _0869_
rlabel metal1 20884 12410 20884 12410 0 _0870_
rlabel metal1 19550 12954 19550 12954 0 _0871_
rlabel metal1 19458 9452 19458 9452 0 _0872_
rlabel metal1 19504 9622 19504 9622 0 _0873_
rlabel metal1 20654 12852 20654 12852 0 _0874_
rlabel metal1 21528 12954 21528 12954 0 _0875_
rlabel metal2 22310 14773 22310 14773 0 _0876_
rlabel metal1 21666 25874 21666 25874 0 _0877_
rlabel metal2 20102 8738 20102 8738 0 _0878_
rlabel metal1 19964 8942 19964 8942 0 _0879_
rlabel metal1 20010 8840 20010 8840 0 _0880_
rlabel metal1 20194 9146 20194 9146 0 _0881_
rlabel metal1 20240 7786 20240 7786 0 _0882_
rlabel metal2 23874 15470 23874 15470 0 _0883_
rlabel metal1 24150 15674 24150 15674 0 _0884_
rlabel metal1 24058 28050 24058 28050 0 _0885_
rlabel metal1 20010 14926 20010 14926 0 _0886_
rlabel metal1 19826 9486 19826 9486 0 _0887_
rlabel metal1 19688 9350 19688 9350 0 _0888_
rlabel metal1 21114 14926 21114 14926 0 _0889_
rlabel metal2 25162 17544 25162 17544 0 _0890_
rlabel metal1 24150 27030 24150 27030 0 _0891_
rlabel metal1 21206 6970 21206 6970 0 _0892_
rlabel metal1 20746 7310 20746 7310 0 _0893_
rlabel metal1 21758 7378 21758 7378 0 _0894_
rlabel metal1 24702 13838 24702 13838 0 _0895_
rlabel metal1 24748 14042 24748 14042 0 _0896_
rlabel metal1 25484 28050 25484 28050 0 _0897_
rlabel metal2 22954 9860 22954 9860 0 _0898_
rlabel metal1 22034 12206 22034 12206 0 _0899_
rlabel metal1 22678 12410 22678 12410 0 _0900_
rlabel metal1 22310 27098 22310 27098 0 _0901_
rlabel metal2 16790 25398 16790 25398 0 _0902_
rlabel metal1 17940 24786 17940 24786 0 _0903_
rlabel metal1 17526 25874 17526 25874 0 _0904_
rlabel via1 15226 20366 15226 20366 0 _0905_
rlabel metal1 15272 22610 15272 22610 0 _0906_
rlabel metal1 15640 20434 15640 20434 0 _0907_
rlabel metal2 14674 21828 14674 21828 0 _0908_
rlabel metal1 12167 20434 12167 20434 0 _0909_
rlabel metal1 10396 20434 10396 20434 0 _0910_
rlabel metal1 10534 23834 10534 23834 0 _0911_
rlabel metal1 13984 25262 13984 25262 0 _0912_
rlabel metal1 9200 23086 9200 23086 0 _0913_
rlabel metal1 10166 25262 10166 25262 0 _0914_
rlabel metal1 8694 25262 8694 25262 0 _0915_
rlabel metal2 18446 35904 18446 35904 0 _0916_
rlabel metal1 19550 29818 19550 29818 0 _0917_
rlabel metal1 20884 31994 20884 31994 0 _0918_
rlabel metal1 23184 31994 23184 31994 0 _0919_
rlabel metal1 24656 33082 24656 33082 0 _0920_
rlabel metal1 22264 31790 22264 31790 0 _0921_
rlabel metal1 24058 35666 24058 35666 0 _0922_
rlabel metal2 22402 35428 22402 35428 0 _0923_
rlabel metal1 19780 35802 19780 35802 0 _0924_
rlabel metal1 17894 38386 17894 38386 0 _0925_
rlabel metal1 17848 37230 17848 37230 0 _0926_
rlabel metal1 16376 37842 16376 37842 0 _0927_
rlabel metal1 14398 38896 14398 38896 0 _0928_
rlabel metal1 7682 38318 7682 38318 0 _0929_
rlabel metal2 7590 34102 7590 34102 0 _0930_
rlabel metal1 2530 34578 2530 34578 0 _0931_
rlabel metal1 2024 32878 2024 32878 0 _0932_
rlabel metal1 5658 33626 5658 33626 0 _0933_
rlabel metal2 2622 39236 2622 39236 0 _0934_
rlabel metal1 5336 37230 5336 37230 0 _0935_
rlabel metal1 19826 43758 19826 43758 0 _0936_
rlabel metal1 9844 44506 9844 44506 0 _0937_
rlabel metal1 11362 44438 11362 44438 0 _0938_
rlabel metal1 13984 43962 13984 43962 0 _0939_
rlabel metal2 16698 43962 16698 43962 0 _0940_
rlabel metal1 19090 43962 19090 43962 0 _0941_
rlabel metal1 23230 36210 23230 36210 0 _0942_
rlabel metal1 20792 36754 20792 36754 0 _0943_
rlabel metal1 19412 36890 19412 36890 0 _0944_
rlabel metal1 18768 37434 18768 37434 0 _0945_
rlabel metal1 15364 39066 15364 39066 0 _0946_
rlabel metal2 12190 39950 12190 39950 0 _0947_
rlabel metal1 11776 38930 11776 38930 0 _0948_
rlabel metal1 8234 37230 8234 37230 0 _0949_
rlabel metal1 7452 32402 7452 32402 0 _0950_
rlabel metal1 3772 35054 3772 35054 0 _0951_
rlabel metal1 3588 33082 3588 33082 0 _0952_
rlabel metal1 3864 33490 3864 33490 0 _0953_
rlabel metal1 3358 37434 3358 37434 0 _0954_
rlabel metal2 7130 37434 7130 37434 0 _0955_
rlabel metal1 8740 41582 8740 41582 0 _0956_
rlabel metal1 11132 41106 11132 41106 0 _0957_
rlabel metal1 13248 41786 13248 41786 0 _0958_
rlabel metal1 15226 41106 15226 41106 0 _0959_
rlabel metal1 18952 41786 18952 41786 0 _0960_
rlabel metal1 24196 34714 24196 34714 0 _0961_
rlabel metal1 21574 33490 21574 33490 0 _0962_
rlabel metal1 19688 34714 19688 34714 0 _0963_
rlabel metal1 17986 35258 17986 35258 0 _0964_
rlabel metal1 16514 35666 16514 35666 0 _0965_
rlabel metal2 12558 43996 12558 43996 0 _0966_
rlabel metal1 13616 40154 13616 40154 0 _0967_
rlabel metal1 9430 37978 9430 37978 0 _0968_
rlabel metal1 8694 33626 8694 33626 0 _0969_
rlabel metal1 3680 30702 3680 30702 0 _0970_
rlabel metal1 2300 31314 2300 31314 0 _0971_
rlabel metal1 6256 32266 6256 32266 0 _0972_
rlabel metal1 2300 37230 2300 37230 0 _0973_
rlabel metal1 5428 35802 5428 35802 0 _0974_
rlabel metal1 9016 45458 9016 45458 0 _0975_
rlabel metal1 11684 44506 11684 44506 0 _0976_
rlabel metal1 14996 44846 14996 44846 0 _0977_
rlabel metal1 16698 45390 16698 45390 0 _0978_
rlabel metal1 18400 43962 18400 43962 0 _0979_
rlabel metal1 18354 3502 18354 3502 0 _0980_
rlabel metal1 18676 3570 18676 3570 0 _0981_
rlabel metal1 17756 3162 17756 3162 0 _0982_
rlabel metal1 20378 4726 20378 4726 0 _0983_
rlabel metal1 16652 3026 16652 3026 0 _0984_
rlabel metal1 14674 3162 14674 3162 0 _0985_
rlabel metal1 14076 3162 14076 3162 0 _0986_
rlabel metal1 13110 3706 13110 3706 0 _0987_
rlabel metal2 12650 4726 12650 4726 0 _0988_
rlabel metal1 13064 2958 13064 2958 0 _0989_
rlabel metal2 13202 4930 13202 4930 0 _0990_
rlabel metal1 19182 4658 19182 4658 0 _0991_
rlabel metal1 20608 4046 20608 4046 0 _0992_
rlabel metal1 20976 4590 20976 4590 0 _0993_
rlabel metal2 25898 44948 25898 44948 0 _0994_
rlabel metal1 24012 44846 24012 44846 0 _0995_
rlabel metal1 22954 43622 22954 43622 0 _0996_
rlabel metal1 22678 41990 22678 41990 0 _0997_
rlabel metal1 28106 38896 28106 38896 0 _0998_
rlabel metal2 27186 40460 27186 40460 0 _0999_
rlabel metal2 28290 39508 28290 39508 0 _1000_
rlabel metal2 30314 40273 30314 40273 0 _1001_
rlabel metal1 22862 40086 22862 40086 0 _1002_
rlabel metal2 18998 41718 18998 41718 0 _1003_
rlabel metal2 34362 36499 34362 36499 0 _1004_
rlabel metal1 9752 18666 9752 18666 0 _1005_
rlabel metal1 35696 14994 35696 14994 0 _1006_
rlabel metal1 22080 3060 22080 3060 0 _1007_
rlabel metal1 30636 3162 30636 3162 0 _1008_
rlabel metal2 26082 3638 26082 3638 0 _1009_
rlabel metal1 15870 17646 15870 17646 0 _1010_
rlabel metal1 36064 16082 36064 16082 0 _1011_
rlabel metal1 10534 18258 10534 18258 0 _1012_
rlabel viali 33166 16556 33166 16556 0 _1013_
rlabel metal1 26910 3162 26910 3162 0 _1014_
rlabel metal1 9568 18258 9568 18258 0 _1015_
rlabel metal1 25300 43758 25300 43758 0 _1016_
rlabel metal1 7176 13498 7176 13498 0 _1017_
rlabel metal1 7314 17170 7314 17170 0 _1018_
rlabel metal1 7774 12784 7774 12784 0 _1019_
rlabel metal1 43654 12818 43654 12818 0 _1020_
rlabel metal1 8142 16048 8142 16048 0 _1021_
rlabel metal1 43976 32402 43976 32402 0 _1022_
rlabel metal1 44068 14994 44068 14994 0 _1023_
rlabel metal1 34730 4148 34730 4148 0 _1024_
rlabel metal1 35190 4046 35190 4046 0 _1025_
rlabel metal1 35190 4250 35190 4250 0 _1026_
rlabel metal1 33626 3978 33626 3978 0 _1027_
rlabel metal1 36202 3978 36202 3978 0 _1028_
rlabel metal1 36938 4080 36938 4080 0 _1029_
rlabel metal2 38042 5236 38042 5236 0 _1030_
rlabel metal2 33994 3774 33994 3774 0 _1031_
rlabel metal2 39606 6290 39606 6290 0 _1032_
rlabel metal1 41584 7378 41584 7378 0 _1033_
rlabel metal1 41308 5338 41308 5338 0 _1034_
rlabel metal1 39698 7310 39698 7310 0 _1035_
rlabel metal1 39330 7412 39330 7412 0 _1036_
rlabel metal2 39146 8364 39146 8364 0 _1037_
rlabel metal1 39192 6970 39192 6970 0 _1038_
rlabel metal1 36202 5202 36202 5202 0 _1039_
rlabel metal1 38686 3536 38686 3536 0 _1040_
rlabel metal1 38502 3468 38502 3468 0 _1041_
rlabel metal1 40526 4522 40526 4522 0 _1042_
rlabel metal1 39606 4692 39606 4692 0 _1043_
rlabel metal1 40020 3706 40020 3706 0 _1044_
rlabel metal1 40480 4250 40480 4250 0 _1045_
rlabel metal1 40802 4658 40802 4658 0 _1046_
rlabel metal1 41078 4080 41078 4080 0 _1047_
rlabel metal1 41308 4114 41308 4114 0 _1048_
rlabel metal1 42458 5338 42458 5338 0 _1049_
rlabel metal1 42244 4522 42244 4522 0 _1050_
rlabel metal1 43010 4624 43010 4624 0 _1051_
rlabel metal1 41998 8976 41998 8976 0 _1052_
rlabel metal1 42964 6426 42964 6426 0 _1053_
rlabel metal2 42918 7888 42918 7888 0 _1054_
rlabel metal1 42182 9350 42182 9350 0 _1055_
rlabel metal2 41906 9384 41906 9384 0 _1056_
rlabel metal1 41584 9554 41584 9554 0 _1057_
rlabel metal1 40388 8466 40388 8466 0 _1058_
rlabel metal1 43102 7242 43102 7242 0 _1059_
rlabel metal2 37766 6732 37766 6732 0 _1060_
rlabel metal1 39698 7956 39698 7956 0 _1061_
rlabel via1 37946 6426 37946 6426 0 _1062_
rlabel metal1 36938 6358 36938 6358 0 _1063_
rlabel metal1 36892 7514 36892 7514 0 _1064_
rlabel metal1 36846 7888 36846 7888 0 _1065_
rlabel metal2 37398 9894 37398 9894 0 _1066_
rlabel metal1 37490 9418 37490 9418 0 _1067_
rlabel metal1 39698 9146 39698 9146 0 _1068_
rlabel metal1 39179 8806 39179 8806 0 _1069_
rlabel metal1 39422 9078 39422 9078 0 _1070_
rlabel metal1 34546 10030 34546 10030 0 _1071_
rlabel metal1 41078 23732 41078 23732 0 _1072_
rlabel metal1 43102 25330 43102 25330 0 _1073_
rlabel via1 40058 24038 40058 24038 0 _1074_
rlabel metal1 41906 23698 41906 23698 0 _1075_
rlabel metal1 39422 24140 39422 24140 0 _1076_
rlabel metal1 39882 24174 39882 24174 0 _1077_
rlabel metal1 38548 24718 38548 24718 0 _1078_
rlabel metal1 38548 24786 38548 24786 0 _1079_
rlabel metal1 38180 24786 38180 24786 0 _1080_
rlabel metal1 23414 41480 23414 41480 0 _1081_
rlabel metal1 23732 41106 23732 41106 0 _1082_
rlabel metal1 18354 42602 18354 42602 0 _1083_
rlabel metal1 25530 41446 25530 41446 0 _1084_
rlabel via1 26722 44506 26722 44506 0 _1085_
rlabel metal1 23920 44506 23920 44506 0 _1086_
rlabel metal1 23506 43826 23506 43826 0 _1087_
rlabel metal1 21942 42126 21942 42126 0 _1088_
rlabel metal1 17250 45458 17250 45458 0 _1089_
rlabel metal2 21206 39712 21206 39712 0 _1090_
rlabel metal1 21666 41140 21666 41140 0 _1091_
rlabel metal1 18032 31450 18032 31450 0 _1092_
rlabel metal2 12282 33626 12282 33626 0 _1093_
rlabel metal2 13662 31212 13662 31212 0 _1094_
rlabel metal2 9614 30532 9614 30532 0 _1095_
rlabel metal2 21574 32504 21574 32504 0 _1096_
rlabel metal2 8326 30974 8326 30974 0 _1097_
rlabel metal1 13110 30906 13110 30906 0 _1098_
rlabel metal1 15272 29614 15272 29614 0 _1099_
rlabel metal1 12742 27914 12742 27914 0 _1100_
rlabel metal1 15272 28730 15272 28730 0 _1101_
rlabel metal1 14260 29274 14260 29274 0 _1102_
rlabel metal1 11270 30634 11270 30634 0 _1103_
rlabel metal1 13202 30702 13202 30702 0 _1104_
rlabel metal1 14168 30770 14168 30770 0 _1105_
rlabel metal1 15456 31382 15456 31382 0 _1106_
rlabel metal2 13846 31552 13846 31552 0 _1107_
rlabel metal2 13570 25568 13570 25568 0 _1108_
rlabel metal1 14582 31994 14582 31994 0 _1109_
rlabel metal1 14950 30906 14950 30906 0 _1110_
rlabel metal1 14352 32470 14352 32470 0 _1111_
rlabel metal1 13772 32402 13772 32402 0 _1112_
rlabel metal1 16514 31994 16514 31994 0 _1113_
rlabel metal1 13616 32198 13616 32198 0 _1114_
rlabel metal2 11270 28934 11270 28934 0 _1115_
rlabel metal1 10488 29478 10488 29478 0 _1116_
rlabel metal1 10626 28730 10626 28730 0 _1117_
rlabel metal2 11362 29750 11362 29750 0 _1118_
rlabel metal1 13662 28730 13662 28730 0 _1119_
rlabel metal1 12742 32470 12742 32470 0 _1120_
rlabel metal1 12696 30022 12696 30022 0 _1121_
rlabel metal2 13110 27540 13110 27540 0 _1122_
rlabel metal1 12144 29206 12144 29206 0 _1123_
rlabel metal2 12926 28900 12926 28900 0 _1124_
rlabel metal1 12696 29274 12696 29274 0 _1125_
rlabel metal1 11408 32878 11408 32878 0 _1126_
rlabel metal1 11868 30702 11868 30702 0 _1127_
rlabel metal1 11776 30294 11776 30294 0 _1128_
rlabel metal1 13478 30090 13478 30090 0 _1129_
rlabel metal2 13202 34833 13202 34833 0 _1130_
rlabel metal1 8418 28594 8418 28594 0 _1131_
rlabel metal1 18354 28730 18354 28730 0 _1132_
rlabel metal1 18040 28390 18040 28390 0 _1133_
rlabel metal1 18676 28662 18676 28662 0 _1134_
rlabel metal1 16284 30022 16284 30022 0 _1135_
rlabel viali 16322 30294 16322 30294 0 _1136_
rlabel metal1 16008 30362 16008 30362 0 _1137_
rlabel metal1 15594 29138 15594 29138 0 _1138_
rlabel metal1 15502 28968 15502 28968 0 _1139_
rlabel metal1 15791 29274 15791 29274 0 _1140_
rlabel metal1 16330 29104 16330 29104 0 _1141_
rlabel metal1 14076 27846 14076 27846 0 _1142_
rlabel metal1 14996 26962 14996 26962 0 _1143_
rlabel metal1 12650 28118 12650 28118 0 _1144_
rlabel metal1 12834 28084 12834 28084 0 _1145_
rlabel metal1 9108 27642 9108 27642 0 _1146_
rlabel metal1 8740 28526 8740 28526 0 _1147_
rlabel metal1 9354 28458 9354 28458 0 _1148_
rlabel metal1 9890 27438 9890 27438 0 _1149_
rlabel metal2 8326 28016 8326 28016 0 _1150_
rlabel metal1 9062 26996 9062 26996 0 _1151_
rlabel metal2 5474 28016 5474 28016 0 _1152_
rlabel metal2 5658 28254 5658 28254 0 _1153_
rlabel metal1 6670 28118 6670 28118 0 _1154_
rlabel metal1 4968 27438 4968 27438 0 _1155_
rlabel metal1 6578 28084 6578 28084 0 _1156_
rlabel metal1 6670 28730 6670 28730 0 _1157_
rlabel metal1 5888 29818 5888 29818 0 _1158_
rlabel metal1 6624 29138 6624 29138 0 _1159_
rlabel metal2 5198 30260 5198 30260 0 _1160_
rlabel metal1 6256 29274 6256 29274 0 _1161_
rlabel metal1 7268 35666 7268 35666 0 _1162_
rlabel metal1 6670 35496 6670 35496 0 _1163_
rlabel metal1 8050 35632 8050 35632 0 _1164_
rlabel metal1 7330 35734 7330 35734 0 _1165_
rlabel metal1 6992 35054 6992 35054 0 _1166_
rlabel metal1 9292 35258 9292 35258 0 _1167_
rlabel metal2 9522 35496 9522 35496 0 _1168_
rlabel metal1 9660 35258 9660 35258 0 _1169_
rlabel metal1 11500 35666 11500 35666 0 _1170_
rlabel metal1 10626 36346 10626 36346 0 _1171_
rlabel metal1 12650 36176 12650 36176 0 _1172_
rlabel metal1 12650 36584 12650 36584 0 _1173_
rlabel metal1 13570 36108 13570 36108 0 _1174_
rlabel metal2 12834 37060 12834 37060 0 _1175_
rlabel metal1 13662 36720 13662 36720 0 _1176_
rlabel metal1 13708 36278 13708 36278 0 _1177_
rlabel metal1 14076 35734 14076 35734 0 _1178_
rlabel metal1 39376 21114 39376 21114 0 _1179_
rlabel metal1 38916 20026 38916 20026 0 _1180_
rlabel metal1 37950 20468 37950 20468 0 _1181_
rlabel metal1 9338 3570 9338 3570 0 _1182_
rlabel metal1 9154 3706 9154 3706 0 _1183_
rlabel metal1 8878 4658 8878 4658 0 _1184_
rlabel metal2 38042 16694 38042 16694 0 _1185_
rlabel metal1 33626 8466 33626 8466 0 _1186_
rlabel metal1 34178 10098 34178 10098 0 _1187_
rlabel metal1 40710 30022 40710 30022 0 _1188_
rlabel metal1 11454 32946 11454 32946 0 _1189_
rlabel metal1 13386 44302 13386 44302 0 _1190_
rlabel metal2 12466 34238 12466 34238 0 _1191_
rlabel metal1 13938 34612 13938 34612 0 _1192_
rlabel via1 12942 33966 12942 33966 0 _1193_
rlabel metal1 13018 33864 13018 33864 0 _1194_
rlabel metal1 11868 33082 11868 33082 0 _1195_
rlabel metal1 7360 30634 7360 30634 0 _1196_
rlabel metal1 9798 31246 9798 31246 0 _1197_
rlabel metal1 10442 31790 10442 31790 0 _1198_
rlabel metal1 10575 32402 10575 32402 0 _1199_
rlabel metal1 9798 32198 9798 32198 0 _1200_
rlabel metal1 9062 31382 9062 31382 0 _1201_
rlabel metal1 8096 31790 8096 31790 0 _1202_
rlabel metal1 10166 31858 10166 31858 0 _1203_
rlabel metal1 10304 31314 10304 31314 0 _1204_
rlabel metal1 10391 31110 10391 31110 0 _1205_
rlabel metal1 10028 31246 10028 31246 0 _1206_
rlabel metal1 10488 32266 10488 32266 0 _1207_
rlabel metal1 10442 31450 10442 31450 0 _1208_
rlabel metal1 11224 31994 11224 31994 0 _1209_
rlabel metal2 14306 33864 14306 33864 0 _1210_
rlabel metal1 11086 33898 11086 33898 0 _1211_
rlabel metal1 13373 33422 13373 33422 0 _1212_
rlabel metal1 17802 32878 17802 32878 0 _1213_
rlabel metal1 18216 32810 18216 32810 0 _1214_
rlabel metal1 17756 33898 17756 33898 0 _1215_
rlabel metal1 17434 32334 17434 32334 0 _1216_
rlabel metal1 18446 32266 18446 32266 0 _1217_
rlabel metal1 17802 32436 17802 32436 0 _1218_
rlabel metal2 17066 33388 17066 33388 0 _1219_
rlabel metal1 16376 32538 16376 32538 0 _1220_
rlabel metal1 17204 32266 17204 32266 0 _1221_
rlabel metal1 16054 32300 16054 32300 0 _1222_
rlabel metal1 15962 32436 15962 32436 0 _1223_
rlabel via1 15778 33898 15778 33898 0 _1224_
rlabel metal1 16422 33286 16422 33286 0 _1225_
rlabel metal1 15456 32538 15456 32538 0 _1226_
rlabel metal2 15134 33388 15134 33388 0 _1227_
rlabel metal1 15042 32844 15042 32844 0 _1228_
rlabel metal1 15318 33014 15318 33014 0 _1229_
rlabel metal1 14766 33082 14766 33082 0 _1230_
rlabel metal1 15180 33354 15180 33354 0 _1231_
rlabel metal1 9660 31790 9660 31790 0 _1232_
rlabel metal1 9614 31926 9614 31926 0 _1233_
rlabel metal1 9798 31824 9798 31824 0 _1234_
rlabel metal1 11362 31790 11362 31790 0 _1235_
rlabel metal1 12834 33558 12834 33558 0 _1236_
rlabel metal2 17158 33813 17158 33813 0 _1237_
rlabel metal1 17521 33966 17521 33966 0 _1238_
rlabel metal1 16376 33626 16376 33626 0 _1239_
rlabel metal1 17388 33626 17388 33626 0 _1240_
rlabel metal1 14950 33592 14950 33592 0 _1241_
rlabel metal1 15686 34000 15686 34000 0 _1242_
rlabel metal1 17434 34068 17434 34068 0 _1243_
rlabel metal1 21114 33898 21114 33898 0 _1244_
rlabel metal1 41262 29682 41262 29682 0 _1245_
rlabel metal1 40434 28594 40434 28594 0 _1246_
rlabel metal1 39974 28934 39974 28934 0 _1247_
rlabel metal1 41078 29682 41078 29682 0 _1248_
rlabel metal1 39468 27642 39468 27642 0 _1249_
rlabel metal1 39836 28526 39836 28526 0 _1250_
rlabel metal2 38962 28356 38962 28356 0 _1251_
rlabel metal2 40158 30022 40158 30022 0 _1252_
rlabel metal1 39376 29274 39376 29274 0 _1253_
rlabel metal1 39284 28662 39284 28662 0 _1254_
rlabel via1 40798 29274 40798 29274 0 _1255_
rlabel metal1 41032 26418 41032 26418 0 _1256_
rlabel metal1 44574 29104 44574 29104 0 _1257_
rlabel metal1 43654 29002 43654 29002 0 _1258_
rlabel metal1 42596 26418 42596 26418 0 _1259_
rlabel metal1 44022 28084 44022 28084 0 _1260_
rlabel metal2 43930 28492 43930 28492 0 _1261_
rlabel metal1 43746 28084 43746 28084 0 _1262_
rlabel metal1 42918 26962 42918 26962 0 _1263_
rlabel metal1 43286 27914 43286 27914 0 _1264_
rlabel metal1 42642 26928 42642 26928 0 _1265_
rlabel metal1 42918 25908 42918 25908 0 _1266_
rlabel metal2 42458 26486 42458 26486 0 _1267_
rlabel metal2 42918 26554 42918 26554 0 _1268_
rlabel metal1 41262 26384 41262 26384 0 _1269_
rlabel metal1 43378 30770 43378 30770 0 _1270_
rlabel metal1 41722 29172 41722 29172 0 _1271_
rlabel metal1 41630 26350 41630 26350 0 _1272_
rlabel metal1 41170 26486 41170 26486 0 _1273_
rlabel metal2 41446 26180 41446 26180 0 _1274_
rlabel metal1 40572 26350 40572 26350 0 _1275_
rlabel metal1 40526 30362 40526 30362 0 _1276_
rlabel metal1 40526 28526 40526 28526 0 _1277_
rlabel metal1 39836 26282 39836 26282 0 _1278_
rlabel metal2 40250 26180 40250 26180 0 _1279_
rlabel metal1 39606 29682 39606 29682 0 _1280_
rlabel metal2 39882 29444 39882 29444 0 _1281_
rlabel metal1 39238 29716 39238 29716 0 _1282_
rlabel metal1 40066 26282 40066 26282 0 _1283_
rlabel metal1 39606 26350 39606 26350 0 _1284_
rlabel metal1 39882 17306 39882 17306 0 _1285_
rlabel metal1 38962 15334 38962 15334 0 _1286_
rlabel metal2 38778 14348 38778 14348 0 _1287_
rlabel metal1 32798 12716 32798 12716 0 _1288_
rlabel metal1 31188 13974 31188 13974 0 _1289_
rlabel metal1 32062 14042 32062 14042 0 _1290_
rlabel metal1 31924 14314 31924 14314 0 _1291_
rlabel metal1 35558 14246 35558 14246 0 _1292_
rlabel metal1 39514 15436 39514 15436 0 _1293_
rlabel metal1 23598 21046 23598 21046 0 _1294_
rlabel metal2 34822 12298 34822 12298 0 clk
rlabel metal2 14766 19115 14766 19115 0 clknet_0_clk
rlabel metal1 12144 20502 12144 20502 0 clknet_2_0__leaf_clk
rlabel metal1 20792 43282 20792 43282 0 clknet_2_1__leaf_clk
rlabel metal1 39882 14008 39882 14008 0 clknet_2_2__leaf_clk
rlabel metal1 35604 38998 35604 38998 0 clknet_2_3__leaf_clk
rlabel metal1 10718 17714 10718 17714 0 clknet_leaf_0_clk
rlabel metal1 21344 37978 21344 37978 0 clknet_leaf_10_clk
rlabel metal2 16790 34646 16790 34646 0 clknet_leaf_11_clk
rlabel metal1 20884 32946 20884 32946 0 clknet_leaf_12_clk
rlabel metal1 24288 26350 24288 26350 0 clknet_leaf_13_clk
rlabel metal1 27922 33558 27922 33558 0 clknet_leaf_14_clk
rlabel metal1 26036 35122 26036 35122 0 clknet_leaf_15_clk
rlabel metal2 24426 43792 24426 43792 0 clknet_leaf_16_clk
rlabel metal1 30130 43826 30130 43826 0 clknet_leaf_17_clk
rlabel metal1 37950 38726 37950 38726 0 clknet_leaf_18_clk
rlabel metal1 42182 37230 42182 37230 0 clknet_leaf_19_clk
rlabel metal1 17388 20910 17388 20910 0 clknet_leaf_1_clk
rlabel metal1 42780 34034 42780 34034 0 clknet_leaf_20_clk
rlabel metal1 43102 28730 43102 28730 0 clknet_leaf_21_clk
rlabel metal2 35696 32980 35696 32980 0 clknet_leaf_22_clk
rlabel metal2 27002 26146 27002 26146 0 clknet_leaf_23_clk
rlabel metal1 32660 17714 32660 17714 0 clknet_leaf_24_clk
rlabel metal1 34776 16626 34776 16626 0 clknet_leaf_25_clk
rlabel metal1 36938 22066 36938 22066 0 clknet_leaf_26_clk
rlabel metal1 44620 24242 44620 24242 0 clknet_leaf_27_clk
rlabel metal1 37812 13906 37812 13906 0 clknet_leaf_28_clk
rlabel metal1 42550 10098 42550 10098 0 clknet_leaf_29_clk
rlabel metal1 15502 27506 15502 27506 0 clknet_leaf_2_clk
rlabel metal1 34454 6766 34454 6766 0 clknet_leaf_30_clk
rlabel metal1 34914 9588 34914 9588 0 clknet_leaf_31_clk
rlabel metal1 32614 3570 32614 3570 0 clknet_leaf_32_clk
rlabel metal1 32890 13940 32890 13940 0 clknet_leaf_33_clk
rlabel metal1 18722 18734 18722 18734 0 clknet_leaf_34_clk
rlabel metal3 22747 12852 22747 12852 0 clknet_leaf_35_clk
rlabel metal1 16514 4522 16514 4522 0 clknet_leaf_36_clk
rlabel metal1 2622 5066 2622 5066 0 clknet_leaf_37_clk
rlabel metal1 7038 14518 7038 14518 0 clknet_leaf_38_clk
rlabel metal1 8970 23154 8970 23154 0 clknet_leaf_39_clk
rlabel metal1 9430 25738 9430 25738 0 clknet_leaf_3_clk
rlabel metal1 2024 31246 2024 31246 0 clknet_leaf_4_clk
rlabel metal1 3036 35598 3036 35598 0 clknet_leaf_5_clk
rlabel metal1 1748 40562 1748 40562 0 clknet_leaf_6_clk
rlabel metal1 10902 39406 10902 39406 0 clknet_leaf_7_clk
rlabel metal1 15962 41514 15962 41514 0 clknet_leaf_8_clk
rlabel metal1 20976 41582 20976 41582 0 clknet_leaf_9_clk
rlabel metal1 45080 44370 45080 44370 0 cs
rlabel metal1 42044 45934 42044 45934 0 gpio[0]
rlabel metal1 23920 45934 23920 45934 0 gpio[10]
rlabel metal3 820 8908 820 8908 0 gpio[11]
rlabel metal3 820 18428 820 18428 0 gpio[12]
rlabel metal1 44850 6324 44850 6324 0 gpio[13]
rlabel metal3 820 36788 820 36788 0 gpio[14]
rlabel metal1 45080 35054 45080 35054 0 gpio[15]
rlabel metal2 46 1588 46 1588 0 gpio[16]
rlabel metal2 8418 1027 8418 1027 0 gpio[1]
rlabel metal2 43838 1588 43838 1588 0 gpio[2]
rlabel metal2 17434 1588 17434 1588 0 gpio[3]
rlabel metal1 14950 45968 14950 45968 0 gpio[4]
rlabel metal1 45080 23698 45080 23698 0 gpio[5]
rlabel metal3 820 46308 820 46308 0 gpio[6]
rlabel metal2 33166 46393 33166 46393 0 gpio[7]
rlabel metal2 26450 1027 26450 1027 0 gpio[8]
rlabel metal3 820 27948 820 27948 0 gpio[9]
rlabel metal1 33304 5746 33304 5746 0 inputs.down.det_edge
rlabel metal1 33724 6970 33724 6970 0 inputs.down.ff_in
rlabel metal1 33350 9010 33350 9010 0 inputs.down.ff_out
rlabel metal1 34454 9486 34454 9486 0 inputs.down.in
rlabel metal1 16560 4182 16560 4182 0 inputs.frequency_lut.rng\[0\]
rlabel metal1 15042 4148 15042 4148 0 inputs.frequency_lut.rng\[1\]
rlabel metal1 13432 5678 13432 5678 0 inputs.frequency_lut.rng\[2\]
rlabel metal1 12558 6664 12558 6664 0 inputs.frequency_lut.rng\[3\]
rlabel metal1 19136 7446 19136 7446 0 inputs.frequency_lut.rng\[4\]
rlabel metal1 20148 15606 20148 15606 0 inputs.frequency_lut.rng\[5\]
rlabel metal2 37858 14212 37858 14212 0 inputs.key_encoder.mode_key
rlabel metal1 37720 13294 37720 13294 0 inputs.key_encoder.octave_key_up
rlabel metal1 33350 13838 33350 13838 0 inputs.key_encoder.sync_keys\[0\]
rlabel metal1 29624 15470 29624 15470 0 inputs.key_encoder.sync_keys\[10\]
rlabel metal2 10718 14297 10718 14297 0 inputs.key_encoder.sync_keys\[11\]
rlabel metal1 11270 13736 11270 13736 0 inputs.key_encoder.sync_keys\[12\]
rlabel metal1 24334 13838 24334 13838 0 inputs.key_encoder.sync_keys\[13\]
rlabel metal1 36340 13294 36340 13294 0 inputs.key_encoder.sync_keys\[14\]
rlabel metal1 35144 13294 35144 13294 0 inputs.key_encoder.sync_keys\[15\]
rlabel metal1 31326 13702 31326 13702 0 inputs.key_encoder.sync_keys\[1\]
rlabel metal1 30590 6766 30590 6766 0 inputs.key_encoder.sync_keys\[2\]
rlabel metal1 31280 5882 31280 5882 0 inputs.key_encoder.sync_keys\[3\]
rlabel metal1 29992 16082 29992 16082 0 inputs.key_encoder.sync_keys\[4\]
rlabel metal1 31786 15402 31786 15402 0 inputs.key_encoder.sync_keys\[5\]
rlabel metal1 31326 16014 31326 16014 0 inputs.key_encoder.sync_keys\[6\]
rlabel metal1 31694 14960 31694 14960 0 inputs.key_encoder.sync_keys\[7\]
rlabel metal1 29532 14994 29532 14994 0 inputs.key_encoder.sync_keys\[8\]
rlabel metal1 13386 17544 13386 17544 0 inputs.key_encoder.sync_keys\[9\]
rlabel metal1 35190 14450 35190 14450 0 inputs.keypad\[0\]
rlabel metal1 26266 43656 26266 43656 0 inputs.keypad\[10\]
rlabel metal1 7360 14042 7360 14042 0 inputs.keypad\[11\]
rlabel metal2 7314 16796 7314 16796 0 inputs.keypad\[12\]
rlabel metal1 8602 12954 8602 12954 0 inputs.keypad\[13\]
rlabel metal1 43700 12954 43700 12954 0 inputs.keypad\[14\]
rlabel metal1 8786 15538 8786 15538 0 inputs.keypad\[15\]
rlabel metal1 42527 13770 42527 13770 0 inputs.keypad\[16\]
rlabel metal1 26302 3706 26302 3706 0 inputs.keypad\[1\]
rlabel metal2 29854 4420 29854 4420 0 inputs.keypad\[2\]
rlabel metal2 27186 4726 27186 4726 0 inputs.keypad\[3\]
rlabel metal1 23874 17646 23874 17646 0 inputs.keypad\[4\]
rlabel metal2 36018 16490 36018 16490 0 inputs.keypad\[5\]
rlabel metal1 11638 17238 11638 17238 0 inputs.keypad\[6\]
rlabel metal1 32614 16184 32614 16184 0 inputs.keypad\[7\]
rlabel metal1 27278 3128 27278 3128 0 inputs.keypad\[8\]
rlabel metal2 10074 17816 10074 17816 0 inputs.keypad\[9\]
rlabel metal1 36110 14586 36110 14586 0 inputs.keypad_synchronizer.half_sync\[0\]
rlabel metal2 27784 35020 27784 35020 0 inputs.keypad_synchronizer.half_sync\[10\]
rlabel metal2 8786 14756 8786 14756 0 inputs.keypad_synchronizer.half_sync\[11\]
rlabel metal1 8970 16626 8970 16626 0 inputs.keypad_synchronizer.half_sync\[12\]
rlabel metal1 13708 13430 13708 13430 0 inputs.keypad_synchronizer.half_sync\[13\]
rlabel metal1 41124 13294 41124 13294 0 inputs.keypad_synchronizer.half_sync\[14\]
rlabel via2 10718 15691 10718 15691 0 inputs.keypad_synchronizer.half_sync\[15\]
rlabel metal1 39744 13362 39744 13362 0 inputs.keypad_synchronizer.half_sync\[16\]
rlabel metal1 28566 3604 28566 3604 0 inputs.keypad_synchronizer.half_sync\[1\]
rlabel metal1 31464 5338 31464 5338 0 inputs.keypad_synchronizer.half_sync\[2\]
rlabel metal1 29440 5882 29440 5882 0 inputs.keypad_synchronizer.half_sync\[3\]
rlabel metal1 28842 17306 28842 17306 0 inputs.keypad_synchronizer.half_sync\[4\]
rlabel metal1 37030 16082 37030 16082 0 inputs.keypad_synchronizer.half_sync\[5\]
rlabel metal2 21850 17306 21850 17306 0 inputs.keypad_synchronizer.half_sync\[6\]
rlabel metal1 34408 15538 34408 15538 0 inputs.keypad_synchronizer.half_sync\[7\]
rlabel metal1 29394 2482 29394 2482 0 inputs.keypad_synchronizer.half_sync\[8\]
rlabel metal1 11638 17850 11638 17850 0 inputs.keypad_synchronizer.half_sync\[9\]
rlabel metal1 39284 19754 39284 19754 0 inputs.mode_edge.det_edge
rlabel metal1 37996 17306 37996 17306 0 inputs.mode_edge.ff_in
rlabel metal1 38916 16626 38916 16626 0 inputs.mode_edge.ff_out
rlabel metal1 33258 5848 33258 5848 0 inputs.octave_fsm.octave_key_up
rlabel metal1 25346 5100 25346 5100 0 inputs.octave_fsm.state\[0\]
rlabel metal1 23736 5542 23736 5542 0 inputs.octave_fsm.state\[1\]
rlabel metal1 27002 6766 27002 6766 0 inputs.octave_fsm.state\[2\]
rlabel metal1 4876 3570 4876 3570 0 inputs.random_note_generator.feedback
rlabel metal1 5635 3434 5635 3434 0 inputs.random_note_generator.out\[0\]
rlabel metal1 8280 2482 8280 2482 0 inputs.random_note_generator.out\[10\]
rlabel metal1 8464 4046 8464 4046 0 inputs.random_note_generator.out\[11\]
rlabel metal2 7222 2621 7222 2621 0 inputs.random_note_generator.out\[12\]
rlabel metal1 9798 3570 9798 3570 0 inputs.random_note_generator.out\[13\]
rlabel metal1 11592 4046 11592 4046 0 inputs.random_note_generator.out\[14\]
rlabel metal1 12696 3026 12696 3026 0 inputs.random_note_generator.out\[15\]
rlabel metal1 4508 3162 4508 3162 0 inputs.random_note_generator.out\[1\]
rlabel metal1 1771 4794 1771 4794 0 inputs.random_note_generator.out\[2\]
rlabel metal1 4692 5134 4692 5134 0 inputs.random_note_generator.out\[3\]
rlabel metal1 5681 5678 5681 5678 0 inputs.random_note_generator.out\[4\]
rlabel metal1 5106 6426 5106 6426 0 inputs.random_note_generator.out\[5\]
rlabel metal1 8855 6426 8855 6426 0 inputs.random_note_generator.out\[6\]
rlabel metal1 6716 6834 6716 6834 0 inputs.random_note_generator.out\[7\]
rlabel metal1 9154 5678 9154 5678 0 inputs.random_note_generator.out\[8\]
rlabel metal1 10166 6222 10166 6222 0 inputs.random_note_generator.out\[9\]
rlabel metal1 34270 3468 34270 3468 0 inputs.random_update_clock.count\[0\]
rlabel metal1 42872 4522 42872 4522 0 inputs.random_update_clock.count\[10\]
rlabel metal2 43010 5576 43010 5576 0 inputs.random_update_clock.count\[11\]
rlabel metal1 42734 6324 42734 6324 0 inputs.random_update_clock.count\[12\]
rlabel metal1 41814 8976 41814 8976 0 inputs.random_update_clock.count\[13\]
rlabel metal1 42136 8262 42136 8262 0 inputs.random_update_clock.count\[14\]
rlabel metal1 41446 7242 41446 7242 0 inputs.random_update_clock.count\[15\]
rlabel metal1 36754 7990 36754 7990 0 inputs.random_update_clock.count\[16\]
rlabel metal1 37444 7310 37444 7310 0 inputs.random_update_clock.count\[17\]
rlabel metal1 37122 6834 37122 6834 0 inputs.random_update_clock.count\[18\]
rlabel metal1 38134 9452 38134 9452 0 inputs.random_update_clock.count\[19\]
rlabel metal1 34408 3366 34408 3366 0 inputs.random_update_clock.count\[1\]
rlabel metal1 38364 11254 38364 11254 0 inputs.random_update_clock.count\[20\]
rlabel metal1 38778 9573 38778 9573 0 inputs.random_update_clock.count\[21\]
rlabel metal1 39468 9486 39468 9486 0 inputs.random_update_clock.count\[22\]
rlabel metal2 34730 3706 34730 3706 0 inputs.random_update_clock.count\[2\]
rlabel metal1 34914 4454 34914 4454 0 inputs.random_update_clock.count\[3\]
rlabel metal1 37306 4182 37306 4182 0 inputs.random_update_clock.count\[4\]
rlabel metal1 36892 4454 36892 4454 0 inputs.random_update_clock.count\[5\]
rlabel metal1 37950 3502 37950 3502 0 inputs.random_update_clock.count\[6\]
rlabel metal1 38502 4760 38502 4760 0 inputs.random_update_clock.count\[7\]
rlabel metal1 41032 4794 41032 4794 0 inputs.random_update_clock.count\[8\]
rlabel metal1 42136 4046 42136 4046 0 inputs.random_update_clock.count\[9\]
rlabel metal1 31142 3162 31142 3162 0 inputs.random_update_clock.next_count\[0\]
rlabel metal1 42780 4046 42780 4046 0 inputs.random_update_clock.next_count\[10\]
rlabel metal1 43286 5338 43286 5338 0 inputs.random_update_clock.next_count\[11\]
rlabel metal2 43378 7820 43378 7820 0 inputs.random_update_clock.next_count\[12\]
rlabel metal1 41906 9690 41906 9690 0 inputs.random_update_clock.next_count\[13\]
rlabel metal1 43240 7786 43240 7786 0 inputs.random_update_clock.next_count\[14\]
rlabel metal1 39882 7786 39882 7786 0 inputs.random_update_clock.next_count\[15\]
rlabel metal1 35236 7310 35236 7310 0 inputs.random_update_clock.next_count\[16\]
rlabel metal1 38456 6154 38456 6154 0 inputs.random_update_clock.next_count\[17\]
rlabel metal1 35965 6970 35965 6970 0 inputs.random_update_clock.next_count\[18\]
rlabel metal1 36938 9486 36938 9486 0 inputs.random_update_clock.next_count\[19\]
rlabel via1 32699 3706 32699 3706 0 inputs.random_update_clock.next_count\[1\]
rlabel metal1 36846 10778 36846 10778 0 inputs.random_update_clock.next_count\[20\]
rlabel metal1 39882 10744 39882 10744 0 inputs.random_update_clock.next_count\[21\]
rlabel metal1 39928 10234 39928 10234 0 inputs.random_update_clock.next_count\[22\]
rlabel metal1 34086 2958 34086 2958 0 inputs.random_update_clock.next_count\[2\]
rlabel metal1 33580 4658 33580 4658 0 inputs.random_update_clock.next_count\[3\]
rlabel metal1 35650 3128 35650 3128 0 inputs.random_update_clock.next_count\[4\]
rlabel metal1 35965 4794 35965 4794 0 inputs.random_update_clock.next_count\[5\]
rlabel metal1 38824 2958 38824 2958 0 inputs.random_update_clock.next_count\[6\]
rlabel metal1 40388 4182 40388 4182 0 inputs.random_update_clock.next_count\[7\]
rlabel metal1 39790 4794 39790 4794 0 inputs.random_update_clock.next_count\[8\]
rlabel metal1 40618 3128 40618 3128 0 inputs.random_update_clock.next_count\[9\]
rlabel metal1 33902 6358 33902 6358 0 inputs.up.ff_in
rlabel metal1 34178 10778 34178 10778 0 inputs.up.ff_out
rlabel metal1 38318 20366 38318 20366 0 inputs.wavetype_fsm.next_state\[0\]
rlabel metal1 38916 21454 38916 21454 0 inputs.wavetype_fsm.next_state\[1\]
rlabel metal1 39468 20910 39468 20910 0 inputs.wavetype_fsm.state\[0\]
rlabel metal1 40020 22066 40020 22066 0 inputs.wavetype_fsm.state\[1\]
rlabel metal1 44482 44302 44482 44302 0 net1
rlabel metal1 9660 2618 9660 2618 0 net10
rlabel metal1 28658 45798 28658 45798 0 net100
rlabel metal1 11730 42330 11730 42330 0 net101
rlabel metal1 12558 42602 12558 42602 0 net102
rlabel metal1 14720 42874 14720 42874 0 net103
rlabel metal1 14076 42262 14076 42262 0 net104
rlabel metal2 41998 34748 41998 34748 0 net105
rlabel metal2 40986 35292 40986 35292 0 net106
rlabel metal1 8602 39066 8602 39066 0 net107
rlabel metal1 7130 40562 7130 40562 0 net108
rlabel metal1 16928 42330 16928 42330 0 net109
rlabel via2 30866 2907 30866 2907 0 net11
rlabel metal1 17578 42874 17578 42874 0 net110
rlabel metal1 14904 25262 14904 25262 0 net111
rlabel metal1 26818 44472 26818 44472 0 net112
rlabel metal1 26151 44370 26151 44370 0 net113
rlabel metal1 29532 44846 29532 44846 0 net114
rlabel metal2 38410 16150 38410 16150 0 net115
rlabel viali 8233 39406 8233 39406 0 net116
rlabel metal1 6808 39610 6808 39610 0 net117
rlabel metal1 5290 41446 5290 41446 0 net118
rlabel metal1 5842 42296 5842 42296 0 net119
rlabel metal1 21804 2618 21804 2618 0 net12
rlabel viali 21297 38930 21297 38930 0 net120
rlabel metal2 22034 39202 22034 39202 0 net121
rlabel metal1 41400 38182 41400 38182 0 net122
rlabel metal1 40289 36346 40289 36346 0 net123
rlabel metal2 6118 39406 6118 39406 0 net124
rlabel metal1 3910 40120 3910 40120 0 net125
rlabel metal1 32016 32946 32016 32946 0 net126
rlabel metal1 6578 40698 6578 40698 0 net127
rlabel metal1 7323 42874 7323 42874 0 net128
rlabel metal1 36846 33286 36846 33286 0 net129
rlabel metal1 14582 45798 14582 45798 0 net13
rlabel metal1 36708 32810 36708 32810 0 net130
rlabel metal1 23920 44778 23920 44778 0 net131
rlabel metal1 22218 43792 22218 43792 0 net132
rlabel metal1 30268 38318 30268 38318 0 net133
rlabel metal1 4738 40698 4738 40698 0 net134
rlabel metal2 1886 40290 1886 40290 0 net135
rlabel viali 23781 37842 23781 37842 0 net136
rlabel metal1 22816 38386 22816 38386 0 net137
rlabel metal2 38778 33218 38778 33218 0 net138
rlabel metal1 37996 33898 37996 33898 0 net139
rlabel metal1 40020 17034 40020 17034 0 net14
rlabel metal1 28520 23154 28520 23154 0 net140
rlabel metal1 22586 45594 22586 45594 0 net141
rlabel metal1 22264 44438 22264 44438 0 net142
rlabel metal1 40526 33626 40526 33626 0 net143
rlabel metal1 40526 33490 40526 33490 0 net144
rlabel metal1 23782 44404 23782 44404 0 net145
rlabel via1 4720 41106 4720 41106 0 net146
rlabel metal1 2944 41242 2944 41242 0 net147
rlabel metal1 38410 25262 38410 25262 0 net148
rlabel metal1 37812 26010 37812 26010 0 net149
rlabel metal2 1748 45540 1748 45540 0 net15
rlabel metal1 11960 40154 11960 40154 0 net150
rlabel metal1 11546 40086 11546 40086 0 net151
rlabel viali 8693 43282 8693 43282 0 net152
rlabel metal1 9200 42262 9200 42262 0 net153
rlabel metal2 36754 19516 36754 19516 0 net154
rlabel metal1 24518 36142 24518 36142 0 net155
rlabel metal1 25668 37298 25668 37298 0 net156
rlabel metal1 32430 2822 32430 2822 0 net157
rlabel metal1 33304 36142 33304 36142 0 net158
rlabel metal1 20056 41786 20056 41786 0 net159
rlabel metal2 31924 19380 31924 19380 0 net16
rlabel metal1 19734 42126 19734 42126 0 net160
rlabel metal1 32062 25942 32062 25942 0 net161
rlabel metal2 26542 40732 26542 40732 0 net162
rlabel metal1 42274 36788 42274 36788 0 net163
rlabel metal1 42780 36346 42780 36346 0 net164
rlabel metal1 33718 28594 33718 28594 0 net165
rlabel metal2 42458 7820 42458 7820 0 net166
rlabel metal1 42918 8602 42918 8602 0 net167
rlabel metal1 36018 7378 36018 7378 0 net168
rlabel metal1 32568 18394 32568 18394 0 net169
rlabel metal1 26680 2618 26680 2618 0 net17
rlabel metal1 30406 41650 30406 41650 0 net170
rlabel metal1 37858 32878 37858 32878 0 net171
rlabel metal1 37858 33422 37858 33422 0 net172
rlabel metal1 34316 18394 34316 18394 0 net173
rlabel metal1 32798 2414 32798 2414 0 net174
rlabel metal2 36202 27404 36202 27404 0 net175
rlabel metal1 36202 3502 36202 3502 0 net176
rlabel metal1 37168 9554 37168 9554 0 net177
rlabel metal1 36938 10608 36938 10608 0 net178
rlabel metal1 35374 29206 35374 29206 0 net179
rlabel metal1 1702 27846 1702 27846 0 net18
rlabel metal1 23920 42194 23920 42194 0 net180
rlabel metal1 32200 23222 32200 23222 0 net181
rlabel metal1 33902 31382 33902 31382 0 net182
rlabel metal1 39606 21522 39606 21522 0 net183
rlabel metal1 38180 21658 38180 21658 0 net184
rlabel metal1 32844 23766 32844 23766 0 net185
rlabel metal2 13938 35972 13938 35972 0 net186
rlabel metal1 40526 8500 40526 8500 0 net187
rlabel metal1 20700 35802 20700 35802 0 net188
rlabel metal1 19918 34578 19918 34578 0 net189
rlabel metal1 10902 12886 10902 12886 0 net19
rlabel metal1 35926 9588 35926 9588 0 net190
rlabel metal1 43378 5202 43378 5202 0 net191
rlabel metal2 34086 33082 34086 33082 0 net192
rlabel metal1 17618 28628 17618 28628 0 net193
rlabel metal1 34638 3434 34638 3434 0 net194
rlabel metal1 24196 31790 24196 31790 0 net195
rlabel metal1 41538 4250 41538 4250 0 net196
rlabel metal1 38962 37434 38962 37434 0 net197
rlabel metal1 33028 4114 33028 4114 0 net198
rlabel metal1 38180 35802 38180 35802 0 net199
rlabel metal1 41906 16184 41906 16184 0 net2
rlabel metal1 44436 15130 44436 15130 0 net20
rlabel metal1 36340 34646 36340 34646 0 net200
rlabel metal1 43010 37842 43010 37842 0 net201
rlabel metal1 42918 37298 42918 37298 0 net202
rlabel metal2 35650 22474 35650 22474 0 net203
rlabel metal1 22402 42228 22402 42228 0 net204
rlabel metal1 9384 33626 9384 33626 0 net205
rlabel metal1 9338 38930 9338 38930 0 net206
rlabel metal1 17112 45390 17112 45390 0 net207
rlabel metal1 18722 18938 18722 18938 0 net208
rlabel metal2 2438 33354 2438 33354 0 net209
rlabel metal1 37398 29036 37398 29036 0 net21
rlabel metal1 39698 38284 39698 38284 0 net210
rlabel metal1 26726 39066 26726 39066 0 net211
rlabel metal2 39330 3978 39330 3978 0 net212
rlabel metal1 38732 38794 38732 38794 0 net213
rlabel metal1 40480 38522 40480 38522 0 net214
rlabel metal2 13018 39508 13018 39508 0 net215
rlabel metal1 37444 3706 37444 3706 0 net216
rlabel metal1 22770 24786 22770 24786 0 net217
rlabel metal1 42550 25262 42550 25262 0 net218
rlabel metal1 44620 25262 44620 25262 0 net219
rlabel metal2 2714 4930 2714 4930 0 net22
rlabel metal1 25392 31790 25392 31790 0 net220
rlabel metal1 7958 32538 7958 32538 0 net221
rlabel metal1 33488 42670 33488 42670 0 net222
rlabel metal1 5980 37162 5980 37162 0 net223
rlabel metal2 14490 19924 14490 19924 0 net224
rlabel metal1 20470 35734 20470 35734 0 net225
rlabel metal1 13202 25874 13202 25874 0 net226
rlabel metal1 40894 24310 40894 24310 0 net227
rlabel metal1 2944 38930 2944 38930 0 net228
rlabel metal1 2438 37842 2438 37842 0 net229
rlabel metal2 12006 3978 12006 3978 0 net23
rlabel metal2 19642 43962 19642 43962 0 net230
rlabel metal2 11914 19890 11914 19890 0 net231
rlabel metal1 10120 45458 10120 45458 0 net232
rlabel metal1 8832 44846 8832 44846 0 net233
rlabel metal1 22632 34986 22632 34986 0 net234
rlabel metal1 21528 34578 21528 34578 0 net235
rlabel metal1 40158 22542 40158 22542 0 net236
rlabel metal2 24794 35360 24794 35360 0 net237
rlabel metal1 14582 44914 14582 44914 0 net238
rlabel metal1 16606 19482 16606 19482 0 net239
rlabel metal1 9798 12614 9798 12614 0 net24
rlabel metal1 16330 19380 16330 19380 0 net240
rlabel metal1 18492 22746 18492 22746 0 net241
rlabel metal1 18124 22202 18124 22202 0 net242
rlabel metal1 6670 33354 6670 33354 0 net243
rlabel metal1 5980 33490 5980 33490 0 net244
rlabel metal2 12558 23936 12558 23936 0 net245
rlabel metal1 11362 26282 11362 26282 0 net246
rlabel metal1 11316 24786 11316 24786 0 net247
rlabel metal2 24150 31552 24150 31552 0 net248
rlabel metal2 17066 37910 17066 37910 0 net249
rlabel metal1 10849 20910 10849 20910 0 net25
rlabel metal1 41722 37876 41722 37876 0 net250
rlabel metal1 16836 21658 16836 21658 0 net251
rlabel metal1 16330 21522 16330 21522 0 net252
rlabel metal1 18216 24242 18216 24242 0 net253
rlabel metal1 10902 44506 10902 44506 0 net254
rlabel metal1 17066 23834 17066 23834 0 net255
rlabel metal1 36018 39066 36018 39066 0 net256
rlabel metal2 15134 20706 15134 20706 0 net257
rlabel metal1 14490 18734 14490 18734 0 net258
rlabel metal1 3082 36890 3082 36890 0 net259
rlabel metal2 16054 21420 16054 21420 0 net26
rlabel metal1 34592 35802 34592 35802 0 net260
rlabel metal1 36938 37638 36938 37638 0 net261
rlabel metal2 18170 36652 18170 36652 0 net262
rlabel metal1 27646 41582 27646 41582 0 net263
rlabel metal2 26266 36652 26266 36652 0 net264
rlabel metal1 27876 34714 27876 34714 0 net265
rlabel metal1 26542 32946 26542 32946 0 net266
rlabel metal2 26542 31994 26542 31994 0 net267
rlabel metal1 42136 24786 42136 24786 0 net268
rlabel metal1 26036 29546 26036 29546 0 net269
rlabel metal1 32522 3434 32522 3434 0 net27
rlabel metal1 22356 29614 22356 29614 0 net270
rlabel metal2 3818 33558 3818 33558 0 net271
rlabel metal2 21758 29002 21758 29002 0 net272
rlabel metal1 12098 44506 12098 44506 0 net273
rlabel metal1 29716 36686 29716 36686 0 net274
rlabel metal2 12650 23970 12650 23970 0 net275
rlabel metal2 17986 26248 17986 26248 0 net276
rlabel metal1 4278 35156 4278 35156 0 net277
rlabel metal1 24104 25806 24104 25806 0 net278
rlabel metal1 18860 20434 18860 20434 0 net279
rlabel metal1 25392 13158 25392 13158 0 net28
rlabel metal1 18032 20434 18032 20434 0 net280
rlabel metal2 33350 42364 33350 42364 0 net281
rlabel metal1 6900 31926 6900 31926 0 net282
rlabel metal2 30682 41599 30682 41599 0 net283
rlabel metal1 38042 6392 38042 6392 0 net284
rlabel metal1 38272 6290 38272 6290 0 net285
rlabel metal1 21114 31892 21114 31892 0 net286
rlabel metal1 20470 31790 20470 31790 0 net287
rlabel metal1 34224 24922 34224 24922 0 net288
rlabel metal1 41538 31824 41538 31824 0 net289
rlabel metal2 33810 3808 33810 3808 0 net29
rlabel metal2 15870 32513 15870 32513 0 net290
rlabel metal1 18998 24378 18998 24378 0 net291
rlabel metal1 26680 21454 26680 21454 0 net292
rlabel metal1 36248 4182 36248 4182 0 net293
rlabel metal1 20010 33626 20010 33626 0 net294
rlabel metal1 35650 40154 35650 40154 0 net295
rlabel metal1 34224 8534 34224 8534 0 net296
rlabel metal1 24702 22542 24702 22542 0 net297
rlabel metal1 26588 28186 26588 28186 0 net298
rlabel metal1 35742 23664 35742 23664 0 net299
rlabel metal2 25070 44676 25070 44676 0 net3
rlabel metal1 42773 4182 42773 4182 0 net30
rlabel metal2 22954 36992 22954 36992 0 net300
rlabel metal1 18308 41446 18308 41446 0 net301
rlabel metal1 9246 41242 9246 41242 0 net302
rlabel metal1 38272 30226 38272 30226 0 net303
rlabel metal1 4462 37230 4462 37230 0 net304
rlabel metal1 35650 11050 35650 11050 0 net305
rlabel metal1 22632 26010 22632 26010 0 net306
rlabel metal1 37352 6970 37352 6970 0 net307
rlabel metal1 25530 24038 25530 24038 0 net308
rlabel metal1 4600 33626 4600 33626 0 net309
rlabel metal1 36524 8534 36524 8534 0 net31
rlabel metal1 22494 20570 22494 20570 0 net310
rlabel metal1 21344 18394 21344 18394 0 net311
rlabel metal1 20608 26282 20608 26282 0 net312
rlabel metal2 27094 30532 27094 30532 0 net313
rlabel metal1 41032 23834 41032 23834 0 net314
rlabel metal1 23920 20570 23920 20570 0 net315
rlabel metal1 21942 19380 21942 19380 0 net316
rlabel metal1 19412 21658 19412 21658 0 net317
rlabel metal1 21988 20434 21988 20434 0 net318
rlabel metal1 8004 2414 8004 2414 0 net319
rlabel metal1 25859 18326 25859 18326 0 net32
rlabel metal1 33074 23127 33074 23127 0 net33
rlabel metal1 38265 18326 38265 18326 0 net34
rlabel metal1 41446 15368 41446 15368 0 net35
rlabel metal1 35052 12954 35052 12954 0 net36
rlabel metal1 9936 34374 9936 34374 0 net37
rlabel metal2 19274 28254 19274 28254 0 net38
rlabel metal1 21022 34102 21022 34102 0 net39
rlabel metal1 4278 9146 4278 9146 0 net4
rlabel via2 21206 33915 21206 33915 0 net40
rlabel metal1 10403 40086 10403 40086 0 net41
rlabel metal2 5566 35904 5566 35904 0 net42
rlabel metal2 22678 44608 22678 44608 0 net43
rlabel metal1 20615 42194 20615 42194 0 net44
rlabel metal2 31878 26962 31878 26962 0 net45
rlabel metal1 27738 32953 27738 32953 0 net46
rlabel metal1 35597 32878 35597 32878 0 net47
rlabel metal2 43470 33320 43470 33320 0 net48
rlabel metal1 41814 32912 41814 32912 0 net49
rlabel metal2 6946 18190 6946 18190 0 net5
rlabel metal1 29302 36040 29302 36040 0 net50
rlabel metal2 25162 45016 25162 45016 0 net51
rlabel metal2 40710 39168 40710 39168 0 net52
rlabel metal1 43838 37155 43838 37155 0 net53
rlabel metal1 25990 42602 25990 42602 0 net54
rlabel metal1 22823 41582 22823 41582 0 net55
rlabel metal1 35144 14926 35144 14926 0 net56
rlabel metal1 37582 15538 37582 15538 0 net57
rlabel metal1 36432 13974 36432 13974 0 net58
rlabel metal1 9752 14450 9752 14450 0 net59
rlabel metal1 44390 12682 44390 12682 0 net6
rlabel metal1 9660 16422 9660 16422 0 net60
rlabel metal1 28007 16762 28007 16762 0 net61
rlabel metal1 42228 15538 42228 15538 0 net62
rlabel metal1 12144 17714 12144 17714 0 net63
rlabel metal1 30268 2618 30268 2618 0 net64
rlabel metal1 29900 5746 29900 5746 0 net65
rlabel metal1 29026 3706 29026 3706 0 net66
rlabel metal1 8105 3706 8105 3706 0 net67
rlabel metal1 8786 5882 8786 5882 0 net68
rlabel metal2 31694 6052 31694 6052 0 net69
rlabel metal1 4554 15946 4554 15946 0 net7
rlabel metal1 6578 6290 6578 6290 0 net70
rlabel metal1 7452 5610 7452 5610 0 net71
rlabel metal1 11270 3570 11270 3570 0 net72
rlabel metal1 4324 5338 4324 5338 0 net73
rlabel metal1 40480 12886 40480 12886 0 net74
rlabel metal2 10350 5644 10350 5644 0 net75
rlabel metal1 3450 4250 3450 4250 0 net76
rlabel metal1 39836 13294 39836 13294 0 net77
rlabel via2 17342 13821 17342 13821 0 net78
rlabel metal1 29118 17238 29118 17238 0 net79
rlabel metal2 44114 34136 44114 34136 0 net8
rlabel metal1 32062 14348 32062 14348 0 net80
rlabel metal1 8473 6970 8473 6970 0 net81
rlabel metal1 5980 3094 5980 3094 0 net82
rlabel metal1 6164 5882 6164 5882 0 net83
rlabel metal1 2714 5270 2714 5270 0 net84
rlabel metal1 7820 2958 7820 2958 0 net85
rlabel metal1 28198 30566 28198 30566 0 net86
rlabel metal2 9614 3876 9614 3876 0 net87
rlabel metal1 36892 11526 36892 11526 0 net88
rlabel metal1 7176 4046 7176 4046 0 net89
rlabel metal2 1610 7650 1610 7650 0 net9
rlabel metal1 43470 25466 43470 25466 0 net90
rlabel metal2 43286 26146 43286 26146 0 net91
rlabel metal1 20102 38998 20102 38998 0 net92
rlabel metal1 20562 39950 20562 39950 0 net93
rlabel metal1 36478 13362 36478 13362 0 net94
rlabel metal2 37306 15946 37306 15946 0 net95
rlabel metal1 39514 9690 39514 9690 0 net96
rlabel metal1 41308 10098 41308 10098 0 net97
rlabel metal1 17388 39066 17388 39066 0 net98
rlabel metal1 18170 40426 18170 40426 0 net99
rlabel metal1 6532 45934 6532 45934 0 nrst
rlabel metal1 29072 23630 29072 23630 0 outputs.div.a\[0\]
rlabel metal2 36754 27812 36754 27812 0 outputs.div.a\[10\]
rlabel metal1 36662 29138 36662 29138 0 outputs.div.a\[11\]
rlabel metal2 32706 28458 32706 28458 0 outputs.div.a\[12\]
rlabel metal1 35052 31790 35052 31790 0 outputs.div.a\[13\]
rlabel metal1 32246 33422 32246 33422 0 outputs.div.a\[14\]
rlabel metal1 33902 33626 33902 33626 0 outputs.div.a\[15\]
rlabel metal1 33258 36720 33258 36720 0 outputs.div.a\[16\]
rlabel metal1 34592 38726 34592 38726 0 outputs.div.a\[17\]
rlabel metal1 34408 38930 34408 38930 0 outputs.div.a\[18\]
rlabel metal2 35926 40188 35926 40188 0 outputs.div.a\[19\]
rlabel metal1 33258 22746 33258 22746 0 outputs.div.a\[1\]
rlabel metal1 35512 42738 35512 42738 0 outputs.div.a\[20\]
rlabel metal2 31878 43248 31878 43248 0 outputs.div.a\[21\]
rlabel metal1 30314 42704 30314 42704 0 outputs.div.a\[22\]
rlabel metal1 30912 42126 30912 42126 0 outputs.div.a\[23\]
rlabel metal1 30498 37876 30498 37876 0 outputs.div.a\[24\]
rlabel metal1 29578 36278 29578 36278 0 outputs.div.a\[25\]
rlabel metal1 37398 22542 37398 22542 0 outputs.div.a\[2\]
rlabel metal1 36018 19788 36018 19788 0 outputs.div.a\[3\]
rlabel metal1 36156 18938 36156 18938 0 outputs.div.a\[4\]
rlabel metal2 33626 18020 33626 18020 0 outputs.div.a\[5\]
rlabel metal2 30958 18020 30958 18020 0 outputs.div.a\[6\]
rlabel metal2 33442 23460 33442 23460 0 outputs.div.a\[7\]
rlabel metal1 32660 26418 32660 26418 0 outputs.div.a\[8\]
rlabel metal1 34914 25126 34914 25126 0 outputs.div.a\[9\]
rlabel viali 28198 41105 28198 41105 0 outputs.div.count\[0\]
rlabel metal1 26864 42194 26864 42194 0 outputs.div.count\[1\]
rlabel metal1 26864 41038 26864 41038 0 outputs.div.count\[2\]
rlabel metal1 27876 40018 27876 40018 0 outputs.div.count\[3\]
rlabel metal1 27278 39916 27278 39916 0 outputs.div.count\[4\]
rlabel metal1 30958 38998 30958 38998 0 outputs.div.div
rlabel metal1 22264 22066 22264 22066 0 outputs.div.divisor\[0\]
rlabel metal1 13662 23766 13662 23766 0 outputs.div.divisor\[10\]
rlabel metal2 20286 25602 20286 25602 0 outputs.div.divisor\[11\]
rlabel metal2 21390 26622 21390 26622 0 outputs.div.divisor\[12\]
rlabel metal1 21965 28458 21965 28458 0 outputs.div.divisor\[13\]
rlabel metal2 24886 29444 24886 29444 0 outputs.div.divisor\[14\]
rlabel metal1 25944 29614 25944 29614 0 outputs.div.divisor\[15\]
rlabel metal1 26404 28730 26404 28730 0 outputs.div.divisor\[16\]
rlabel metal2 23138 32198 23138 32198 0 outputs.div.divisor\[17\]
rlabel metal1 18814 22610 18814 22610 0 outputs.div.divisor\[1\]
rlabel metal1 19826 20468 19826 20468 0 outputs.div.divisor\[2\]
rlabel metal1 19090 21352 19090 21352 0 outputs.div.divisor\[3\]
rlabel metal1 20930 19414 20930 19414 0 outputs.div.divisor\[4\]
rlabel metal1 21666 18768 21666 18768 0 outputs.div.divisor\[5\]
rlabel metal1 19504 18734 19504 18734 0 outputs.div.divisor\[6\]
rlabel metal1 12052 19278 12052 19278 0 outputs.div.divisor\[7\]
rlabel metal1 12466 23562 12466 23562 0 outputs.div.divisor\[8\]
rlabel metal1 21574 23562 21574 23562 0 outputs.div.divisor\[9\]
rlabel metal1 29072 21998 29072 21998 0 outputs.div.m\[0\]
rlabel metal1 28888 25670 28888 25670 0 outputs.div.m\[10\]
rlabel metal2 26174 26112 26174 26112 0 outputs.div.m\[11\]
rlabel metal2 28474 27200 28474 27200 0 outputs.div.m\[12\]
rlabel metal1 28704 29002 28704 29002 0 outputs.div.m\[13\]
rlabel metal1 28888 30158 28888 30158 0 outputs.div.m\[14\]
rlabel metal1 29118 32402 29118 32402 0 outputs.div.m\[15\]
rlabel metal1 27738 32742 27738 32742 0 outputs.div.m\[16\]
rlabel metal1 29624 33286 29624 33286 0 outputs.div.m\[17\]
rlabel metal2 25162 21760 25162 21760 0 outputs.div.m\[1\]
rlabel metal1 25392 20774 25392 20774 0 outputs.div.m\[2\]
rlabel metal1 28658 21522 28658 21522 0 outputs.div.m\[3\]
rlabel metal1 29049 18258 29049 18258 0 outputs.div.m\[4\]
rlabel metal2 25622 18564 25622 18564 0 outputs.div.m\[5\]
rlabel metal1 25576 19142 25576 19142 0 outputs.div.m\[6\]
rlabel metal1 29440 19822 29440 19822 0 outputs.div.m\[7\]
rlabel metal2 26726 24344 26726 24344 0 outputs.div.m\[8\]
rlabel metal1 22724 24922 22724 24922 0 outputs.div.m\[9\]
rlabel metal1 33948 32810 33948 32810 0 outputs.div.next_div
rlabel metal1 27094 36890 27094 36890 0 outputs.div.next_start
rlabel metal1 23920 36890 23920 36890 0 outputs.div.oscillator_out\[0\]
rlabel metal1 5290 34578 5290 34578 0 outputs.div.oscillator_out\[10\]
rlabel metal1 5152 38386 5152 38386 0 outputs.div.oscillator_out\[11\]
rlabel metal2 5106 39508 5106 39508 0 outputs.div.oscillator_out\[12\]
rlabel metal1 9292 41106 9292 41106 0 outputs.div.oscillator_out\[13\]
rlabel metal2 11546 41956 11546 41956 0 outputs.div.oscillator_out\[14\]
rlabel metal1 13800 42330 13800 42330 0 outputs.div.oscillator_out\[15\]
rlabel metal2 17342 41956 17342 41956 0 outputs.div.oscillator_out\[16\]
rlabel metal1 20562 41718 20562 41718 0 outputs.div.oscillator_out\[17\]
rlabel metal1 22678 37094 22678 37094 0 outputs.div.oscillator_out\[1\]
rlabel metal1 21620 37094 21620 37094 0 outputs.div.oscillator_out\[2\]
rlabel metal1 19458 38862 19458 38862 0 outputs.div.oscillator_out\[3\]
rlabel metal1 16974 39610 16974 39610 0 outputs.div.oscillator_out\[4\]
rlabel metal2 12466 39780 12466 39780 0 outputs.div.oscillator_out\[5\]
rlabel metal1 8786 37978 8786 37978 0 outputs.div.oscillator_out\[6\]
rlabel metal2 8142 36176 8142 36176 0 outputs.div.oscillator_out\[7\]
rlabel metal1 4600 35802 4600 35802 0 outputs.div.oscillator_out\[8\]
rlabel metal2 2530 33116 2530 33116 0 outputs.div.oscillator_out\[9\]
rlabel metal2 37306 35292 37306 35292 0 outputs.div.q\[0\]
rlabel metal1 20746 39610 20746 39610 0 outputs.div.q\[10\]
rlabel metal2 18814 39406 18814 39406 0 outputs.div.q\[11\]
rlabel metal1 15088 40562 15088 40562 0 outputs.div.q\[12\]
rlabel via1 10074 39950 10074 39950 0 outputs.div.q\[13\]
rlabel metal1 8464 40562 8464 40562 0 outputs.div.q\[14\]
rlabel metal1 8142 40018 8142 40018 0 outputs.div.q\[15\]
rlabel metal1 5428 39950 5428 39950 0 outputs.div.q\[16\]
rlabel metal1 5382 40596 5382 40596 0 outputs.div.q\[17\]
rlabel metal1 3818 42194 3818 42194 0 outputs.div.q\[18\]
rlabel metal1 5382 41718 5382 41718 0 outputs.div.q\[19\]
rlabel metal1 41722 34612 41722 34612 0 outputs.div.q\[1\]
rlabel viali 6486 42194 6486 42194 0 outputs.div.q\[20\]
rlabel metal2 10718 42602 10718 42602 0 outputs.div.q\[21\]
rlabel metal1 13478 42602 13478 42602 0 outputs.div.q\[22\]
rlabel metal1 15410 41990 15410 41990 0 outputs.div.q\[23\]
rlabel metal1 17986 42772 17986 42772 0 outputs.div.q\[24\]
rlabel metal1 20930 42296 20930 42296 0 outputs.div.q\[25\]
rlabel metal1 26542 34544 26542 34544 0 outputs.div.q\[26\]
rlabel metal1 41860 37842 41860 37842 0 outputs.div.q\[2\]
rlabel metal2 42090 38012 42090 38012 0 outputs.div.q\[3\]
rlabel metal1 40572 38318 40572 38318 0 outputs.div.q\[4\]
rlabel metal1 39330 37196 39330 37196 0 outputs.div.q\[5\]
rlabel metal1 37950 35598 37950 35598 0 outputs.div.q\[6\]
rlabel metal1 36662 34646 36662 34646 0 outputs.div.q\[7\]
rlabel metal2 36202 36975 36202 36975 0 outputs.div.q\[8\]
rlabel metal1 23874 38522 23874 38522 0 outputs.div.q\[9\]
rlabel metal1 35650 33082 35650 33082 0 outputs.div.q_out\[0\]
rlabel metal1 42780 35122 42780 35122 0 outputs.div.q_out\[1\]
rlabel metal1 44344 37434 44344 37434 0 outputs.div.q_out\[2\]
rlabel metal2 44206 37332 44206 37332 0 outputs.div.q_out\[3\]
rlabel metal1 41906 36006 41906 36006 0 outputs.div.q_out\[4\]
rlabel metal1 40940 34510 40940 34510 0 outputs.div.q_out\[5\]
rlabel metal1 39744 34170 39744 34170 0 outputs.div.q_out\[6\]
rlabel metal1 38870 32946 38870 32946 0 outputs.div.q_out\[7\]
rlabel metal1 28658 38930 28658 38930 0 outputs.div.start
rlabel metal1 17066 23698 17066 23698 0 outputs.divider_buffer2\[0\]
rlabel metal1 13294 22746 13294 22746 0 outputs.divider_buffer2\[10\]
rlabel metal1 11730 25364 11730 25364 0 outputs.divider_buffer2\[11\]
rlabel metal1 12006 24786 12006 24786 0 outputs.divider_buffer2\[12\]
rlabel metal1 21735 27914 21735 27914 0 outputs.divider_buffer2\[13\]
rlabel metal1 23046 29274 23046 29274 0 outputs.divider_buffer2\[14\]
rlabel metal1 26082 31178 26082 31178 0 outputs.divider_buffer2\[15\]
rlabel metal1 26174 30804 26174 30804 0 outputs.divider_buffer2\[16\]
rlabel metal2 24242 30396 24242 30396 0 outputs.divider_buffer2\[17\]
rlabel metal1 19228 22610 19228 22610 0 outputs.divider_buffer2\[1\]
rlabel metal1 18584 20570 18584 20570 0 outputs.divider_buffer2\[2\]
rlabel metal1 16836 21862 16836 21862 0 outputs.divider_buffer2\[3\]
rlabel metal1 17572 18938 17572 18938 0 outputs.divider_buffer2\[4\]
rlabel metal1 14720 19482 14720 19482 0 outputs.divider_buffer2\[5\]
rlabel metal1 13846 19958 13846 19958 0 outputs.divider_buffer2\[6\]
rlabel metal1 11684 18802 11684 18802 0 outputs.divider_buffer2\[7\]
rlabel metal1 11454 23290 11454 23290 0 outputs.divider_buffer2\[8\]
rlabel metal2 16238 25364 16238 25364 0 outputs.divider_buffer2\[9\]
rlabel metal1 16882 25466 16882 25466 0 outputs.divider_buffer\[0\]
rlabel metal2 9798 23392 9798 23392 0 outputs.divider_buffer\[10\]
rlabel metal1 8648 31314 8648 31314 0 outputs.divider_buffer\[11\]
rlabel metal1 9292 25670 9292 25670 0 outputs.divider_buffer\[12\]
rlabel metal1 20010 31926 20010 31926 0 outputs.divider_buffer\[13\]
rlabel metal1 21160 31790 21160 31790 0 outputs.divider_buffer\[14\]
rlabel metal1 20838 31722 20838 31722 0 outputs.divider_buffer\[15\]
rlabel metal2 24426 33847 24426 33847 0 outputs.divider_buffer\[16\]
rlabel metal1 21942 31178 21942 31178 0 outputs.divider_buffer\[17\]
rlabel metal1 18722 25466 18722 25466 0 outputs.divider_buffer\[1\]
rlabel metal1 18492 26554 18492 26554 0 outputs.divider_buffer\[2\]
rlabel metal1 16284 32402 16284 32402 0 outputs.divider_buffer\[3\]
rlabel metal1 16008 20570 16008 20570 0 outputs.divider_buffer\[4\]
rlabel metal1 14536 21658 14536 21658 0 outputs.divider_buffer\[5\]
rlabel metal1 13800 21114 13800 21114 0 outputs.divider_buffer\[6\]
rlabel metal1 11362 21114 11362 21114 0 outputs.divider_buffer\[7\]
rlabel metal1 10672 33422 10672 33422 0 outputs.divider_buffer\[8\]
rlabel metal2 14950 29410 14950 29410 0 outputs.divider_buffer\[9\]
rlabel via1 42834 24854 42834 24854 0 outputs.output_gen.count\[0\]
rlabel metal1 43976 26962 43976 26962 0 outputs.output_gen.count\[1\]
rlabel metal1 42642 26282 42642 26282 0 outputs.output_gen.count\[2\]
rlabel metal1 42136 24242 42136 24242 0 outputs.output_gen.count\[3\]
rlabel metal2 41170 26078 41170 26078 0 outputs.output_gen.count\[4\]
rlabel metal1 39974 25840 39974 25840 0 outputs.output_gen.count\[5\]
rlabel metal1 39698 25840 39698 25840 0 outputs.output_gen.count\[6\]
rlabel metal1 39698 26418 39698 26418 0 outputs.output_gen.count\[7\]
rlabel metal2 43286 23460 43286 23460 0 outputs.output_gen.next_count\[0\]
rlabel metal1 43470 25874 43470 25874 0 outputs.output_gen.next_count\[1\]
rlabel metal2 44390 24684 44390 24684 0 outputs.output_gen.next_count\[2\]
rlabel metal1 41354 24072 41354 24072 0 outputs.output_gen.next_count\[3\]
rlabel metal1 40526 22644 40526 22644 0 outputs.output_gen.next_count\[4\]
rlabel metal1 39054 23800 39054 23800 0 outputs.output_gen.next_count\[5\]
rlabel metal1 37713 24378 37713 24378 0 outputs.output_gen.next_count\[6\]
rlabel metal1 38134 25466 38134 25466 0 outputs.output_gen.next_count\[7\]
rlabel metal2 41630 15844 41630 15844 0 outputs.output_gen.pwm_ff
rlabel metal1 39928 15402 39928 15402 0 outputs.output_gen.pwm_unff
rlabel metal1 43746 15674 43746 15674 0 outputs.pwm_output
rlabel metal1 27646 44166 27646 44166 0 outputs.sample_rate.count\[0\]
rlabel metal1 29026 45254 29026 45254 0 outputs.sample_rate.count\[1\]
rlabel metal1 28060 45050 28060 45050 0 outputs.sample_rate.count\[2\]
rlabel metal1 25760 44302 25760 44302 0 outputs.sample_rate.count\[3\]
rlabel metal1 23552 44506 23552 44506 0 outputs.sample_rate.count\[4\]
rlabel metal1 23506 44846 23506 44846 0 outputs.sample_rate.count\[5\]
rlabel metal1 23138 42738 23138 42738 0 outputs.sample_rate.count\[6\]
rlabel metal1 23276 41786 23276 41786 0 outputs.sample_rate.count\[7\]
rlabel metal1 27416 44438 27416 44438 0 outputs.sample_rate.next_count\[0\]
rlabel metal1 29532 45050 29532 45050 0 outputs.sample_rate.next_count\[1\]
rlabel metal2 26542 44642 26542 44642 0 outputs.sample_rate.next_count\[2\]
rlabel metal1 24380 44914 24380 44914 0 outputs.sample_rate.next_count\[3\]
rlabel metal2 22034 45499 22034 45499 0 outputs.sample_rate.next_count\[4\]
rlabel metal2 22218 44438 22218 44438 0 outputs.sample_rate.next_count\[5\]
rlabel metal1 21804 42330 21804 42330 0 outputs.sample_rate.next_count\[6\]
rlabel metal1 21528 41242 21528 41242 0 outputs.sample_rate.next_count\[7\]
rlabel metal2 43378 30532 43378 30532 0 outputs.scaled_buffer\[0\]
rlabel metal1 42688 33830 42688 33830 0 outputs.scaled_buffer\[1\]
rlabel metal1 44206 31178 44206 31178 0 outputs.scaled_buffer\[2\]
rlabel metal1 43010 33524 43010 33524 0 outputs.scaled_buffer\[3\]
rlabel metal2 41262 31994 41262 31994 0 outputs.scaled_buffer\[4\]
rlabel metal1 40940 33082 40940 33082 0 outputs.scaled_buffer\[5\]
rlabel metal2 39514 31552 39514 31552 0 outputs.scaled_buffer\[6\]
rlabel metal1 39376 30158 39376 30158 0 outputs.scaled_buffer\[7\]
rlabel metal1 19550 33456 19550 33456 0 outputs.shaper.count\[0\]
rlabel metal1 7268 31858 7268 31858 0 outputs.shaper.count\[10\]
rlabel metal1 3588 36686 3588 36686 0 outputs.shaper.count\[11\]
rlabel metal1 6716 34918 6716 34918 0 outputs.shaper.count\[12\]
rlabel metal1 10350 32368 10350 32368 0 outputs.shaper.count\[13\]
rlabel metal1 13156 44914 13156 44914 0 outputs.shaper.count\[14\]
rlabel metal1 13156 44166 13156 44166 0 outputs.shaper.count\[15\]
rlabel metal1 16974 45458 16974 45458 0 outputs.shaper.count\[16\]
rlabel metal1 18584 43622 18584 43622 0 outputs.shaper.count\[17\]
rlabel metal2 22034 33286 22034 33286 0 outputs.shaper.count\[1\]
rlabel metal1 20654 34170 20654 34170 0 outputs.shaper.count\[2\]
rlabel metal1 18722 35054 18722 35054 0 outputs.shaper.count\[3\]
rlabel metal2 16054 36550 16054 36550 0 outputs.shaper.count\[4\]
rlabel metal1 14766 40154 14766 40154 0 outputs.shaper.count\[5\]
rlabel metal2 11270 38046 11270 38046 0 outputs.shaper.count\[6\]
rlabel metal1 9936 33830 9936 33830 0 outputs.shaper.count\[7\]
rlabel metal2 4186 30617 4186 30617 0 outputs.shaper.count\[8\]
rlabel metal2 3266 31246 3266 31246 0 outputs.shaper.count\[9\]
rlabel metal1 21620 36006 21620 36006 0 outputs.sig_gen.count\[0\]
rlabel metal1 5014 33354 5014 33354 0 outputs.sig_gen.count\[10\]
rlabel metal1 4692 37094 4692 37094 0 outputs.sig_gen.count\[11\]
rlabel metal1 7728 35666 7728 35666 0 outputs.sig_gen.count\[12\]
rlabel metal1 9338 36074 9338 36074 0 outputs.sig_gen.count\[13\]
rlabel metal2 12466 32946 12466 32946 0 outputs.sig_gen.count\[14\]
rlabel metal1 13478 41446 13478 41446 0 outputs.sig_gen.count\[15\]
rlabel metal1 15778 37978 15778 37978 0 outputs.sig_gen.count\[16\]
rlabel metal1 14398 36346 14398 36346 0 outputs.sig_gen.count\[17\]
rlabel metal2 21298 29359 21298 29359 0 outputs.sig_gen.count\[1\]
rlabel metal1 18492 31858 18492 31858 0 outputs.sig_gen.count\[2\]
rlabel metal1 18400 37230 18400 37230 0 outputs.sig_gen.count\[3\]
rlabel metal2 16422 36210 16422 36210 0 outputs.sig_gen.count\[4\]
rlabel metal1 13984 31178 13984 31178 0 outputs.sig_gen.count\[5\]
rlabel metal1 13064 33014 13064 33014 0 outputs.sig_gen.count\[6\]
rlabel metal1 7820 32334 7820 32334 0 outputs.sig_gen.count\[7\]
rlabel metal1 4876 34918 4876 34918 0 outputs.sig_gen.count\[8\]
rlabel metal1 12512 28050 12512 28050 0 outputs.sig_gen.count\[9\]
rlabel metal1 17940 28050 17940 28050 0 outputs.sig_gen.next_count\[0\]
rlabel metal1 4462 30328 4462 30328 0 outputs.sig_gen.next_count\[10\]
rlabel metal1 6164 29546 6164 29546 0 outputs.sig_gen.next_count\[11\]
rlabel metal1 6716 35258 6716 35258 0 outputs.sig_gen.next_count\[12\]
rlabel metal1 9476 35598 9476 35598 0 outputs.sig_gen.next_count\[13\]
rlabel metal1 11040 36210 11040 36210 0 outputs.sig_gen.next_count\[14\]
rlabel metal1 12512 37434 12512 37434 0 outputs.sig_gen.next_count\[15\]
rlabel metal1 14168 36890 14168 36890 0 outputs.sig_gen.next_count\[16\]
rlabel metal1 14904 35530 14904 35530 0 outputs.sig_gen.next_count\[17\]
rlabel metal1 19504 28458 19504 28458 0 outputs.sig_gen.next_count\[1\]
rlabel metal1 16882 30770 16882 30770 0 outputs.sig_gen.next_count\[2\]
rlabel metal1 16974 29240 16974 29240 0 outputs.sig_gen.next_count\[3\]
rlabel metal1 14766 27098 14766 27098 0 outputs.sig_gen.next_count\[4\]
rlabel metal2 12834 27744 12834 27744 0 outputs.sig_gen.next_count\[5\]
rlabel metal1 10672 27574 10672 27574 0 outputs.sig_gen.next_count\[6\]
rlabel metal1 9016 27098 9016 27098 0 outputs.sig_gen.next_count\[7\]
rlabel metal2 4830 27812 4830 27812 0 outputs.sig_gen.next_count\[8\]
rlabel metal1 6808 27030 6808 27030 0 outputs.sig_gen.next_count\[9\]
rlabel metal1 25576 35802 25576 35802 0 outputs.signal_buffer2\[0\]
rlabel metal1 6118 33082 6118 33082 0 outputs.signal_buffer2\[10\]
rlabel metal1 3496 38522 3496 38522 0 outputs.signal_buffer2\[11\]
rlabel metal1 6394 37298 6394 37298 0 outputs.signal_buffer2\[12\]
rlabel metal1 9706 44472 9706 44472 0 outputs.signal_buffer2\[13\]
rlabel metal1 9982 43860 9982 43860 0 outputs.signal_buffer2\[14\]
rlabel metal1 14674 45356 14674 45356 0 outputs.signal_buffer2\[15\]
rlabel metal1 17342 44472 17342 44472 0 outputs.signal_buffer2\[16\]
rlabel metal1 20378 44268 20378 44268 0 outputs.signal_buffer2\[17\]
rlabel metal1 23322 34714 23322 34714 0 outputs.signal_buffer2\[1\]
rlabel metal1 21206 35666 21206 35666 0 outputs.signal_buffer2\[2\]
rlabel metal1 19044 37978 19044 37978 0 outputs.signal_buffer2\[3\]
rlabel metal1 17388 38522 17388 38522 0 outputs.signal_buffer2\[4\]
rlabel metal1 13938 38930 13938 38930 0 outputs.signal_buffer2\[5\]
rlabel metal1 9108 38522 9108 38522 0 outputs.signal_buffer2\[6\]
rlabel metal1 8694 34170 8694 34170 0 outputs.signal_buffer2\[7\]
rlabel metal1 3128 32402 3128 32402 0 outputs.signal_buffer2\[8\]
rlabel metal1 3082 32538 3082 32538 0 outputs.signal_buffer2\[9\]
rlabel via2 44758 16405 44758 16405 0 pwm
<< properties >>
string FIXED_BBOX 0 0 46337 48481
<< end >>
