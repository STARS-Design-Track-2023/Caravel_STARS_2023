magic
tech sky130A
magscale 1 2
timestamp 1691548399
<< obsli1 >>
rect 1104 2159 62376 63121
<< obsm1 >>
rect 14 2128 62454 63152
<< metal2 >>
rect 5170 64909 5226 65709
rect 12254 64909 12310 65709
rect 19338 64909 19394 65709
rect 25778 64909 25834 65709
rect 32862 64909 32918 65709
rect 39302 64909 39358 65709
rect 46386 64909 46442 65709
rect 53470 64909 53526 65709
rect 59910 64909 59966 65709
rect 18 0 74 800
rect 6458 0 6514 800
rect 13542 0 13598 800
rect 19982 0 20038 800
rect 27066 0 27122 800
rect 33506 0 33562 800
rect 40590 0 40646 800
rect 47674 0 47730 800
rect 54114 0 54170 800
rect 61198 0 61254 800
<< obsm2 >>
rect 20 64853 5114 64909
rect 5282 64853 12198 64909
rect 12366 64853 19282 64909
rect 19450 64853 25722 64909
rect 25890 64853 32806 64909
rect 32974 64853 39246 64909
rect 39414 64853 46330 64909
rect 46498 64853 53414 64909
rect 53582 64853 59854 64909
rect 60022 64853 62450 64909
rect 20 856 62450 64853
rect 130 734 6402 856
rect 6570 734 13486 856
rect 13654 734 19926 856
rect 20094 734 27010 856
rect 27178 734 33450 856
rect 33618 734 40534 856
rect 40702 734 47618 856
rect 47786 734 54058 856
rect 54226 734 61142 856
rect 61310 734 62450 856
<< metal3 >>
rect 0 64608 800 64728
rect 62765 61888 63565 62008
rect 0 57128 800 57248
rect 62765 55088 63565 55208
rect 0 50328 800 50448
rect 62765 47608 63565 47728
rect 0 42848 800 42968
rect 62765 40128 63565 40248
rect 0 35368 800 35488
rect 62765 33328 63565 33448
rect 0 28568 800 28688
rect 62765 25848 63565 25968
rect 0 21088 800 21208
rect 62765 19048 63565 19168
rect 0 14288 800 14408
rect 62765 11568 63565 11688
rect 0 6808 800 6928
rect 62765 4088 63565 4208
<< obsm3 >>
rect 880 64528 62765 64701
rect 798 62088 62765 64528
rect 798 61808 62685 62088
rect 798 57328 62765 61808
rect 880 57048 62765 57328
rect 798 55288 62765 57048
rect 798 55008 62685 55288
rect 798 50528 62765 55008
rect 880 50248 62765 50528
rect 798 47808 62765 50248
rect 798 47528 62685 47808
rect 798 43048 62765 47528
rect 880 42768 62765 43048
rect 798 40328 62765 42768
rect 798 40048 62685 40328
rect 798 35568 62765 40048
rect 880 35288 62765 35568
rect 798 33528 62765 35288
rect 798 33248 62685 33528
rect 798 28768 62765 33248
rect 880 28488 62765 28768
rect 798 26048 62765 28488
rect 798 25768 62685 26048
rect 798 21288 62765 25768
rect 880 21008 62765 21288
rect 798 19248 62765 21008
rect 798 18968 62685 19248
rect 798 14488 62765 18968
rect 880 14208 62765 14488
rect 798 11768 62765 14208
rect 798 11488 62685 11768
rect 798 7008 62765 11488
rect 880 6728 62765 7008
rect 798 4288 62765 6728
rect 798 4008 62685 4288
rect 798 2143 62765 4008
<< metal4 >>
rect 4208 2128 4528 63152
rect 4868 2128 5188 63152
rect 34928 2128 35248 63152
rect 35588 2128 35908 63152
<< obsm4 >>
rect 12203 20299 34848 62389
rect 35328 20299 35508 62389
rect 35988 20299 56061 62389
<< metal5 >>
rect 1056 36642 62424 36962
rect 1056 35982 62424 36302
rect 1056 6006 62424 6326
rect 1056 5346 62424 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 63152 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 63152 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 62424 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 62424 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 63152 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 63152 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 62424 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 62424 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 33506 0 33562 800 6 bottom_row[0]
port 3 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 bottom_row[1]
port 4 nsew signal output
rlabel metal2 s 12254 64909 12310 65709 6 bottom_row[2]
port 5 nsew signal output
rlabel metal2 s 53470 64909 53526 65709 6 bottom_row[3]
port 6 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 bottom_row[4]
port 7 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 bottom_row[5]
port 8 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 bottom_row[6]
port 9 nsew signal output
rlabel metal2 s 46386 64909 46442 65709 6 button[0]
port 10 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 button[1]
port 11 nsew signal input
rlabel metal3 s 62765 40128 63565 40248 6 button[2]
port 12 nsew signal input
rlabel metal2 s 39302 64909 39358 65709 6 button[3]
port 13 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 chip_select
port 14 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 clk
port 15 nsew signal input
rlabel metal3 s 62765 4088 63565 4208 6 green_disp
port 16 nsew signal output
rlabel metal3 s 62765 33328 63565 33448 6 n_rst
port 17 nsew signal input
rlabel metal3 s 62765 47608 63565 47728 6 red_disp
port 18 nsew signal output
rlabel metal2 s 18 0 74 800 6 ss0[0]
port 19 nsew signal output
rlabel metal2 s 32862 64909 32918 65709 6 ss0[1]
port 20 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 ss0[2]
port 21 nsew signal output
rlabel metal2 s 19338 64909 19394 65709 6 ss0[3]
port 22 nsew signal output
rlabel metal2 s 5170 64909 5226 65709 6 ss0[4]
port 23 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 ss0[5]
port 24 nsew signal output
rlabel metal2 s 59910 64909 59966 65709 6 ss0[6]
port 25 nsew signal output
rlabel metal3 s 62765 11568 63565 11688 6 ss1[0]
port 26 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 ss1[1]
port 27 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 ss1[2]
port 28 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 ss1[3]
port 29 nsew signal output
rlabel metal3 s 62765 19048 63565 19168 6 ss1[4]
port 30 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 ss1[5]
port 31 nsew signal output
rlabel metal3 s 62765 55088 63565 55208 6 ss1[6]
port 32 nsew signal output
rlabel metal3 s 62765 61888 63565 62008 6 top_row[0]
port 33 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 top_row[1]
port 34 nsew signal output
rlabel metal2 s 25778 64909 25834 65709 6 top_row[2]
port 35 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 top_row[3]
port 36 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 top_row[4]
port 37 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 top_row[5]
port 38 nsew signal output
rlabel metal3 s 62765 25848 63565 25968 6 top_row[6]
port 39 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 63565 65709
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10142850
string GDS_FILE /home/designer-25/CUP/openlane/GuitarVillans/runs/23_08_08_19_26/results/signoff/Guitar_Villains.magic.gds
string GDS_START 1091252
<< end >>

