// This is the unpowered netlist.
module z23 (clk,
    interrupt_gpio_in,
    memory_wr,
    nrst,
    keypad_input,
    memory_address_out,
    memory_data_in,
    memory_data_out,
    programmable_gpio_in,
    programmable_gpio_out,
    programmable_gpio_wr,
    ss0,
    ss1,
    ss2,
    ss3,
    ss4,
    ss5,
    ss6,
    ss7);
 input clk;
 input interrupt_gpio_in;
 output memory_wr;
 input nrst;
 input [15:0] keypad_input;
 output [15:0] memory_address_out;
 input [7:0] memory_data_in;
 output [7:0] memory_data_out;
 input [7:0] programmable_gpio_in;
 output [7:0] programmable_gpio_out;
 output [7:0] programmable_gpio_wr;
 output [7:0] ss0;
 output [7:0] ss1;
 output [7:0] ss2;
 output [7:0] ss3;
 output [7:0] ss4;
 output [7:0] ss5;
 output [7:0] ss6;
 output [7:0] ss7;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire \alu.Cin ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \cu.alu_f[1] ;
 wire \cu.alu_f[2] ;
 wire \cu.alu_f[3] ;
 wire \cu.alu_f[4] ;
 wire \cu.alu_f[5] ;
 wire \cu.alu_f[6] ;
 wire \cu.alu_f[7] ;
 wire \cu.id.alu_opcode[0] ;
 wire \cu.id.alu_opcode[1] ;
 wire \cu.id.alu_opcode[3] ;
 wire \cu.id.can_be_interrupted ;
 wire \cu.id.cb_opcode_x[0] ;
 wire \cu.id.cb_opcode_x[1] ;
 wire \cu.id.cb_opcode_y[0] ;
 wire \cu.id.cb_opcode_y[1] ;
 wire \cu.id.cb_opcode_y[2] ;
 wire \cu.id.cb_opcode_z[0] ;
 wire \cu.id.cb_opcode_z[1] ;
 wire \cu.id.cb_opcode_z[2] ;
 wire \cu.id.imm_i[10] ;
 wire \cu.id.imm_i[11] ;
 wire \cu.id.imm_i[12] ;
 wire \cu.id.imm_i[13] ;
 wire \cu.id.imm_i[14] ;
 wire \cu.id.imm_i[15] ;
 wire \cu.id.imm_i[8] ;
 wire \cu.id.imm_i[9] ;
 wire \cu.id.interrupt_requested ;
 wire \cu.id.is_halted ;
 wire \cu.id.is_interrupted ;
 wire \cu.id.opcode[0] ;
 wire \cu.id.opcode[1] ;
 wire \cu.id.opcode[2] ;
 wire \cu.id.opcode[6] ;
 wire \cu.id.opcode[7] ;
 wire \cu.id.starting_int_service ;
 wire \cu.id.state[0] ;
 wire \cu.id.state[1] ;
 wire \cu.id.state[2] ;
 wire \cu.ir.idx[0] ;
 wire \cu.ir.idx[1] ;
 wire \cu.pc.pc_o[0] ;
 wire \cu.pc.pc_o[10] ;
 wire \cu.pc.pc_o[11] ;
 wire \cu.pc.pc_o[12] ;
 wire \cu.pc.pc_o[13] ;
 wire \cu.pc.pc_o[14] ;
 wire \cu.pc.pc_o[15] ;
 wire \cu.pc.pc_o[1] ;
 wire \cu.pc.pc_o[2] ;
 wire \cu.pc.pc_o[3] ;
 wire \cu.pc.pc_o[4] ;
 wire \cu.pc.pc_o[5] ;
 wire \cu.pc.pc_o[6] ;
 wire \cu.pc.pc_o[7] ;
 wire \cu.pc.pc_o[8] ;
 wire \cu.pc.pc_o[9] ;
 wire \cu.reg_file.reg_a[0] ;
 wire \cu.reg_file.reg_a[1] ;
 wire \cu.reg_file.reg_a[2] ;
 wire \cu.reg_file.reg_a[3] ;
 wire \cu.reg_file.reg_a[4] ;
 wire \cu.reg_file.reg_a[5] ;
 wire \cu.reg_file.reg_a[6] ;
 wire \cu.reg_file.reg_a[7] ;
 wire \cu.reg_file.reg_b[0] ;
 wire \cu.reg_file.reg_b[1] ;
 wire \cu.reg_file.reg_b[2] ;
 wire \cu.reg_file.reg_b[3] ;
 wire \cu.reg_file.reg_b[4] ;
 wire \cu.reg_file.reg_b[5] ;
 wire \cu.reg_file.reg_b[6] ;
 wire \cu.reg_file.reg_b[7] ;
 wire \cu.reg_file.reg_c[0] ;
 wire \cu.reg_file.reg_c[1] ;
 wire \cu.reg_file.reg_c[2] ;
 wire \cu.reg_file.reg_c[3] ;
 wire \cu.reg_file.reg_c[4] ;
 wire \cu.reg_file.reg_c[5] ;
 wire \cu.reg_file.reg_c[6] ;
 wire \cu.reg_file.reg_c[7] ;
 wire \cu.reg_file.reg_d[0] ;
 wire \cu.reg_file.reg_d[1] ;
 wire \cu.reg_file.reg_d[2] ;
 wire \cu.reg_file.reg_d[3] ;
 wire \cu.reg_file.reg_d[4] ;
 wire \cu.reg_file.reg_d[5] ;
 wire \cu.reg_file.reg_d[6] ;
 wire \cu.reg_file.reg_d[7] ;
 wire \cu.reg_file.reg_e[0] ;
 wire \cu.reg_file.reg_e[1] ;
 wire \cu.reg_file.reg_e[2] ;
 wire \cu.reg_file.reg_e[3] ;
 wire \cu.reg_file.reg_e[4] ;
 wire \cu.reg_file.reg_e[5] ;
 wire \cu.reg_file.reg_e[6] ;
 wire \cu.reg_file.reg_e[7] ;
 wire \cu.reg_file.reg_h[0] ;
 wire \cu.reg_file.reg_h[1] ;
 wire \cu.reg_file.reg_h[2] ;
 wire \cu.reg_file.reg_h[3] ;
 wire \cu.reg_file.reg_h[4] ;
 wire \cu.reg_file.reg_h[5] ;
 wire \cu.reg_file.reg_h[6] ;
 wire \cu.reg_file.reg_h[7] ;
 wire \cu.reg_file.reg_l[0] ;
 wire \cu.reg_file.reg_l[1] ;
 wire \cu.reg_file.reg_l[2] ;
 wire \cu.reg_file.reg_l[3] ;
 wire \cu.reg_file.reg_l[4] ;
 wire \cu.reg_file.reg_l[5] ;
 wire \cu.reg_file.reg_l[6] ;
 wire \cu.reg_file.reg_l[7] ;
 wire \cu.reg_file.reg_mem[0] ;
 wire \cu.reg_file.reg_mem[10] ;
 wire \cu.reg_file.reg_mem[11] ;
 wire \cu.reg_file.reg_mem[12] ;
 wire \cu.reg_file.reg_mem[13] ;
 wire \cu.reg_file.reg_mem[14] ;
 wire \cu.reg_file.reg_mem[15] ;
 wire \cu.reg_file.reg_mem[1] ;
 wire \cu.reg_file.reg_mem[2] ;
 wire \cu.reg_file.reg_mem[3] ;
 wire \cu.reg_file.reg_mem[4] ;
 wire \cu.reg_file.reg_mem[5] ;
 wire \cu.reg_file.reg_mem[6] ;
 wire \cu.reg_file.reg_mem[7] ;
 wire \cu.reg_file.reg_mem[8] ;
 wire \cu.reg_file.reg_mem[9] ;
 wire \cu.reg_file.reg_sp[0] ;
 wire \cu.reg_file.reg_sp[10] ;
 wire \cu.reg_file.reg_sp[11] ;
 wire \cu.reg_file.reg_sp[12] ;
 wire \cu.reg_file.reg_sp[13] ;
 wire \cu.reg_file.reg_sp[14] ;
 wire \cu.reg_file.reg_sp[15] ;
 wire \cu.reg_file.reg_sp[1] ;
 wire \cu.reg_file.reg_sp[2] ;
 wire \cu.reg_file.reg_sp[3] ;
 wire \cu.reg_file.reg_sp[4] ;
 wire \cu.reg_file.reg_sp[5] ;
 wire \cu.reg_file.reg_sp[6] ;
 wire \cu.reg_file.reg_sp[7] ;
 wire \cu.reg_file.reg_sp[8] ;
 wire \cu.reg_file.reg_sp[9] ;
 wire \ih.gpio_interrupt_mask[0] ;
 wire \ih.gpio_interrupt_mask[1] ;
 wire \ih.gpio_interrupt_mask[2] ;
 wire \ih.gpio_interrupt_mask[3] ;
 wire \ih.gpio_interrupt_mask[4] ;
 wire \ih.gpio_interrupt_mask[5] ;
 wire \ih.gpio_interrupt_mask[6] ;
 wire \ih.gpio_interrupt_mask[7] ;
 wire \ih.ih.ih.prev_data[0] ;
 wire \ih.ih.ih.prev_data[10] ;
 wire \ih.ih.ih.prev_data[11] ;
 wire \ih.ih.ih.prev_data[12] ;
 wire \ih.ih.ih.prev_data[13] ;
 wire \ih.ih.ih.prev_data[14] ;
 wire \ih.ih.ih.prev_data[15] ;
 wire \ih.ih.ih.prev_data[1] ;
 wire \ih.ih.ih.prev_data[2] ;
 wire \ih.ih.ih.prev_data[3] ;
 wire \ih.ih.ih.prev_data[4] ;
 wire \ih.ih.ih.prev_data[5] ;
 wire \ih.ih.ih.prev_data[6] ;
 wire \ih.ih.ih.prev_data[7] ;
 wire \ih.ih.ih.prev_data[8] ;
 wire \ih.ih.ih.prev_data[9] ;
 wire \ih.ih.int_f.data_in ;
 wire \ih.ih.int_f.prev_data ;
 wire \ih.input_handler_enable ;
 wire \ih.interrupt_source[1] ;
 wire \ih.interrupt_source[2] ;
 wire \ih.interrupt_source[3] ;
 wire \ih.ip_ed.prev_data ;
 wire \ih.t.count[0] ;
 wire \ih.t.count[10] ;
 wire \ih.t.count[11] ;
 wire \ih.t.count[12] ;
 wire \ih.t.count[13] ;
 wire \ih.t.count[14] ;
 wire \ih.t.count[15] ;
 wire \ih.t.count[16] ;
 wire \ih.t.count[17] ;
 wire \ih.t.count[18] ;
 wire \ih.t.count[19] ;
 wire \ih.t.count[1] ;
 wire \ih.t.count[20] ;
 wire \ih.t.count[21] ;
 wire \ih.t.count[22] ;
 wire \ih.t.count[23] ;
 wire \ih.t.count[24] ;
 wire \ih.t.count[25] ;
 wire \ih.t.count[26] ;
 wire \ih.t.count[27] ;
 wire \ih.t.count[28] ;
 wire \ih.t.count[29] ;
 wire \ih.t.count[2] ;
 wire \ih.t.count[30] ;
 wire \ih.t.count[31] ;
 wire \ih.t.count[3] ;
 wire \ih.t.count[4] ;
 wire \ih.t.count[5] ;
 wire \ih.t.count[6] ;
 wire \ih.t.count[7] ;
 wire \ih.t.count[8] ;
 wire \ih.t.count[9] ;
 wire \ih.t.enable ;
 wire \ih.t.next_count[0] ;
 wire \ih.t.next_count[10] ;
 wire \ih.t.next_count[11] ;
 wire \ih.t.next_count[12] ;
 wire \ih.t.next_count[13] ;
 wire \ih.t.next_count[14] ;
 wire \ih.t.next_count[15] ;
 wire \ih.t.next_count[16] ;
 wire \ih.t.next_count[17] ;
 wire \ih.t.next_count[18] ;
 wire \ih.t.next_count[19] ;
 wire \ih.t.next_count[1] ;
 wire \ih.t.next_count[20] ;
 wire \ih.t.next_count[21] ;
 wire \ih.t.next_count[22] ;
 wire \ih.t.next_count[23] ;
 wire \ih.t.next_count[24] ;
 wire \ih.t.next_count[25] ;
 wire \ih.t.next_count[26] ;
 wire \ih.t.next_count[27] ;
 wire \ih.t.next_count[28] ;
 wire \ih.t.next_count[29] ;
 wire \ih.t.next_count[2] ;
 wire \ih.t.next_count[30] ;
 wire \ih.t.next_count[31] ;
 wire \ih.t.next_count[3] ;
 wire \ih.t.next_count[4] ;
 wire \ih.t.next_count[5] ;
 wire \ih.t.next_count[6] ;
 wire \ih.t.next_count[7] ;
 wire \ih.t.next_count[8] ;
 wire \ih.t.next_count[9] ;
 wire \ih.t.timer_max[0] ;
 wire \ih.t.timer_max[10] ;
 wire \ih.t.timer_max[11] ;
 wire \ih.t.timer_max[12] ;
 wire \ih.t.timer_max[13] ;
 wire \ih.t.timer_max[14] ;
 wire \ih.t.timer_max[15] ;
 wire \ih.t.timer_max[16] ;
 wire \ih.t.timer_max[17] ;
 wire \ih.t.timer_max[18] ;
 wire \ih.t.timer_max[19] ;
 wire \ih.t.timer_max[1] ;
 wire \ih.t.timer_max[20] ;
 wire \ih.t.timer_max[21] ;
 wire \ih.t.timer_max[22] ;
 wire \ih.t.timer_max[23] ;
 wire \ih.t.timer_max[24] ;
 wire \ih.t.timer_max[25] ;
 wire \ih.t.timer_max[26] ;
 wire \ih.t.timer_max[27] ;
 wire \ih.t.timer_max[28] ;
 wire \ih.t.timer_max[29] ;
 wire \ih.t.timer_max[2] ;
 wire \ih.t.timer_max[30] ;
 wire \ih.t.timer_max[31] ;
 wire \ih.t.timer_max[3] ;
 wire \ih.t.timer_max[4] ;
 wire \ih.t.timer_max[5] ;
 wire \ih.t.timer_max[6] ;
 wire \ih.t.timer_max[7] ;
 wire \ih.t.timer_max[8] ;
 wire \ih.t.timer_max[9] ;
 wire \mc.cc.count[0] ;
 wire \mc.cc.count[1] ;
 wire \mc.cc.count[2] ;
 wire \mc.cc.count[3] ;
 wire \mc.cc.enable ;
 wire \mc.cc.enable_edge_detector.prev_data ;
 wire \mc.cl.cmp_o ;
 wire \mc.cl.next_data[0] ;
 wire \mc.cl.next_data[10] ;
 wire \mc.cl.next_data[11] ;
 wire \mc.cl.next_data[12] ;
 wire \mc.cl.next_data[13] ;
 wire \mc.cl.next_data[14] ;
 wire \mc.cl.next_data[15] ;
 wire \mc.cl.next_data[1] ;
 wire \mc.cl.next_data[2] ;
 wire \mc.cl.next_data[3] ;
 wire \mc.cl.next_data[4] ;
 wire \mc.cl.next_data[5] ;
 wire \mc.cl.next_data[6] ;
 wire \mc.cl.next_data[7] ;
 wire \mc.cl.next_data[8] ;
 wire \mc.cl.next_data[9] ;
 wire \mc.count ;
 wire \mc.rw.cmp_check ;
 wire \mc.rw.next_state[0] ;
 wire \mc.rw.next_state[1] ;
 wire \mc.rw.next_state[2] ;
 wire \mc.rw.state[0] ;
 wire \mc.rw.state[1] ;
 wire \mc.rw.state[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0306_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\cu.pc.pc_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\ih.t.timer_max[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\ih.t.timer_max[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(keypad_input[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(memory_data_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(programmable_gpio_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(programmable_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__B (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__B (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__B (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__B (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__B (.DIODE(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A (.DIODE(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A (.DIODE(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__B1 (.DIODE(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__B1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B1 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__A2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A_N (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A_N (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__B_N (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__B (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A1 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__B (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A1 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__B1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__B1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__C1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__C (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__C1 (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B1_N (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A1_N (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__B1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__D1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__B (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A1 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__B (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__B (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__B1 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A1 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__B1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__B1 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__C1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A1 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B2 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__B1 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__B1 (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B1 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B1 (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__B_N (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B1 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A_N (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__B1_N (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A_N (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__D (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__C (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A_N (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__B2 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__C_N (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A1 (.DIODE(\cu.reg_file.reg_mem[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A1 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A1 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__B2 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B1_N (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A1 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A2 (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A2 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__C1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__B1 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__C1 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B2 (.DIODE(\cu.reg_file.reg_mem[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A (.DIODE(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A1 (.DIODE(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__B2 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B2 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A1 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__C1 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__C1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__C1 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__B (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A1 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__B2 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A1 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A1 (.DIODE(\cu.reg_file.reg_mem[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B_N (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A1 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B2 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B2 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B2 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B2 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B2 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A1 (.DIODE(\cu.reg_file.reg_mem[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B2 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(\cu.reg_file.reg_mem[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__B2 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A1 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B2 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B2 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B2 (.DIODE(\cu.reg_file.reg_mem[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B2 (.DIODE(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A1 (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A2 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__B (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B2 (.DIODE(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A1 (.DIODE(\cu.reg_file.reg_mem[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B2 (.DIODE(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B2 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__C_N (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B2 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B2 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(\cu.reg_file.reg_mem[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__S (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B2 (.DIODE(\cu.reg_file.reg_mem[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A1 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__C_N (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B2 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B2 (.DIODE(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A0 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__S (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B2 (.DIODE(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B2 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B2 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__B2 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A1 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A1 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B2 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__D1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B2 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B2 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__B2 (.DIODE(\cu.reg_file.reg_mem[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B2 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B2 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__B (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B2 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__D1 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A1 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B2 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A1 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A1_N (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__B (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B2 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B2 (.DIODE(\cu.reg_file.reg_mem[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A1 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A1 (.DIODE(\cu.reg_file.reg_mem[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A_N (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B2 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A1 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B2 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B2 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A1 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B2 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A1 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A1 (.DIODE(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B2 (.DIODE(\cu.reg_file.reg_mem[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A1 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B2 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(\cu.reg_file.reg_mem[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B2 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A1 (.DIODE(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B2 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__B2 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A1 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B2 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A1 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B2 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A1 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A1 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B2 (.DIODE(\cu.reg_file.reg_mem[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A1 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(\cu.reg_file.reg_mem[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B2 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B2 (.DIODE(\cu.reg_file.reg_mem[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(\cu.reg_file.reg_mem[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B2 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__B1 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__C1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__C1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B2 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__D (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__C (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A1 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B1 (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__D (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B1 (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B (.DIODE(_0529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__C1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A2 (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A2 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A1_N (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A2 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B2 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A1_N (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A2_N (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A2_N (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__C1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__C1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A1_N (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__B1 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__B1 (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A2 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A2 (.DIODE(_1185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B2 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(_1185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__B2 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A2 (.DIODE(_1185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__B2 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B2 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__C1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__B1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__C (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A3 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A1 (.DIODE(_1032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__C (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__C (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__B (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__C (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__D (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A0 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A0 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A0 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A2 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A2 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__C (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__C1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__C1 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A1 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B2 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A (.DIODE(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B2 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__C1 (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A1 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A3 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__C1 (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A_N (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__C (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B_N (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__D_N (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A2 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__B2 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__B2 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__B1_N (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__C (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B2 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A1 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B2 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A1 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B2 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A1 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__C1 (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__B2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A1 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B2 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__B2 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__B2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__B1 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__C1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__B1 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__B1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__B2 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B2 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A1 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__B2 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B2 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B2 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__B (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A_N (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__B (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A1 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B2 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__B2 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B2 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B2 (.DIODE(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__B2 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B2 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__C1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A1 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__B2 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__C1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B2 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A2 (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A2 (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B2 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__B2 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__C1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A1 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B2 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__B2 (.DIODE(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B2 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__B2 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A1 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__B2 (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A1 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A1 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B2 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A1 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__B2 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B2 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B2 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__C1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__B2 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A1 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__B2 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A2 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B2 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B2 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__C1 (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A1 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B2 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B2 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A1 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A1 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B2 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A1 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__B2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B2 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__C1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__B2 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__B2 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B2 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A1 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B2 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A1 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__B2 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__B2 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__B2 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B2 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A1 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B2 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B2 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__C1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B2 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__C1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B2 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A1 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B2 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A1 (.DIODE(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__B2 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__C1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B2 (.DIODE(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__C1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B2 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B2 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A1 (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__B (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A1 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__B1 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__B2 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A1 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B2 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__B1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__B2 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__B2 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__B2 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__B (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__B (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__B (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A2 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B1 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B2 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A1 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B2 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A1 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__B2 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A1 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B2 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A1 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B2 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__B2 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__B (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A3 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A2 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A2 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A2 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A2 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A2 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A2 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A2 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__C (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__D (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__D (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__C1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A (.DIODE(\mc.cl.cmp_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__C (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A (.DIODE(\mc.cl.cmp_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__C (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A0 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A2 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__C (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A1 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A2 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A3 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A0 (.DIODE(\cu.alu_f[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A1 (.DIODE(\alu.Cin ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B1 (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__B1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A3 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B1 (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(\cu.id.is_halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A2 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A3 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__C (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__B1 (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A2 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1 (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A (.DIODE(_1185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A0 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__C1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A0 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A0 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A0 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__C (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__B1 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A2 (.DIODE(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A0 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A0 (.DIODE(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A0 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A0 (.DIODE(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A0 (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A0 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A1 (.DIODE(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B1 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A0 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A0 (.DIODE(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A0 (.DIODE(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A0 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A0 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B1 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A (.DIODE(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__B1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A0 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A0 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A0 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A1 (.DIODE(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A2 (.DIODE(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A0 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__B1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A0 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A0 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A0 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A0 (.DIODE(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A0 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A0 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B1_N (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A0 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A0 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A1 (.DIODE(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A0 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A0 (.DIODE(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A0 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A0 (.DIODE(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A0 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A0 (.DIODE(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A0 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A0 (.DIODE(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A0 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A0 (.DIODE(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A0 (.DIODE(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A0 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__S (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A0 (.DIODE(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__S (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A0 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A1 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A0 (.DIODE(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A0 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A0 (.DIODE(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A0 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A0 (.DIODE(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A0 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A0 (.DIODE(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A0 (.DIODE(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A0 (.DIODE(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A0 (.DIODE(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A0 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A0 (.DIODE(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B1 (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A0 (.DIODE(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A0 (.DIODE(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A1 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A0 (.DIODE(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A0 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B1 (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A0 (.DIODE(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A0 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A0 (.DIODE(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A0 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A0 (.DIODE(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A0 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A0 (.DIODE(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A0 (.DIODE(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A0 (.DIODE(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A0 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A0 (.DIODE(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A0 (.DIODE(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A0 (.DIODE(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A0 (.DIODE(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A0 (.DIODE(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A0 (.DIODE(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A0 (.DIODE(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B1_N (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A0 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1 (.DIODE(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A0 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A0 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A1 (.DIODE(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A0 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A0 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A0 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A0 (.DIODE(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A0 (.DIODE(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A1 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__S (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__C_N (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__C1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__C (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A0 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__S (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A0 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__S (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A0 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__S (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A0 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__S (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A0 (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__S (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A0 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A0 (.DIODE(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_2162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A0 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__S (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A0 (.DIODE(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__S (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__S (.DIODE(_2167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__S (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__S (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__S (.DIODE(_2203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__S (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__S (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A0 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__S (.DIODE(_2234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A0 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A0 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A0 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A0 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__S (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__C (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__S0 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__S1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A2 (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(\mc.cl.cmp_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B2 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(\ih.t.enable ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C1 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__C1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__D1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__C (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__S0 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__S1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B2 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A0 (.DIODE(\cu.reg_file.reg_mem[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B2 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__C1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__C (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A0 (.DIODE(\cu.reg_file.reg_mem[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__C1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A0 (.DIODE(\cu.reg_file.reg_mem[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__C1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A0 (.DIODE(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__C1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A0 (.DIODE(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(_2425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__C1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A0 (.DIODE(\cu.reg_file.reg_mem[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__S (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B1 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__C1 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A0 (.DIODE(\cu.reg_file.reg_mem[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__B (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B1 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A1 (.DIODE(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B2 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A_N (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__C1 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B2 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__C (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B1 (.DIODE(\cu.reg_file.reg_mem[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B1 (.DIODE(\cu.reg_file.reg_mem[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B2 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B1 (.DIODE(\cu.reg_file.reg_mem[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B2 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B1 (.DIODE(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B1 (.DIODE(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__B2 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B1 (.DIODE(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B2 (.DIODE(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B1 (.DIODE(\cu.reg_file.reg_mem[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__B2 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A2_N (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B1 (.DIODE(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A3 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__B (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B1 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B1 (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A0 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A0 (.DIODE(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A0 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A0 (.DIODE(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A0 (.DIODE(_1159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A0 (.DIODE(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A0 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A0 (.DIODE(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A0 (.DIODE(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A0 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A0 (.DIODE(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A0 (.DIODE(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A0 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A0 (.DIODE(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__S (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A2 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A0 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__S (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A0 (.DIODE(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__S (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A0 (.DIODE(_1212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__S (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__S (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__B (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A0 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__S (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__S (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A0 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__S (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__S (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A0 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__S (.DIODE(_2119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A0 (.DIODE(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__S (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A1 (.DIODE(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A1 (.DIODE(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A0 (.DIODE(_2162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A2 (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A0 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A0 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A0 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A0 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A0 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A0 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A0 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__S (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A2 (.DIODE(_2202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A1 (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A1 (.DIODE(_1186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A1 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A0 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A0 (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(_2425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A0 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A1 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A0 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A0 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A0 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A0 (.DIODE(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A0 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(_2425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A0 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A0 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A0 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A0 (.DIODE(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A0 (.DIODE(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A0 (.DIODE(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A0 (.DIODE(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A0 (.DIODE(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(_2425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A0 (.DIODE(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A1 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A0 (.DIODE(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A0 (.DIODE(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__RESET_B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__SET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__D (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__RESET_B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__RESET_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__RESET_B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__RESET_B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1_A (.DIODE(\cu.id.is_halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire143_A (.DIODE(net144));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2957_ (.A(\mc.rw.state[1] ),
    .Y(_2697_));
 sky130_fd_sc_hd__and3_1 _2958_ (.A(\mc.rw.state[2] ),
    .B(_2697_),
    .C(\mc.rw.state[0] ),
    .X(_2698_));
 sky130_fd_sc_hd__clkbuf_8 _2959_ (.A(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__inv_2 _2960_ (.A(\mc.rw.state[2] ),
    .Y(_2700_));
 sky130_fd_sc_hd__nor2_2 _2961_ (.A(_2697_),
    .B(\mc.rw.state[0] ),
    .Y(_2701_));
 sky130_fd_sc_hd__and3b_1 _2962_ (.A_N(\mc.rw.state[0] ),
    .B(\mc.rw.state[2] ),
    .C(_2697_),
    .X(_2702_));
 sky130_fd_sc_hd__clkbuf_2 _2963_ (.A(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a21o_4 _2964_ (.A1(_2700_),
    .A2(_2701_),
    .B1(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__or2_1 _2965_ (.A(_2699_),
    .B(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_2705_),
    .X(net59));
 sky130_fd_sc_hd__or3_2 _2967_ (.A(_2700_),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .X(_2706_));
 sky130_fd_sc_hd__and2_1 _2968_ (.A(_2697_),
    .B(\mc.rw.state[0] ),
    .X(_2707_));
 sky130_fd_sc_hd__nor2_1 _2969_ (.A(_2707_),
    .B(_2701_),
    .Y(_2708_));
 sky130_fd_sc_hd__and3_2 _2970_ (.A(_2700_),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .X(_2709_));
 sky130_fd_sc_hd__inv_2 _2971_ (.A(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__and3_2 _2972_ (.A(_2706_),
    .B(_2708_),
    .C(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__inv_2 _2973_ (.A(_2711_),
    .Y(\mc.cc.enable ));
 sky130_fd_sc_hd__inv_2 _2974_ (.A(net9),
    .Y(_2712_));
 sky130_fd_sc_hd__inv_2 _2975_ (.A(net4),
    .Y(_2713_));
 sky130_fd_sc_hd__inv_2 _2976_ (.A(net10),
    .Y(_2714_));
 sky130_fd_sc_hd__inv_2 _2977_ (.A(net11),
    .Y(_2715_));
 sky130_fd_sc_hd__o22a_1 _2978_ (.A1(_2714_),
    .A2(\ih.ih.ih.prev_data[2] ),
    .B1(_2715_),
    .B2(\ih.ih.ih.prev_data[3] ),
    .X(_2716_));
 sky130_fd_sc_hd__o221a_1 _2979_ (.A1(_2712_),
    .A2(\ih.ih.ih.prev_data[1] ),
    .B1(_2713_),
    .B2(net225),
    .C1(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__inv_2 _2980_ (.A(net14),
    .Y(_2718_));
 sky130_fd_sc_hd__inv_2 _2981_ (.A(net5),
    .Y(_2719_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(net12),
    .Y(_2720_));
 sky130_fd_sc_hd__inv_2 _2983_ (.A(net6),
    .Y(_2721_));
 sky130_fd_sc_hd__o22a_1 _2984_ (.A1(_2720_),
    .A2(\ih.ih.ih.prev_data[4] ),
    .B1(_2721_),
    .B2(\ih.ih.ih.prev_data[13] ),
    .X(_2722_));
 sky130_fd_sc_hd__o221a_1 _2985_ (.A1(_2718_),
    .A2(\ih.ih.ih.prev_data[6] ),
    .B1(_2719_),
    .B2(\ih.ih.ih.prev_data[12] ),
    .C1(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__inv_2 _2986_ (.A(net17),
    .Y(_2724_));
 sky130_fd_sc_hd__inv_2 _2987_ (.A(net7),
    .Y(_2725_));
 sky130_fd_sc_hd__inv_2 _2988_ (.A(net13),
    .Y(_2726_));
 sky130_fd_sc_hd__inv_2 _2989_ (.A(net3),
    .Y(_2727_));
 sky130_fd_sc_hd__o22a_1 _2990_ (.A1(_2726_),
    .A2(\ih.ih.ih.prev_data[5] ),
    .B1(_2727_),
    .B2(\ih.ih.ih.prev_data[10] ),
    .X(_2728_));
 sky130_fd_sc_hd__o221a_1 _2991_ (.A1(_2724_),
    .A2(\ih.ih.ih.prev_data[9] ),
    .B1(_2725_),
    .B2(\ih.ih.ih.prev_data[14] ),
    .C1(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__inv_2 _2992_ (.A(net2),
    .Y(_2730_));
 sky130_fd_sc_hd__inv_2 _2993_ (.A(net8),
    .Y(_2731_));
 sky130_fd_sc_hd__inv_2 _2994_ (.A(net15),
    .Y(_2732_));
 sky130_fd_sc_hd__inv_2 _2995_ (.A(net16),
    .Y(_2733_));
 sky130_fd_sc_hd__o22a_1 _2996_ (.A1(_2732_),
    .A2(\ih.ih.ih.prev_data[7] ),
    .B1(_2733_),
    .B2(\ih.ih.ih.prev_data[8] ),
    .X(_2734_));
 sky130_fd_sc_hd__o221a_1 _2997_ (.A1(_2730_),
    .A2(\ih.ih.ih.prev_data[0] ),
    .B1(_2731_),
    .B2(\ih.ih.ih.prev_data[15] ),
    .C1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__and3_1 _2998_ (.A(_2723_),
    .B(_2729_),
    .C(_2735_),
    .X(_2736_));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(net226),
    .B(_2736_),
    .Y(\ih.ih.int_f.data_in ));
 sky130_fd_sc_hd__or3_1 _3000_ (.A(\ih.t.timer_max[0] ),
    .B(\ih.t.timer_max[1] ),
    .C(\ih.t.timer_max[2] ),
    .X(_2737_));
 sky130_fd_sc_hd__or2_1 _3001_ (.A(\ih.t.timer_max[3] ),
    .B(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__or2_1 _3002_ (.A(\ih.t.timer_max[4] ),
    .B(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3003_ (.A(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__or3_2 _3004_ (.A(\ih.t.timer_max[5] ),
    .B(\ih.t.timer_max[6] ),
    .C(_2740_),
    .X(_2741_));
 sky130_fd_sc_hd__or3_1 _3005_ (.A(\ih.t.timer_max[7] ),
    .B(\ih.t.timer_max[8] ),
    .C(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__or2_2 _3006_ (.A(\ih.t.timer_max[9] ),
    .B(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__or3_1 _3007_ (.A(\ih.t.timer_max[10] ),
    .B(\ih.t.timer_max[11] ),
    .C(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__or2_2 _3008_ (.A(\ih.t.timer_max[12] ),
    .B(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__or3_1 _3009_ (.A(\ih.t.timer_max[13] ),
    .B(\ih.t.timer_max[14] ),
    .C(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__or2_2 _3010_ (.A(\ih.t.timer_max[15] ),
    .B(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__or3_1 _3011_ (.A(\ih.t.timer_max[16] ),
    .B(\ih.t.timer_max[17] ),
    .C(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__or2_2 _3012_ (.A(\ih.t.timer_max[18] ),
    .B(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__or3_1 _3013_ (.A(\ih.t.timer_max[19] ),
    .B(\ih.t.timer_max[20] ),
    .C(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__or2_2 _3014_ (.A(\ih.t.timer_max[21] ),
    .B(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__or3_1 _3015_ (.A(\ih.t.timer_max[22] ),
    .B(\ih.t.timer_max[23] ),
    .C(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__or2_2 _3016_ (.A(\ih.t.timer_max[24] ),
    .B(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__or3_1 _3017_ (.A(\ih.t.timer_max[25] ),
    .B(\ih.t.timer_max[26] ),
    .C(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__or2_2 _3018_ (.A(\ih.t.timer_max[27] ),
    .B(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__or3_1 _3019_ (.A(\ih.t.timer_max[28] ),
    .B(\ih.t.timer_max[29] ),
    .C(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__nor2_1 _3020_ (.A(\ih.t.timer_max[30] ),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__xnor2_1 _3021_ (.A(\ih.t.count[31] ),
    .B(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__xnor2_1 _3022_ (.A(\ih.t.timer_max[31] ),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__o21ai_1 _3023_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2755_),
    .B1(\ih.t.timer_max[29] ),
    .Y(_2760_));
 sky130_fd_sc_hd__and3_1 _3024_ (.A(\ih.t.count[29] ),
    .B(_2756_),
    .C(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__a21oi_1 _3025_ (.A1(_2756_),
    .A2(_2760_),
    .B1(\ih.t.count[29] ),
    .Y(_2762_));
 sky130_fd_sc_hd__xor2_1 _3026_ (.A(\ih.t.timer_max[28] ),
    .B(_2755_),
    .X(_2763_));
 sky130_fd_sc_hd__xnor2_1 _3027_ (.A(\ih.t.count[28] ),
    .B(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand2_1 _3028_ (.A(\ih.t.timer_max[27] ),
    .B(_2754_),
    .Y(_2765_));
 sky130_fd_sc_hd__a21oi_1 _3029_ (.A1(_2755_),
    .A2(_2765_),
    .B1(\ih.t.count[27] ),
    .Y(_2766_));
 sky130_fd_sc_hd__and3_1 _3030_ (.A(\ih.t.count[27] ),
    .B(_2755_),
    .C(_2765_),
    .X(_2767_));
 sky130_fd_sc_hd__o21ai_1 _3031_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2753_),
    .B1(\ih.t.timer_max[26] ),
    .Y(_2768_));
 sky130_fd_sc_hd__and3_1 _3032_ (.A(\ih.t.count[26] ),
    .B(_2754_),
    .C(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__a21oi_1 _3033_ (.A1(_2754_),
    .A2(_2768_),
    .B1(\ih.t.count[26] ),
    .Y(_2770_));
 sky130_fd_sc_hd__xor2_1 _3034_ (.A(\ih.t.timer_max[25] ),
    .B(_2753_),
    .X(_2771_));
 sky130_fd_sc_hd__xnor2_1 _3035_ (.A(\ih.t.count[25] ),
    .B(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__nand2_1 _3036_ (.A(\ih.t.timer_max[24] ),
    .B(_2752_),
    .Y(_2773_));
 sky130_fd_sc_hd__and3_1 _3037_ (.A(\ih.t.count[24] ),
    .B(_2753_),
    .C(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__a21oi_1 _3038_ (.A1(_2753_),
    .A2(_2773_),
    .B1(\ih.t.count[24] ),
    .Y(_2775_));
 sky130_fd_sc_hd__o21ai_1 _3039_ (.A1(\ih.t.timer_max[22] ),
    .A2(_2751_),
    .B1(\ih.t.timer_max[23] ),
    .Y(_2776_));
 sky130_fd_sc_hd__and3_1 _3040_ (.A(\ih.t.count[23] ),
    .B(_2752_),
    .C(_2776_),
    .X(_2777_));
 sky130_fd_sc_hd__a21oi_1 _3041_ (.A1(_2752_),
    .A2(_2776_),
    .B1(\ih.t.count[23] ),
    .Y(_2778_));
 sky130_fd_sc_hd__xor2_1 _3042_ (.A(\ih.t.timer_max[22] ),
    .B(_2751_),
    .X(_2779_));
 sky130_fd_sc_hd__xnor2_1 _3043_ (.A(\ih.t.count[22] ),
    .B(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(\ih.t.timer_max[21] ),
    .B(_2750_),
    .Y(_2781_));
 sky130_fd_sc_hd__and3_1 _3045_ (.A(\ih.t.count[21] ),
    .B(_2751_),
    .C(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__a21oi_1 _3046_ (.A1(_2751_),
    .A2(_2781_),
    .B1(\ih.t.count[21] ),
    .Y(_2783_));
 sky130_fd_sc_hd__o21ai_1 _3047_ (.A1(\ih.t.timer_max[19] ),
    .A2(_2749_),
    .B1(\ih.t.timer_max[20] ),
    .Y(_2784_));
 sky130_fd_sc_hd__a21oi_1 _3048_ (.A1(_2750_),
    .A2(_2784_),
    .B1(\ih.t.count[20] ),
    .Y(_2785_));
 sky130_fd_sc_hd__and3_1 _3049_ (.A(\ih.t.count[20] ),
    .B(_2750_),
    .C(_2784_),
    .X(_2786_));
 sky130_fd_sc_hd__xor2_1 _3050_ (.A(\ih.t.timer_max[19] ),
    .B(_2749_),
    .X(_2787_));
 sky130_fd_sc_hd__xnor2_1 _3051_ (.A(\ih.t.count[19] ),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nand2_1 _3052_ (.A(\ih.t.timer_max[18] ),
    .B(_2748_),
    .Y(_2789_));
 sky130_fd_sc_hd__a21oi_1 _3053_ (.A1(_2749_),
    .A2(_2789_),
    .B1(\ih.t.count[18] ),
    .Y(_2790_));
 sky130_fd_sc_hd__and3_1 _3054_ (.A(\ih.t.count[18] ),
    .B(_2749_),
    .C(_2789_),
    .X(_2791_));
 sky130_fd_sc_hd__o21ai_1 _3055_ (.A1(\ih.t.timer_max[16] ),
    .A2(_2747_),
    .B1(\ih.t.timer_max[17] ),
    .Y(_2792_));
 sky130_fd_sc_hd__a21oi_1 _3056_ (.A1(_2748_),
    .A2(_2792_),
    .B1(\ih.t.count[17] ),
    .Y(_2793_));
 sky130_fd_sc_hd__and3_1 _3057_ (.A(\ih.t.count[17] ),
    .B(_2748_),
    .C(_2792_),
    .X(_2794_));
 sky130_fd_sc_hd__xor2_1 _3058_ (.A(\ih.t.timer_max[16] ),
    .B(_2747_),
    .X(_2795_));
 sky130_fd_sc_hd__xnor2_1 _3059_ (.A(\ih.t.count[16] ),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand2_1 _3060_ (.A(\ih.t.timer_max[15] ),
    .B(_2746_),
    .Y(_2797_));
 sky130_fd_sc_hd__a21oi_1 _3061_ (.A1(_2747_),
    .A2(_2797_),
    .B1(\ih.t.count[15] ),
    .Y(_2798_));
 sky130_fd_sc_hd__and3_1 _3062_ (.A(\ih.t.count[15] ),
    .B(_2747_),
    .C(_2797_),
    .X(_2799_));
 sky130_fd_sc_hd__o21ai_1 _3063_ (.A1(\ih.t.timer_max[13] ),
    .A2(_2745_),
    .B1(\ih.t.timer_max[14] ),
    .Y(_2800_));
 sky130_fd_sc_hd__and3_1 _3064_ (.A(\ih.t.count[14] ),
    .B(_2746_),
    .C(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__a21oi_1 _3065_ (.A1(_2746_),
    .A2(_2800_),
    .B1(\ih.t.count[14] ),
    .Y(_2802_));
 sky130_fd_sc_hd__xor2_1 _3066_ (.A(\ih.t.timer_max[13] ),
    .B(_2745_),
    .X(_2803_));
 sky130_fd_sc_hd__xnor2_1 _3067_ (.A(\ih.t.count[13] ),
    .B(_2803_),
    .Y(_2804_));
 sky130_fd_sc_hd__nand2_1 _3068_ (.A(\ih.t.timer_max[12] ),
    .B(_2744_),
    .Y(_2805_));
 sky130_fd_sc_hd__and3_1 _3069_ (.A(\ih.t.count[12] ),
    .B(_2745_),
    .C(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__a21oi_1 _3070_ (.A1(_2745_),
    .A2(_2805_),
    .B1(\ih.t.count[12] ),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_1 _3071_ (.A1(\ih.t.timer_max[10] ),
    .A2(_2743_),
    .B1(\ih.t.timer_max[11] ),
    .Y(_2808_));
 sky130_fd_sc_hd__a21oi_1 _3072_ (.A1(_2744_),
    .A2(_2808_),
    .B1(\ih.t.count[11] ),
    .Y(_2809_));
 sky130_fd_sc_hd__and3_1 _3073_ (.A(\ih.t.count[11] ),
    .B(_2744_),
    .C(_2808_),
    .X(_2810_));
 sky130_fd_sc_hd__xor2_1 _3074_ (.A(\ih.t.timer_max[10] ),
    .B(_2743_),
    .X(_2811_));
 sky130_fd_sc_hd__xnor2_1 _3075_ (.A(\ih.t.count[10] ),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(\ih.t.timer_max[9] ),
    .B(_2742_),
    .Y(_2813_));
 sky130_fd_sc_hd__and3_1 _3077_ (.A(\ih.t.count[9] ),
    .B(_2743_),
    .C(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__a21oi_1 _3078_ (.A1(_2743_),
    .A2(_2813_),
    .B1(\ih.t.count[9] ),
    .Y(_2815_));
 sky130_fd_sc_hd__o21ai_1 _3079_ (.A1(\ih.t.timer_max[7] ),
    .A2(_2741_),
    .B1(\ih.t.timer_max[8] ),
    .Y(_2816_));
 sky130_fd_sc_hd__and3_1 _3080_ (.A(\ih.t.count[8] ),
    .B(_2742_),
    .C(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__a21oi_1 _3081_ (.A1(_2742_),
    .A2(_2816_),
    .B1(\ih.t.count[8] ),
    .Y(_2818_));
 sky130_fd_sc_hd__xor2_1 _3082_ (.A(\ih.t.timer_max[7] ),
    .B(_2741_),
    .X(_2819_));
 sky130_fd_sc_hd__xnor2_1 _3083_ (.A(\ih.t.count[7] ),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__o21ai_1 _3084_ (.A1(\ih.t.timer_max[5] ),
    .A2(_2740_),
    .B1(\ih.t.timer_max[6] ),
    .Y(_2821_));
 sky130_fd_sc_hd__and3_1 _3085_ (.A(\ih.t.count[6] ),
    .B(_2741_),
    .C(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__a21oi_1 _3086_ (.A1(_2741_),
    .A2(_2821_),
    .B1(\ih.t.count[6] ),
    .Y(_2823_));
 sky130_fd_sc_hd__xor2_1 _3087_ (.A(\ih.t.timer_max[5] ),
    .B(_2740_),
    .X(_2824_));
 sky130_fd_sc_hd__xnor2_1 _3088_ (.A(\ih.t.count[5] ),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _3089_ (.A(\ih.t.timer_max[4] ),
    .B(_2738_),
    .Y(_2826_));
 sky130_fd_sc_hd__and2_1 _3090_ (.A(\ih.t.timer_max[0] ),
    .B(\ih.t.count[0] ),
    .X(_2827_));
 sky130_fd_sc_hd__o21ai_1 _3091_ (.A1(\ih.t.timer_max[0] ),
    .A2(\ih.t.timer_max[1] ),
    .B1(\ih.t.timer_max[2] ),
    .Y(_2828_));
 sky130_fd_sc_hd__and3_1 _3092_ (.A(\ih.t.count[2] ),
    .B(_2737_),
    .C(_2828_),
    .X(_2829_));
 sky130_fd_sc_hd__a21oi_1 _3093_ (.A1(_2737_),
    .A2(_2828_),
    .B1(\ih.t.count[2] ),
    .Y(_2830_));
 sky130_fd_sc_hd__xor2_1 _3094_ (.A(\ih.t.timer_max[1] ),
    .B(\ih.t.count[1] ),
    .X(_2831_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(\ih.t.timer_max[0] ),
    .A1(\ih.t.count[0] ),
    .S(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__or4b_1 _3096_ (.A(_2827_),
    .B(_2829_),
    .C(_2830_),
    .D_N(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__a31o_1 _3097_ (.A1(\ih.t.count[4] ),
    .A2(_2740_),
    .A3(_2826_),
    .B1(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__a21oi_1 _3098_ (.A1(_2740_),
    .A2(_2826_),
    .B1(\ih.t.count[4] ),
    .Y(_2835_));
 sky130_fd_sc_hd__nand2_1 _3099_ (.A(\ih.t.timer_max[3] ),
    .B(_2737_),
    .Y(_2836_));
 sky130_fd_sc_hd__nand2_1 _3100_ (.A(_2738_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__xor2_1 _3101_ (.A(\ih.t.count[3] ),
    .B(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__or4_1 _3102_ (.A(_2825_),
    .B(_2834_),
    .C(_2835_),
    .D(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__or4_1 _3103_ (.A(_2820_),
    .B(_2822_),
    .C(_2823_),
    .D(_2839_),
    .X(_2840_));
 sky130_fd_sc_hd__or3_1 _3104_ (.A(_2817_),
    .B(_2818_),
    .C(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__or4_1 _3105_ (.A(_2812_),
    .B(_2814_),
    .C(_2815_),
    .D(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__or3_1 _3106_ (.A(_2809_),
    .B(_2810_),
    .C(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__or4_1 _3107_ (.A(_2804_),
    .B(_2806_),
    .C(_2807_),
    .D(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__or3_1 _3108_ (.A(_2801_),
    .B(_2802_),
    .C(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__or4_1 _3109_ (.A(_2796_),
    .B(_2798_),
    .C(_2799_),
    .D(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__or3_1 _3110_ (.A(_2793_),
    .B(_2794_),
    .C(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__or4_1 _3111_ (.A(_2788_),
    .B(_2790_),
    .C(_2791_),
    .D(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__or3_1 _3112_ (.A(_2785_),
    .B(_2786_),
    .C(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__or4_1 _3113_ (.A(_2780_),
    .B(_2782_),
    .C(_2783_),
    .D(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__or3_1 _3114_ (.A(_2777_),
    .B(_2778_),
    .C(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__or4_1 _3115_ (.A(_2772_),
    .B(_2774_),
    .C(_2775_),
    .D(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__or3_1 _3116_ (.A(_2769_),
    .B(_2770_),
    .C(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__or4_1 _3117_ (.A(_2764_),
    .B(_2766_),
    .C(_2767_),
    .D(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__or3_1 _3118_ (.A(_2761_),
    .B(_2762_),
    .C(_2854_),
    .X(_2855_));
 sky130_fd_sc_hd__and2_1 _3119_ (.A(\ih.t.timer_max[30] ),
    .B(_2756_),
    .X(_2856_));
 sky130_fd_sc_hd__nor2_1 _3120_ (.A(_2757_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__nor2_1 _3121_ (.A(\ih.t.count[30] ),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand2_1 _3122_ (.A(\ih.t.count[30] ),
    .B(_2857_),
    .Y(_2859_));
 sky130_fd_sc_hd__or4b_4 _3123_ (.A(_2759_),
    .B(_2855_),
    .C(_2858_),
    .D_N(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__inv_2 _3124_ (.A(net69),
    .Y(_2861_));
 sky130_fd_sc_hd__and3b_1 _3125_ (.A_N(net68),
    .B(net27),
    .C(\ih.gpio_interrupt_mask[0] ),
    .X(_2862_));
 sky130_fd_sc_hd__a31o_1 _3126_ (.A1(_2861_),
    .A2(net28),
    .A3(\ih.gpio_interrupt_mask[1] ),
    .B1(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__and3b_1 _3127_ (.A_N(net70),
    .B(net29),
    .C(\ih.gpio_interrupt_mask[2] ),
    .X(_2864_));
 sky130_fd_sc_hd__and3b_1 _3128_ (.A_N(net71),
    .B(net30),
    .C(\ih.gpio_interrupt_mask[3] ),
    .X(_2865_));
 sky130_fd_sc_hd__inv_2 _3129_ (.A(net74),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _3130_ (.A(net73),
    .Y(_2867_));
 sky130_fd_sc_hd__and3b_1 _3131_ (.A_N(net72),
    .B(net31),
    .C(\ih.gpio_interrupt_mask[4] ),
    .X(_2868_));
 sky130_fd_sc_hd__a31o_1 _3132_ (.A1(_2867_),
    .A2(net32),
    .A3(\ih.gpio_interrupt_mask[5] ),
    .B1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__and3b_1 _3133_ (.A_N(net75),
    .B(net34),
    .C(\ih.gpio_interrupt_mask[7] ),
    .X(_2870_));
 sky130_fd_sc_hd__a311o_1 _3134_ (.A1(_2866_),
    .A2(net33),
    .A3(\ih.gpio_interrupt_mask[6] ),
    .B1(_2869_),
    .C1(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__or4_4 _3135_ (.A(_2863_),
    .B(_2864_),
    .C(_2865_),
    .D(_2871_),
    .X(_2872_));
 sky130_fd_sc_hd__and3b_2 _3136_ (.A_N(\ih.ih.int_f.prev_data ),
    .B(\ih.ih.int_f.data_in ),
    .C(\ih.input_handler_enable ),
    .X(_2873_));
 sky130_fd_sc_hd__inv_2 _3137_ (.A(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__or2b_1 _3138_ (.A(_2872_),
    .B_N(_2860_),
    .X(_2875_));
 sky130_fd_sc_hd__nor3_1 _3139_ (.A(net1),
    .B(_2873_),
    .C(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__a32o_1 _3140_ (.A1(_2860_),
    .A2(_2872_),
    .A3(_2874_),
    .B1(_2876_),
    .B2(net204),
    .X(_0000_));
 sky130_fd_sc_hd__and3_2 _3141_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[0] ),
    .C(\cu.id.alu_opcode[3] ),
    .X(_2877_));
 sky130_fd_sc_hd__buf_2 _3142_ (.A(\cu.id.opcode[6] ),
    .X(_2878_));
 sky130_fd_sc_hd__clkbuf_4 _3143_ (.A(\cu.id.opcode[7] ),
    .X(_2879_));
 sky130_fd_sc_hd__nand2b_4 _3144_ (.A_N(_2878_),
    .B(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand3b_4 _3145_ (.A_N(\cu.id.opcode[0] ),
    .B(\cu.id.opcode[2] ),
    .C(\cu.id.opcode[1] ),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_1 _3146_ (.A(_2878_),
    .B(_2879_),
    .Y(_2882_));
 sky130_fd_sc_hd__or2_2 _3147_ (.A(_2881_),
    .B(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__and2_1 _3148_ (.A(_2880_),
    .B(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__nor2_1 _3149_ (.A(_2877_),
    .B(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__inv_2 _3150_ (.A(\cu.id.alu_opcode[1] ),
    .Y(_2886_));
 sky130_fd_sc_hd__buf_4 _3151_ (.A(\cu.id.alu_opcode[3] ),
    .X(_2887_));
 sky130_fd_sc_hd__and2_2 _3152_ (.A(\cu.id.alu_opcode[0] ),
    .B(\cu.id.opcode[0] ),
    .X(_2888_));
 sky130_fd_sc_hd__and4bb_1 _3153_ (.A_N(\cu.id.opcode[6] ),
    .B_N(\cu.id.opcode[7] ),
    .C(\cu.id.opcode[2] ),
    .D(\cu.id.opcode[1] ),
    .X(_2889_));
 sky130_fd_sc_hd__and4_2 _3154_ (.A(_2886_),
    .B(_2887_),
    .C(_2888_),
    .D(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__nor2_2 _3155_ (.A(\cu.id.opcode[6] ),
    .B(_2879_),
    .Y(_2891_));
 sky130_fd_sc_hd__and3_1 _3156_ (.A(\cu.id.opcode[0] ),
    .B(\cu.id.opcode[2] ),
    .C(\cu.id.opcode[1] ),
    .X(_2892_));
 sky130_fd_sc_hd__and2b_1 _3157_ (.A_N(\cu.id.alu_opcode[3] ),
    .B(\cu.id.alu_opcode[1] ),
    .X(_2893_));
 sky130_fd_sc_hd__and3_1 _3158_ (.A(_2891_),
    .B(_2892_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__buf_2 _3159_ (.A(\cu.id.alu_opcode[0] ),
    .X(_2895_));
 sky130_fd_sc_hd__clkbuf_4 _3160_ (.A(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__clkbuf_4 _3161_ (.A(\cu.id.opcode[0] ),
    .X(_2897_));
 sky130_fd_sc_hd__nor4b_2 _3162_ (.A(\cu.id.opcode[2] ),
    .B(\cu.id.opcode[6] ),
    .C(\cu.id.opcode[7] ),
    .D_N(\cu.id.opcode[1] ),
    .Y(_2898_));
 sky130_fd_sc_hd__nand2_4 _3163_ (.A(_2897_),
    .B(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__inv_2 _3164_ (.A(\cu.id.opcode[0] ),
    .Y(_2900_));
 sky130_fd_sc_hd__nand2_1 _3165_ (.A(_2896_),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__buf_2 _3166_ (.A(\cu.id.opcode[2] ),
    .X(_2902_));
 sky130_fd_sc_hd__buf_2 _3167_ (.A(\cu.id.opcode[1] ),
    .X(_2903_));
 sky130_fd_sc_hd__or4b_4 _3168_ (.A(_2902_),
    .B(_2878_),
    .C(_2879_),
    .D_N(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__buf_4 _3169_ (.A(\cu.id.alu_opcode[1] ),
    .X(_2905_));
 sky130_fd_sc_hd__or3b_2 _3170_ (.A(_2904_),
    .B(_2905_),
    .C_N(_2887_),
    .X(_2906_));
 sky130_fd_sc_hd__or2_1 _3171_ (.A(_2901_),
    .B(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__o21ai_1 _3172_ (.A1(_2896_),
    .A2(_2899_),
    .B1(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__or3_1 _3173_ (.A(_2890_),
    .B(_2894_),
    .C(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__nand2_4 _3174_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .Y(_2910_));
 sky130_fd_sc_hd__nor2_2 _3175_ (.A(_2896_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__and2b_2 _3176_ (.A_N(_2879_),
    .B(_2878_),
    .X(_2912_));
 sky130_fd_sc_hd__or4b_2 _3177_ (.A(_2903_),
    .B(_2878_),
    .C(_2879_),
    .D_N(_2902_),
    .X(_2913_));
 sky130_fd_sc_hd__clkbuf_4 _3178_ (.A(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__or2_1 _3179_ (.A(\cu.id.opcode[6] ),
    .B(\cu.id.opcode[7] ),
    .X(_2915_));
 sky130_fd_sc_hd__or2_2 _3180_ (.A(_2915_),
    .B(_2881_),
    .X(_2916_));
 sky130_fd_sc_hd__nand2_2 _3181_ (.A(_2914_),
    .B(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__nor2_2 _3182_ (.A(_2912_),
    .B(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__or2b_1 _3183_ (.A(_2895_),
    .B_N(_2897_),
    .X(_2919_));
 sky130_fd_sc_hd__or4bb_4 _3184_ (.A(\cu.id.opcode[2] ),
    .B(\cu.id.opcode[1] ),
    .C_N(_2878_),
    .D_N(_2879_),
    .X(_2920_));
 sky130_fd_sc_hd__nor2_1 _3185_ (.A(_2919_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__clkbuf_4 _3186_ (.A(_2887_),
    .X(_2922_));
 sky130_fd_sc_hd__and4bb_2 _3187_ (.A_N(\cu.id.opcode[2] ),
    .B_N(\cu.id.opcode[1] ),
    .C(\cu.id.opcode[6] ),
    .D(\cu.id.opcode[7] ),
    .X(_2923_));
 sky130_fd_sc_hd__nand3_2 _3188_ (.A(_2922_),
    .B(_2888_),
    .C(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__nor2_2 _3189_ (.A(_2886_),
    .B(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__nor2_1 _3190_ (.A(_2921_),
    .B(_2925_),
    .Y(_2926_));
 sky130_fd_sc_hd__or4bb_4 _3191_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .C_N(\cu.id.opcode[0] ),
    .D_N(\cu.id.alu_opcode[0] ),
    .X(_2927_));
 sky130_fd_sc_hd__and4b_2 _3192_ (.A_N(_2902_),
    .B(_2903_),
    .C(_2878_),
    .D(_2879_),
    .X(_2928_));
 sky130_fd_sc_hd__nand2b_4 _3193_ (.A_N(_2927_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__and3b_1 _3194_ (.A_N(\cu.id.cb_opcode_z[0] ),
    .B(\cu.id.cb_opcode_z[1] ),
    .C(\cu.id.cb_opcode_z[2] ),
    .X(_2930_));
 sky130_fd_sc_hd__buf_4 _3195_ (.A(\cu.id.cb_opcode_x[1] ),
    .X(_2931_));
 sky130_fd_sc_hd__inv_2 _3196_ (.A(\cu.id.cb_opcode_x[0] ),
    .Y(_2932_));
 sky130_fd_sc_hd__nor2_1 _3197_ (.A(_2931_),
    .B(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__buf_2 _3198_ (.A(_2897_),
    .X(_2934_));
 sky130_fd_sc_hd__or3b_1 _3199_ (.A(_2904_),
    .B(_2934_),
    .C_N(_2877_),
    .X(_2935_));
 sky130_fd_sc_hd__nand2_2 _3200_ (.A(_2895_),
    .B(_2897_),
    .Y(_2936_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(_2936_),
    .B(_2904_),
    .Y(_2937_));
 sky130_fd_sc_hd__nor2_2 _3202_ (.A(_2905_),
    .B(_2887_),
    .Y(_2938_));
 sky130_fd_sc_hd__and3_1 _3203_ (.A(_2891_),
    .B(_2892_),
    .C(_2938_),
    .X(_2939_));
 sky130_fd_sc_hd__nor2_1 _3204_ (.A(_2937_),
    .B(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__o311a_1 _3205_ (.A1(_2929_),
    .A2(_2930_),
    .A3(_2933_),
    .B1(_2935_),
    .C1(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__or4_1 _3206_ (.A(\cu.id.opcode[2] ),
    .B(\cu.id.opcode[1] ),
    .C(\cu.id.opcode[6] ),
    .D(\cu.id.opcode[7] ),
    .X(_2942_));
 sky130_fd_sc_hd__buf_2 _3207_ (.A(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__nor2_2 _3208_ (.A(_2902_),
    .B(_2903_),
    .Y(_2944_));
 sky130_fd_sc_hd__nor2_2 _3209_ (.A(\cu.id.alu_opcode[0] ),
    .B(\cu.id.opcode[0] ),
    .Y(_2945_));
 sky130_fd_sc_hd__nand4_4 _3210_ (.A(_2891_),
    .B(_2893_),
    .C(_2944_),
    .D(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__or3_2 _3211_ (.A(_2922_),
    .B(_2904_),
    .C(_2901_),
    .X(_2947_));
 sky130_fd_sc_hd__o211a_1 _3212_ (.A1(_2900_),
    .A2(_2943_),
    .B1(_2946_),
    .C1(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__o2111ai_4 _3213_ (.A1(_2911_),
    .A2(_2918_),
    .B1(_2926_),
    .C1(_2941_),
    .D1(_2948_),
    .Y(_2949_));
 sky130_fd_sc_hd__inv_2 _3214_ (.A(\cu.id.state[2] ),
    .Y(_2950_));
 sky130_fd_sc_hd__nand2_2 _3215_ (.A(\cu.id.state[1] ),
    .B(\cu.id.state[0] ),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_8 _3216_ (.A(_2950_),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(\cu.id.starting_int_service ),
    .Y(_2953_));
 sky130_fd_sc_hd__buf_4 _3218_ (.A(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__o311a_4 _3219_ (.A1(_2885_),
    .A2(_2909_),
    .A3(_2949_),
    .B1(_2952_),
    .C1(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__or2_2 _3220_ (.A(_2919_),
    .B(_2943_),
    .X(_2956_));
 sky130_fd_sc_hd__nand2_4 _3221_ (.A(_2899_),
    .B(_2956_),
    .Y(_0292_));
 sky130_fd_sc_hd__clkbuf_4 _3222_ (.A(\cu.id.starting_int_service ),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _3223_ (.A(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_4 _3224_ (.A(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_4 _3225_ (.A(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_4 _3226_ (.A(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__o21ai_2 _3227_ (.A1(_2936_),
    .A2(_2943_),
    .B1(_2907_),
    .Y(_0298_));
 sky130_fd_sc_hd__nand3b_2 _3228_ (.A_N(\cu.id.alu_opcode[0] ),
    .B(\cu.id.alu_opcode[3] ),
    .C(_2905_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2b_2 _3229_ (.A_N(\cu.id.opcode[7] ),
    .B(_2878_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _3230_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__and3b_1 _3231_ (.A_N(_2927_),
    .B(_2928_),
    .C(_2930_),
    .X(_0302_));
 sky130_fd_sc_hd__or4bb_1 _3232_ (.A(_2905_),
    .B(_2887_),
    .C_N(_2878_),
    .D_N(_2879_),
    .X(_0303_));
 sky130_fd_sc_hd__or4bb_1 _3233_ (.A(_2895_),
    .B(_2902_),
    .C_N(_2903_),
    .D_N(_2934_),
    .X(_0304_));
 sky130_fd_sc_hd__o2bb2a_2 _3234_ (.A1_N(_2900_),
    .A2_N(_2928_),
    .B1(_0303_),
    .B2(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__o21ai_2 _3235_ (.A1(_2905_),
    .A2(_2924_),
    .B1(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__and4b_2 _3236_ (.A_N(\cu.id.opcode[1] ),
    .B(\cu.id.opcode[6] ),
    .C(\cu.id.opcode[7] ),
    .D(\cu.id.opcode[2] ),
    .X(_0307_));
 sky130_fd_sc_hd__and3_1 _3237_ (.A(_2934_),
    .B(_2877_),
    .C(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__and3_1 _3238_ (.A(_2888_),
    .B(_2938_),
    .C(_0307_),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_4 _3239_ (.A1(_2897_),
    .A2(_2927_),
    .B1(_2920_),
    .Y(_0310_));
 sky130_fd_sc_hd__or2b_1 _3240_ (.A(\cu.id.opcode[1] ),
    .B_N(_2902_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_2 _3241_ (.A(_2895_),
    .B(_2897_),
    .X(_0312_));
 sky130_fd_sc_hd__or3_1 _3242_ (.A(_0311_),
    .B(_0312_),
    .C(_0303_),
    .X(_0313_));
 sky130_fd_sc_hd__or4b_4 _3243_ (.A(_0308_),
    .B(_0309_),
    .C(_0310_),
    .D_N(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_1 _3244_ (.A(_0306_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _3245_ (.A(_2926_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nor2_1 _3246_ (.A(_2919_),
    .B(_2942_),
    .Y(_0317_));
 sky130_fd_sc_hd__o211a_1 _3247_ (.A1(_2895_),
    .A2(_2887_),
    .B1(net150),
    .C1(_2900_),
    .X(_0318_));
 sky130_fd_sc_hd__and3b_2 _3248_ (.A_N(_2887_),
    .B(net150),
    .C(_2945_),
    .X(_0319_));
 sky130_fd_sc_hd__or4b_4 _3249_ (.A(_0317_),
    .B(_0318_),
    .C(_0319_),
    .D_N(_2916_),
    .X(_0320_));
 sky130_fd_sc_hd__nand3_2 _3250_ (.A(_2899_),
    .B(_2913_),
    .C(_2946_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor3_2 _3251_ (.A(_2881_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0322_));
 sky130_fd_sc_hd__or2_1 _3252_ (.A(\cu.id.alu_opcode[1] ),
    .B(\cu.id.alu_opcode[3] ),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _3253_ (.A(_2902_),
    .B(_2903_),
    .Y(_0324_));
 sky130_fd_sc_hd__a2111o_1 _3254_ (.A1(_2910_),
    .A2(_0323_),
    .B1(_2900_),
    .C1(_2915_),
    .D1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or4b_2 _3255_ (.A(_2890_),
    .B(_2894_),
    .C(_0322_),
    .D_N(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _3256_ (.A(_2936_),
    .B(_2943_),
    .Y(_0327_));
 sky130_fd_sc_hd__or2b_1 _3257_ (.A(_2897_),
    .B_N(_2887_),
    .X(_0328_));
 sky130_fd_sc_hd__or4bb_1 _3258_ (.A(\cu.id.opcode[0] ),
    .B(\cu.id.alu_opcode[3] ),
    .C_N(\cu.id.alu_opcode[1] ),
    .D_N(_2895_),
    .X(_0329_));
 sky130_fd_sc_hd__a21oi_1 _3259_ (.A1(_0328_),
    .A2(_0329_),
    .B1(_2943_),
    .Y(_0330_));
 sky130_fd_sc_hd__and4_1 _3260_ (.A(_2891_),
    .B(_2938_),
    .C(_2944_),
    .D(_2945_),
    .X(_0331_));
 sky130_fd_sc_hd__or3_1 _3261_ (.A(_0327_),
    .B(_0330_),
    .C(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nor4_1 _3262_ (.A(_0320_),
    .B(_0321_),
    .C(_0326_),
    .D(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _3263_ (.A(net147),
    .X(_0334_));
 sky130_fd_sc_hd__o31a_1 _3264_ (.A1(_0301_),
    .A2(_0302_),
    .A3(_0316_),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _3265_ (.A(_2911_),
    .B(_2917_),
    .X(_0336_));
 sky130_fd_sc_hd__or4_2 _3266_ (.A(_0297_),
    .B(_0298_),
    .C(_0335_),
    .D(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_2 _3267_ (.A(_0326_),
    .B(_0332_),
    .X(_0338_));
 sky130_fd_sc_hd__or3_4 _3268_ (.A(_0320_),
    .B(_0321_),
    .C(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _3269_ (.A(_2877_),
    .B(_2938_),
    .X(_0340_));
 sky130_fd_sc_hd__buf_4 _3270_ (.A(\cu.id.cb_opcode_z[1] ),
    .X(_0341_));
 sky130_fd_sc_hd__buf_4 _3271_ (.A(\cu.id.cb_opcode_z[2] ),
    .X(_0342_));
 sky130_fd_sc_hd__and3_1 _3272_ (.A(_2888_),
    .B(_2938_),
    .C(_2928_),
    .X(_0343_));
 sky130_fd_sc_hd__buf_4 _3273_ (.A(\cu.id.cb_opcode_z[0] ),
    .X(_0344_));
 sky130_fd_sc_hd__nand3_1 _3274_ (.A(_0344_),
    .B(\cu.id.cb_opcode_z[1] ),
    .C(\cu.id.cb_opcode_z[2] ),
    .Y(_0345_));
 sky130_fd_sc_hd__o211a_1 _3275_ (.A1(_0341_),
    .A2(_0342_),
    .B1(_0343_),
    .C1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_1 _3276_ (.A(_2925_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__o211a_1 _3277_ (.A1(_0300_),
    .A2(_0340_),
    .B1(_0347_),
    .C1(_0315_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_1 _3278_ (.A(_2905_),
    .B(_2922_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _3279_ (.A(_2877_),
    .B(_2938_),
    .Y(_0350_));
 sky130_fd_sc_hd__a221o_1 _3280_ (.A1(_0349_),
    .A2(_0292_),
    .B1(_0350_),
    .B2(_2917_),
    .C1(_0297_),
    .X(_0351_));
 sky130_fd_sc_hd__o21ba_2 _3281_ (.A1(_0339_),
    .A2(_0348_),
    .B1_N(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(_2895_),
    .B(_2910_),
    .Y(_0353_));
 sky130_fd_sc_hd__or2_1 _3283_ (.A(_2886_),
    .B(_2922_),
    .X(_0354_));
 sky130_fd_sc_hd__a21bo_1 _3284_ (.A1(_0341_),
    .A2(_0342_),
    .B1_N(_0344_),
    .X(_0355_));
 sky130_fd_sc_hd__a2bb2o_1 _3285_ (.A1_N(_2929_),
    .A2_N(_0355_),
    .B1(_2886_),
    .B2(_2921_),
    .X(_0356_));
 sky130_fd_sc_hd__a2111o_1 _3286_ (.A1(_0354_),
    .A2(_0292_),
    .B1(_0298_),
    .C1(_0356_),
    .D1(_2925_),
    .X(_0357_));
 sky130_fd_sc_hd__o21ba_1 _3287_ (.A1(_2918_),
    .A2(_0353_),
    .B1_N(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_4 _3288_ (.A(_2905_),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _3289_ (.A(_0341_),
    .Y(_0360_));
 sky130_fd_sc_hd__clkbuf_4 _3290_ (.A(_0343_),
    .X(_0361_));
 sky130_fd_sc_hd__and4_1 _3291_ (.A(_2891_),
    .B(_2893_),
    .C(_2944_),
    .D(_2945_),
    .X(_0362_));
 sky130_fd_sc_hd__a2111oi_1 _3292_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0362_),
    .C1(_0298_),
    .D1(_0296_),
    .Y(_0363_));
 sky130_fd_sc_hd__xnor2_4 _3293_ (.A(_2905_),
    .B(_2887_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21bai_1 _3294_ (.A1(_2921_),
    .A2(_0292_),
    .B1_N(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__o2111a_1 _3295_ (.A1(_0359_),
    .A2(_2918_),
    .B1(_0315_),
    .C1(_0363_),
    .D1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__o21a_1 _3296_ (.A1(_0297_),
    .A2(_0358_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_4 _3297_ (.A1(_0292_),
    .A2(_0337_),
    .B1(_0352_),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _3298_ (.A(_2955_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_2 _3299_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_2 _3300_ (.A(_2954_),
    .B(_0361_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _3301_ (.A(\cu.id.cb_opcode_x[1] ),
    .Y(_0372_));
 sky130_fd_sc_hd__buf_4 _3302_ (.A(\cu.id.cb_opcode_y[2] ),
    .X(_0373_));
 sky130_fd_sc_hd__buf_4 _3303_ (.A(\cu.id.cb_opcode_y[1] ),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _3304_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__and3_1 _3305_ (.A(_0372_),
    .B(_2932_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _3306_ (.A(_0371_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__and2b_1 _3307_ (.A_N(_2895_),
    .B(_2897_),
    .X(_0378_));
 sky130_fd_sc_hd__and2_2 _3308_ (.A(_0378_),
    .B(_0307_),
    .X(_0379_));
 sky130_fd_sc_hd__or3_1 _3309_ (.A(_0296_),
    .B(_2894_),
    .C(_0317_),
    .X(_0380_));
 sky130_fd_sc_hd__a211o_1 _3310_ (.A1(_0361_),
    .A2(_0376_),
    .B1(_2937_),
    .C1(_2939_),
    .X(_0381_));
 sky130_fd_sc_hd__o21bai_4 _3311_ (.A1(_2906_),
    .A2(_0312_),
    .B1_N(_0327_),
    .Y(_0382_));
 sky130_fd_sc_hd__or4_1 _3312_ (.A(_2908_),
    .B(_0380_),
    .C(_0381_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or3_2 _3313_ (.A(_0316_),
    .B(_0379_),
    .C(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _3314_ (.A(_0359_),
    .B(_2896_),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_2 _3315_ (.A(_2880_),
    .B(_2883_),
    .Y(_0386_));
 sky130_fd_sc_hd__buf_4 _3316_ (.A(\cu.id.cb_opcode_x[0] ),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _3317_ (.A(\cu.id.cb_opcode_x[1] ),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__or3_1 _3318_ (.A(_0374_),
    .B(\cu.id.cb_opcode_x[1] ),
    .C(\cu.id.cb_opcode_x[0] ),
    .X(_0389_));
 sky130_fd_sc_hd__a21oi_1 _3319_ (.A1(_0388_),
    .A2(_0389_),
    .B1(_2929_),
    .Y(_0390_));
 sky130_fd_sc_hd__a311o_1 _3320_ (.A1(_2922_),
    .A2(_0385_),
    .A3(_0386_),
    .B1(_2939_),
    .C1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__o21ai_2 _3321_ (.A1(_2890_),
    .A2(_0391_),
    .B1(_2954_),
    .Y(_0392_));
 sky130_fd_sc_hd__or2b_1 _3322_ (.A(_0384_),
    .B_N(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _3323_ (.A(_0377_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_2 _3324_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _3325_ (.A(_0373_),
    .B(_0374_),
    .X(_0396_));
 sky130_fd_sc_hd__a211o_1 _3326_ (.A1(_0375_),
    .A2(_0396_),
    .B1(\cu.id.cb_opcode_x[1] ),
    .C1(_0387_),
    .X(_0397_));
 sky130_fd_sc_hd__a311o_1 _3327_ (.A1(_0361_),
    .A2(_0388_),
    .A3(_0397_),
    .B1(_2894_),
    .C1(_2890_),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_2 _3328_ (.A1(_2896_),
    .A2(_0386_),
    .A3(_2910_),
    .B1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_2 _3329_ (.A(_2954_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_2 _3330_ (.A(_0395_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(_0378_),
    .B(_0307_),
    .Y(_0402_));
 sky130_fd_sc_hd__nor2_1 _3332_ (.A(_2912_),
    .B(_0343_),
    .Y(_0403_));
 sky130_fd_sc_hd__and4_2 _3333_ (.A(_2926_),
    .B(_0315_),
    .C(_0402_),
    .D(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__a21oi_1 _3334_ (.A1(_2883_),
    .A2(_0404_),
    .B1(_0322_),
    .Y(_0405_));
 sky130_fd_sc_hd__or3_1 _3335_ (.A(net150),
    .B(_2917_),
    .C(_0317_),
    .X(_0406_));
 sky130_fd_sc_hd__or4_4 _3336_ (.A(_0293_),
    .B(_0362_),
    .C(_0405_),
    .D(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_4 _3337_ (.A(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _3338_ (.A(_2892_),
    .B(_2944_),
    .X(_0409_));
 sky130_fd_sc_hd__o2bb2a_2 _3339_ (.A1_N(_0349_),
    .A2_N(_0327_),
    .B1(_0409_),
    .B2(_2880_),
    .X(_0410_));
 sky130_fd_sc_hd__o22a_1 _3340_ (.A1(_2880_),
    .A2(_2881_),
    .B1(_2943_),
    .B2(_2936_),
    .X(_0411_));
 sky130_fd_sc_hd__or3b_4 _3341_ (.A(_0293_),
    .B(_0410_),
    .C_N(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_2 _3342_ (.A(\cu.id.starting_int_service ),
    .B(_0411_),
    .Y(_0413_));
 sky130_fd_sc_hd__nand2_4 _3343_ (.A(_0413_),
    .B(_0410_),
    .Y(_0414_));
 sky130_fd_sc_hd__or3_1 _3344_ (.A(_2936_),
    .B(_2943_),
    .C(_0364_),
    .X(_0415_));
 sky130_fd_sc_hd__a21o_1 _3345_ (.A1(_2903_),
    .A2(_2881_),
    .B1(_2880_),
    .X(_0416_));
 sky130_fd_sc_hd__a21o_2 _3346_ (.A1(_0415_),
    .A2(_0416_),
    .B1(\cu.id.starting_int_service ),
    .X(_0417_));
 sky130_fd_sc_hd__a21bo_1 _3347_ (.A1(_2902_),
    .A2(_2903_),
    .B1_N(_2897_),
    .X(_0418_));
 sky130_fd_sc_hd__a21o_1 _3348_ (.A1(_2881_),
    .A2(_0418_),
    .B1(_2880_),
    .X(_0419_));
 sky130_fd_sc_hd__or3_1 _3349_ (.A(_2936_),
    .B(_2893_),
    .C(_2943_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_2 _3350_ (.A1(_0419_),
    .A2(_0420_),
    .B1(\cu.id.starting_int_service ),
    .X(_0421_));
 sky130_fd_sc_hd__or2_2 _3351_ (.A(_0417_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__a21oi_4 _3352_ (.A1(_0412_),
    .A2(_0414_),
    .B1(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _3353_ (.A(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__a21o_1 _3354_ (.A1(_0411_),
    .A2(_0410_),
    .B1(_0293_),
    .X(_0425_));
 sky130_fd_sc_hd__or2b_2 _3355_ (.A(_0421_),
    .B_N(_0417_),
    .X(_0426_));
 sky130_fd_sc_hd__nor2_4 _3356_ (.A(_0426_),
    .B(_0414_),
    .Y(_0427_));
 sky130_fd_sc_hd__a21o_2 _3357_ (.A1(_0424_),
    .A2(_0425_),
    .B1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__and4b_1 _3358_ (.A_N(_0417_),
    .B(_0421_),
    .C(_0413_),
    .D(_0410_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_4 _3359_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__o21bai_4 _3360_ (.A1(_0426_),
    .A2(_0412_),
    .B1_N(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a22o_1 _3361_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[0] ),
    .X(_0432_));
 sky130_fd_sc_hd__and4bb_2 _3362_ (.A_N(_0421_),
    .B_N(_0410_),
    .C(_0413_),
    .D(_0417_),
    .X(_0433_));
 sky130_fd_sc_hd__and3b_4 _3363_ (.A_N(_0412_),
    .B(_0421_),
    .C(_0417_),
    .X(_0434_));
 sky130_fd_sc_hd__and3b_2 _3364_ (.A_N(_0417_),
    .B(_0421_),
    .C(_0425_),
    .X(_0435_));
 sky130_fd_sc_hd__and3_2 _3365_ (.A(_0417_),
    .B(_0421_),
    .C(_0425_),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _3366_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0435_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[0] ),
    .X(_0437_));
 sky130_fd_sc_hd__a221o_1 _3367_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0433_),
    .B1(_0434_),
    .B2(\cu.reg_file.reg_d[0] ),
    .C1(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__and3b_4 _3368_ (.A_N(_0410_),
    .B(_0424_),
    .C(_0413_),
    .X(_0439_));
 sky130_fd_sc_hd__nor3b_4 _3369_ (.A(_0417_),
    .B(_0412_),
    .C_N(_0421_),
    .Y(_0440_));
 sky130_fd_sc_hd__a22o_1 _3370_ (.A1(\cu.reg_file.reg_mem[0] ),
    .A2(_0439_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0441_));
 sky130_fd_sc_hd__a2111o_1 _3371_ (.A1(\cu.reg_file.reg_l[0] ),
    .A2(_0423_),
    .B1(_0432_),
    .C1(_0438_),
    .D1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(_0320_),
    .Y(_0443_));
 sky130_fd_sc_hd__a21o_1 _3373_ (.A1(_0443_),
    .A2(_0404_),
    .B1(_0338_),
    .X(_0444_));
 sky130_fd_sc_hd__a221o_1 _3374_ (.A1(\cu.id.cb_opcode_y[0] ),
    .A2(_0361_),
    .B1(_0444_),
    .B2(_0344_),
    .C1(_0321_),
    .X(_0445_));
 sky130_fd_sc_hd__a21bo_1 _3375_ (.A1(_2953_),
    .A2(_0445_),
    .B1_N(_0407_),
    .X(_0446_));
 sky130_fd_sc_hd__o21ai_4 _3376_ (.A1(_0408_),
    .A2(_0442_),
    .B1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__a2111oi_1 _3377_ (.A1(_2936_),
    .A2(_0312_),
    .B1(_0323_),
    .C1(_0311_),
    .D1(_2882_),
    .Y(_0448_));
 sky130_fd_sc_hd__a32o_2 _3378_ (.A1(_2897_),
    .A2(_2877_),
    .A3(_0307_),
    .B1(_2923_),
    .B2(_0378_),
    .X(_0449_));
 sky130_fd_sc_hd__or3_1 _3379_ (.A(_0310_),
    .B(net148),
    .C(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _3380_ (.A(_2881_),
    .B(_0300_),
    .Y(_0451_));
 sky130_fd_sc_hd__and3_1 _3381_ (.A(_2887_),
    .B(_2888_),
    .C(_2923_),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _3382_ (.A(_0452_),
    .B(_0302_),
    .Y(_0453_));
 sky130_fd_sc_hd__or4b_2 _3383_ (.A(_0379_),
    .B(_0450_),
    .C(_0451_),
    .D_N(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__inv_2 _3384_ (.A(_2895_),
    .Y(_0455_));
 sky130_fd_sc_hd__or3_1 _3385_ (.A(_0455_),
    .B(_2934_),
    .C(_2904_),
    .X(_0456_));
 sky130_fd_sc_hd__or2_1 _3386_ (.A(_0299_),
    .B(_2913_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _3387_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__or4b_2 _3388_ (.A(\cu.id.starting_int_service ),
    .B(_0382_),
    .C(_0458_),
    .D_N(_2899_),
    .X(_0459_));
 sky130_fd_sc_hd__a21oi_4 _3389_ (.A1(_0334_),
    .A2(_0454_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__or3_1 _3390_ (.A(_2892_),
    .B(_0300_),
    .C(_2944_),
    .X(_0461_));
 sky130_fd_sc_hd__or3b_2 _3391_ (.A(_0346_),
    .B(_0450_),
    .C_N(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__o221a_1 _3392_ (.A1(_2899_),
    .A2(_2910_),
    .B1(_2914_),
    .B2(_0340_),
    .C1(_2953_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _3393_ (.A(_0456_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21o_1 _3394_ (.A1(_0334_),
    .A2(_0462_),
    .B1(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__nor2_2 _3395_ (.A(_0460_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__and3_2 _3396_ (.A(_2896_),
    .B(_2900_),
    .C(net150),
    .X(_0467_));
 sky130_fd_sc_hd__a21oi_1 _3397_ (.A1(_0299_),
    .A2(_0353_),
    .B1(_2914_),
    .Y(_0468_));
 sky130_fd_sc_hd__a311o_1 _3398_ (.A1(_2934_),
    .A2(_0354_),
    .A3(net150),
    .B1(_0382_),
    .C1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__nor3_4 _3399_ (.A(_0467_),
    .B(net146),
    .C(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_4 _3400_ (.A(_0310_),
    .B(_0449_),
    .Y(_0471_));
 sky130_fd_sc_hd__a21o_1 _3401_ (.A1(_2881_),
    .A2(_0418_),
    .B1(_0300_),
    .X(_0472_));
 sky130_fd_sc_hd__o221a_1 _3402_ (.A1(_2929_),
    .A2(_0355_),
    .B1(_0402_),
    .B2(_2905_),
    .C1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__a41o_4 _3403_ (.A1(net240),
    .A2(_0471_),
    .A3(_0453_),
    .A4(_0473_),
    .B1(_0293_),
    .X(_0474_));
 sky130_fd_sc_hd__a21o_1 _3404_ (.A1(_2903_),
    .A2(_2881_),
    .B1(_0300_),
    .X(_0475_));
 sky130_fd_sc_hd__o221a_1 _3405_ (.A1(\cu.id.cb_opcode_z[1] ),
    .A2(_2929_),
    .B1(_0364_),
    .B2(_0402_),
    .C1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__or4b_1 _3406_ (.A(_0452_),
    .B(_0302_),
    .C(_0450_),
    .D_N(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__a21o_1 _3407_ (.A1(_2905_),
    .A2(_0299_),
    .B1(_2914_),
    .X(_0478_));
 sky130_fd_sc_hd__o2111ai_2 _3408_ (.A1(_2899_),
    .A2(_0364_),
    .B1(_0478_),
    .C1(_2946_),
    .D1(_2953_),
    .Y(_0479_));
 sky130_fd_sc_hd__a2111o_2 _3409_ (.A1(net240),
    .A2(_0477_),
    .B1(_0479_),
    .C1(_0382_),
    .D1(_0467_),
    .X(_0480_));
 sky130_fd_sc_hd__nor3_2 _3410_ (.A(_0470_),
    .B(_0474_),
    .C(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__a2111oi_1 _3411_ (.A1(net240),
    .A2(_0477_),
    .B1(_0479_),
    .C1(_0382_),
    .D1(_0467_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor3_4 _3412_ (.A(_0470_),
    .B(_0474_),
    .C(net145),
    .Y(_0483_));
 sky130_fd_sc_hd__a21o_1 _3413_ (.A1(net147),
    .A2(_0454_),
    .B1(_0459_),
    .X(_0484_));
 sky130_fd_sc_hd__nor2_1 _3414_ (.A(_0484_),
    .B(_0465_),
    .Y(_0485_));
 sky130_fd_sc_hd__a22o_2 _3415_ (.A1(_0466_),
    .A2(_0481_),
    .B1(_0483_),
    .B2(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a21oi_4 _3416_ (.A1(net147),
    .A2(_0462_),
    .B1(_0464_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_2 _3417_ (.A(_0484_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__o2111a_4 _3418_ (.A1(_0470_),
    .A2(_0474_),
    .B1(_0480_),
    .C1(_0487_),
    .D1(_0484_),
    .X(_0489_));
 sky130_fd_sc_hd__a21o_2 _3419_ (.A1(_0481_),
    .A2(_0488_),
    .B1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__o211a_1 _3420_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .C1(\cu.reg_file.reg_l[0] ),
    .X(_0491_));
 sky130_fd_sc_hd__a221o_1 _3421_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_0486_),
    .B1(_0490_),
    .B2(\cu.reg_file.reg_e[0] ),
    .C1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__o2111a_2 _3422_ (.A1(_0470_),
    .A2(_0474_),
    .B1(net145),
    .C1(_0465_),
    .D1(_0460_),
    .X(_0493_));
 sky130_fd_sc_hd__nor2_1 _3423_ (.A(_0460_),
    .B(_0487_),
    .Y(_0494_));
 sky130_fd_sc_hd__and2_2 _3424_ (.A(_0483_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__o2111a_2 _3425_ (.A1(_0470_),
    .A2(_0474_),
    .B1(_0480_),
    .C1(_0465_),
    .D1(_0460_),
    .X(_0496_));
 sky130_fd_sc_hd__a32o_1 _3426_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0481_),
    .A3(_0494_),
    .B1(_0496_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0497_));
 sky130_fd_sc_hd__a221o_1 _3427_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_mem[0] ),
    .C1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o2111a_2 _3428_ (.A1(_0470_),
    .A2(_0474_),
    .B1(net238),
    .C1(_0487_),
    .D1(_0484_),
    .X(_0499_));
 sky130_fd_sc_hd__o2111a_2 _3429_ (.A1(_0470_),
    .A2(_0474_),
    .B1(net145),
    .C1(_0487_),
    .D1(_0460_),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _3430_ (.A(\cu.id.starting_int_service ),
    .B(net148),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_4 _3431_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__o2111a_2 _3432_ (.A1(_0470_),
    .A2(_0474_),
    .B1(_0480_),
    .C1(_0487_),
    .D1(_0460_),
    .X(_0503_));
 sky130_fd_sc_hd__a31o_1 _3433_ (.A1(_2916_),
    .A2(_2956_),
    .A3(_0305_),
    .B1(_0293_),
    .X(_0504_));
 sky130_fd_sc_hd__a21bo_2 _3434_ (.A1(_2952_),
    .A2(_0502_),
    .B1_N(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__a221o_1 _3435_ (.A1(\cu.pc.pc_o[0] ),
    .A2(_0502_),
    .B1(_0503_),
    .B2(\cu.reg_file.reg_b[0] ),
    .C1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__a221o_1 _3436_ (.A1(\alu.Cin ),
    .A2(_0499_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[0] ),
    .C1(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__inv_2 _3437_ (.A(_0505_),
    .Y(_0508_));
 sky130_fd_sc_hd__a21o_1 _3438_ (.A1(_0344_),
    .A2(_2953_),
    .B1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__o31ai_2 _3439_ (.A1(_0492_),
    .A2(_0498_),
    .A3(_0507_),
    .B1(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__xor2_2 _3440_ (.A(_0447_),
    .B(net142),
    .X(_0511_));
 sky130_fd_sc_hd__nand2_1 _3441_ (.A(\alu.Cin ),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_2 _3442_ (.A(_0395_),
    .B(_0400_),
    .Y(_0513_));
 sky130_fd_sc_hd__a21o_1 _3443_ (.A1(\alu.Cin ),
    .A2(_0513_),
    .B1(_0511_),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _3444_ (.A(_0384_),
    .B(_0392_),
    .Y(_0515_));
 sky130_fd_sc_hd__or2b_1 _3445_ (.A(_0515_),
    .B_N(_0400_),
    .X(_0516_));
 sky130_fd_sc_hd__buf_6 _3446_ (.A(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_2 _3447_ (.A(_0395_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__o211a_1 _3448_ (.A1(_0401_),
    .A2(_0512_),
    .B1(_0514_),
    .C1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_2 _3449_ (.A(_0384_),
    .B(_0392_),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _3450_ (.A(_2889_),
    .B(_0378_),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_1 _3451_ (.A(_2922_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _3452_ (.A(_0373_),
    .B(\cu.id.cb_opcode_y[0] ),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_1 _3453_ (.A(_0373_),
    .B(\cu.id.cb_opcode_y[0] ),
    .X(_0524_));
 sky130_fd_sc_hd__a311o_1 _3454_ (.A1(_0372_),
    .A2(_0523_),
    .A3(_0524_),
    .B1(_0387_),
    .C1(_2929_),
    .X(_0525_));
 sky130_fd_sc_hd__a21oi_1 _3455_ (.A1(_0359_),
    .A2(_0386_),
    .B1(_2890_),
    .Y(_0526_));
 sky130_fd_sc_hd__o221a_2 _3456_ (.A1(_2936_),
    .A2(_2904_),
    .B1(_2914_),
    .B2(_2900_),
    .C1(_2946_),
    .X(_0527_));
 sky130_fd_sc_hd__and4b_1 _3457_ (.A_N(_0522_),
    .B(_0525_),
    .C(_0526_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__buf_2 _3458_ (.A(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__or2_1 _3459_ (.A(_0400_),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _3460_ (.A(_0520_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__buf_2 _3461_ (.A(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o211a_1 _3463_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .C1(\cu.reg_file.reg_l[1] ),
    .X(_0534_));
 sky130_fd_sc_hd__and2_1 _3464_ (.A(\cu.pc.pc_o[1] ),
    .B(_0502_),
    .X(_0535_));
 sky130_fd_sc_hd__a221o_1 _3465_ (.A1(\cu.reg_file.reg_e[1] ),
    .A2(_0489_),
    .B1(_0503_),
    .B2(\cu.reg_file.reg_b[1] ),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_4 _3466_ (.A(_0505_),
    .X(_0537_));
 sky130_fd_sc_hd__a2111o_1 _3467_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_0486_),
    .B1(_0534_),
    .C1(_0536_),
    .D1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _3468_ (.A1(\cu.reg_file.reg_d[1] ),
    .A2(_0493_),
    .B1(_0499_),
    .B2(\cu.alu_f[1] ),
    .X(_0539_));
 sky130_fd_sc_hd__and2_2 _3469_ (.A(_0481_),
    .B(_0494_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _3470_ (.A(\cu.reg_file.reg_a[1] ),
    .B(_0500_),
    .X(_0541_));
 sky130_fd_sc_hd__and3_1 _3471_ (.A(\cu.reg_file.reg_e[1] ),
    .B(_0481_),
    .C(_0488_),
    .X(_0542_));
 sky130_fd_sc_hd__a32o_1 _3472_ (.A1(\cu.reg_file.reg_mem[1] ),
    .A2(_0483_),
    .A3(_0494_),
    .B1(_0496_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_0543_));
 sky130_fd_sc_hd__a2111o_1 _3473_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0540_),
    .B1(_0541_),
    .C1(_0542_),
    .D1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o21ai_1 _3474_ (.A1(_0294_),
    .A2(_0360_),
    .B1(_0537_),
    .Y(_0545_));
 sky130_fd_sc_hd__o31a_4 _3475_ (.A1(_0538_),
    .A2(_0539_),
    .A3(_0544_),
    .B1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or2_2 _3476_ (.A(_0296_),
    .B(_0529_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_2 _3477_ (.A(_0399_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__or2_2 _3478_ (.A(_0371_),
    .B(_0376_),
    .X(_0549_));
 sky130_fd_sc_hd__nor2_1 _3479_ (.A(_0549_),
    .B(_0393_),
    .Y(_0550_));
 sky130_fd_sc_hd__and2b_1 _3480_ (.A_N(_0392_),
    .B(_0384_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(_0399_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _3482_ (.A(_0529_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__or2b_1 _3483_ (.A(_0400_),
    .B_N(_0529_),
    .X(_0554_));
 sky130_fd_sc_hd__nor2_1 _3484_ (.A(_0515_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__and2_1 _3485_ (.A(_0400_),
    .B(_0547_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_0551_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _3487_ (.A(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__a2111o_4 _3488_ (.A1(_0548_),
    .A2(_0550_),
    .B1(_0553_),
    .C1(_0555_),
    .D1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__o211a_1 _3489_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .C1(\cu.reg_file.reg_l[7] ),
    .X(_0560_));
 sky130_fd_sc_hd__a221o_1 _3490_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_0486_),
    .B1(_0490_),
    .B2(\cu.reg_file.reg_e[7] ),
    .C1(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _3491_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0503_),
    .B1(_0493_),
    .B2(\cu.reg_file.reg_d[7] ),
    .X(_0562_));
 sky130_fd_sc_hd__a221o_1 _3492_ (.A1(\cu.reg_file.reg_h[7] ),
    .A2(_0496_),
    .B1(_0540_),
    .B2(\cu.reg_file.reg_sp[7] ),
    .C1(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a221o_1 _3493_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_0502_),
    .B1(_0499_),
    .B2(\cu.alu_f[7] ),
    .C1(_0505_),
    .X(_0564_));
 sky130_fd_sc_hd__a221o_1 _3494_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_0500_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_mem[7] ),
    .C1(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__o21ai_1 _3495_ (.A1(_0294_),
    .A2(_0372_),
    .B1(_0537_),
    .Y(_0566_));
 sky130_fd_sc_hd__o31a_4 _3496_ (.A1(_0561_),
    .A2(_0563_),
    .A3(_0565_),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__and3_1 _3497_ (.A(_0567_),
    .B(_0548_),
    .C(_0551_),
    .X(_0568_));
 sky130_fd_sc_hd__a221o_1 _3498_ (.A1(net142),
    .A2(_0533_),
    .B1(_0546_),
    .B2(_0559_),
    .C1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__or2_1 _3499_ (.A(_0520_),
    .B(_0554_),
    .X(_0570_));
 sky130_fd_sc_hd__buf_2 _3500_ (.A(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__and2b_1 _3501_ (.A_N(_0571_),
    .B(_0511_),
    .X(_0572_));
 sky130_fd_sc_hd__inv_2 _3502_ (.A(\alu.Cin ),
    .Y(_0573_));
 sky130_fd_sc_hd__or2_1 _3503_ (.A(_0515_),
    .B(_0530_),
    .X(_0574_));
 sky130_fd_sc_hd__a22o_1 _3504_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[2] ),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _3505_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0435_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[2] ),
    .X(_0576_));
 sky130_fd_sc_hd__a221o_1 _3506_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0433_),
    .B1(_0434_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__a22o_1 _3507_ (.A1(\cu.reg_file.reg_mem[2] ),
    .A2(_0439_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0578_));
 sky130_fd_sc_hd__a2111o_1 _3508_ (.A1(\cu.reg_file.reg_l[2] ),
    .A2(_0423_),
    .B1(_0575_),
    .C1(_0577_),
    .D1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a21oi_1 _3509_ (.A1(_0342_),
    .A2(_0338_),
    .B1(_0334_),
    .Y(_0580_));
 sky130_fd_sc_hd__a221o_1 _3510_ (.A1(\cu.id.cb_opcode_y[2] ),
    .A2(_0361_),
    .B1(_0404_),
    .B2(_0342_),
    .C1(_0339_),
    .X(_0581_));
 sky130_fd_sc_hd__or3b_1 _3511_ (.A(_0294_),
    .B(_0580_),
    .C_N(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _3512_ (.A(_0408_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__o21ai_2 _3513_ (.A1(_0408_),
    .A2(_0579_),
    .B1(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__buf_2 _3514_ (.A(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _3515_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[1] ),
    .X(_0586_));
 sky130_fd_sc_hd__a22o_1 _3516_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0433_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_0587_));
 sky130_fd_sc_hd__a221o_1 _3517_ (.A1(\cu.reg_file.reg_mem[1] ),
    .A2(_0439_),
    .B1(_0434_),
    .B2(\cu.reg_file.reg_d[1] ),
    .C1(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _3518_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0435_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[1] ),
    .X(_0589_));
 sky130_fd_sc_hd__a21o_1 _3519_ (.A1(\cu.reg_file.reg_l[1] ),
    .A2(_0423_),
    .B1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _3520_ (.A1(_0341_),
    .A2(_0338_),
    .B1(_0334_),
    .Y(_0591_));
 sky130_fd_sc_hd__a221o_1 _3521_ (.A1(\cu.id.cb_opcode_y[1] ),
    .A2(_0361_),
    .B1(_0404_),
    .B2(_0341_),
    .C1(_0339_),
    .X(_0592_));
 sky130_fd_sc_hd__or3b_1 _3522_ (.A(_0293_),
    .B(_0591_),
    .C_N(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__nand2_1 _3523_ (.A(_0407_),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__o41a_4 _3524_ (.A1(_0407_),
    .A2(_0586_),
    .A3(_0588_),
    .A4(_0590_),
    .B1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_4 _3525_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__and3_1 _3527_ (.A(_0447_),
    .B(_0585_),
    .C(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or2b_1 _3528_ (.A(_0520_),
    .B_N(_0556_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_4 _3529_ (.A(_0549_),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _3530_ (.A(_0598_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__or2_1 _3531_ (.A(_0447_),
    .B(_0600_),
    .X(_0602_));
 sky130_fd_sc_hd__or2_2 _3532_ (.A(_0399_),
    .B(_0547_),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_4 _3533_ (.A(_0520_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__nor2_2 _3534_ (.A(_0600_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__a31o_1 _3535_ (.A1(net142),
    .A2(_0601_),
    .A3(_0602_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_2 _3536_ (.A(_0377_),
    .B(_0599_),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _3537_ (.A(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__or3_1 _3538_ (.A(_0549_),
    .B(_0393_),
    .C(_0530_),
    .X(_0609_));
 sky130_fd_sc_hd__buf_2 _3539_ (.A(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__o21a_1 _3540_ (.A1(_0447_),
    .A2(_0608_),
    .B1(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__or3_1 _3541_ (.A(net142),
    .B(_0598_),
    .C(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_1 _3542_ (.A(_0550_),
    .B(_0556_),
    .Y(_0613_));
 sky130_fd_sc_hd__o2111a_1 _3543_ (.A1(_0573_),
    .A2(_0574_),
    .B1(_0606_),
    .C1(_0612_),
    .D1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or4b_1 _3544_ (.A(_0519_),
    .B(_0569_),
    .C(_0572_),
    .D_N(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__buf_4 _3545_ (.A(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_4 _3546_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_1 _3548_ (.A(_0377_),
    .B(_0393_),
    .Y(_0619_));
 sky130_fd_sc_hd__o21a_1 _3549_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _3550_ (.A1(\cu.reg_file.reg_e[6] ),
    .A2(_0490_),
    .B1(_0620_),
    .B2(\cu.reg_file.reg_l[6] ),
    .X(_0621_));
 sky130_fd_sc_hd__a21o_1 _3551_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_0486_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_4 _3552_ (.A(_0540_),
    .X(_0623_));
 sky130_fd_sc_hd__buf_2 _3553_ (.A(_0499_),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _3554_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0493_),
    .B1(_0624_),
    .B2(\cu.alu_f[6] ),
    .X(_0625_));
 sky130_fd_sc_hd__a221o_1 _3555_ (.A1(\cu.reg_file.reg_h[6] ),
    .A2(_0496_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[6] ),
    .C1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__buf_2 _3556_ (.A(_0495_),
    .X(_0627_));
 sky130_fd_sc_hd__a221o_1 _3557_ (.A1(\cu.pc.pc_o[6] ),
    .A2(_0502_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[6] ),
    .C1(_0537_),
    .X(_0628_));
 sky130_fd_sc_hd__a221o_1 _3558_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0503_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[6] ),
    .C1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__o21ai_1 _3559_ (.A1(_0295_),
    .A2(_2932_),
    .B1(_0537_),
    .Y(_0630_));
 sky130_fd_sc_hd__o31a_4 _3560_ (.A1(_0622_),
    .A2(_0626_),
    .A3(_0629_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _3561_ (.A(_0443_),
    .B(_0404_),
    .Y(_0632_));
 sky130_fd_sc_hd__o21ba_1 _3562_ (.A1(_0321_),
    .A2(_0632_),
    .B1_N(_0338_),
    .X(_0633_));
 sky130_fd_sc_hd__or3_1 _3563_ (.A(_0295_),
    .B(_2932_),
    .C(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _3564_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[6] ),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_8 _3565_ (.A(_0439_),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _3566_ (.A1(\cu.reg_file.reg_mem[6] ),
    .A2(_0636_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[6] ),
    .X(_0637_));
 sky130_fd_sc_hd__a2111o_1 _3567_ (.A1(\cu.reg_file.reg_l[6] ),
    .A2(_0423_),
    .B1(_0635_),
    .C1(_0637_),
    .D1(_0408_),
    .X(_0638_));
 sky130_fd_sc_hd__buf_2 _3568_ (.A(_0433_),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _3569_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0434_),
    .B1(_0435_),
    .B2(\cu.reg_file.reg_b[6] ),
    .X(_0640_));
 sky130_fd_sc_hd__a221o_1 _3570_ (.A1(\cu.reg_file.reg_sp[6] ),
    .A2(_0639_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[6] ),
    .C1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__o2bb2a_2 _3571_ (.A1_N(_0408_),
    .A2_N(_0634_),
    .B1(_0638_),
    .B2(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__xnor2_2 _3572_ (.A(_0631_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _3573_ (.A(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__or3b_1 _3574_ (.A(_0295_),
    .B(_0633_),
    .C_N(_0373_),
    .X(_0645_));
 sky130_fd_sc_hd__a22o_1 _3575_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0434_),
    .B1(_0435_),
    .B2(\cu.reg_file.reg_b[5] ),
    .X(_0646_));
 sky130_fd_sc_hd__a221o_1 _3576_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0639_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_1 _3577_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[5] ),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _3578_ (.A1(\cu.reg_file.reg_mem[5] ),
    .A2(_0636_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[5] ),
    .X(_0649_));
 sky130_fd_sc_hd__a2111o_1 _3579_ (.A1(\cu.reg_file.reg_l[5] ),
    .A2(_0423_),
    .B1(_0648_),
    .C1(_0649_),
    .D1(_0408_),
    .X(_0650_));
 sky130_fd_sc_hd__o2bb2a_2 _3580_ (.A1_N(_0408_),
    .A2_N(_0645_),
    .B1(_0647_),
    .B2(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__clkbuf_8 _3581_ (.A(_0508_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_1 _3582_ (.A(\ih.interrupt_source[3] ),
    .B(\ih.interrupt_source[1] ),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(\cu.id.cb_opcode_y[2] ),
    .A1(_0653_),
    .S(_0294_),
    .X(_0654_));
 sky130_fd_sc_hd__and2_1 _3584_ (.A(\cu.pc.pc_o[5] ),
    .B(_0502_),
    .X(_0655_));
 sky130_fd_sc_hd__a221o_1 _3585_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0493_),
    .B1(_0624_),
    .B2(\cu.alu_f[5] ),
    .C1(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _3586_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0503_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[5] ),
    .X(_0657_));
 sky130_fd_sc_hd__a221o_1 _3587_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0540_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_mem[5] ),
    .C1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a221o_1 _3588_ (.A1(\cu.reg_file.reg_e[5] ),
    .A2(_0490_),
    .B1(_0496_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_0537_),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _3589_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_0486_),
    .B1(_0620_),
    .B2(\cu.reg_file.reg_l[5] ),
    .X(_0660_));
 sky130_fd_sc_hd__or3_1 _3590_ (.A(_0658_),
    .B(_0659_),
    .C(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__o22a_4 _3591_ (.A1(_0652_),
    .A2(_0654_),
    .B1(_0656_),
    .B2(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__xnor2_4 _3592_ (.A(_0651_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__or3b_1 _3593_ (.A(_0294_),
    .B(_0633_),
    .C_N(_0374_),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _3594_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_0434_),
    .B1(_0435_),
    .B2(\cu.reg_file.reg_b[4] ),
    .X(_0665_));
 sky130_fd_sc_hd__a221o_1 _3595_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0433_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[4] ),
    .C1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__a22o_1 _3596_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[4] ),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _3597_ (.A1(\cu.reg_file.reg_mem[4] ),
    .A2(_0439_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[4] ),
    .X(_0668_));
 sky130_fd_sc_hd__a2111o_1 _3598_ (.A1(\cu.reg_file.reg_l[4] ),
    .A2(_0423_),
    .B1(_0667_),
    .C1(_0668_),
    .D1(_0408_),
    .X(_0669_));
 sky130_fd_sc_hd__o2bb2a_1 _3599_ (.A1_N(_0408_),
    .A2_N(_0664_),
    .B1(_0666_),
    .B2(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(\ih.interrupt_source[2] ),
    .B(\ih.interrupt_source[3] ),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(_0374_),
    .A1(_0671_),
    .S(_0294_),
    .X(_0672_));
 sky130_fd_sc_hd__a22o_1 _3602_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_0486_),
    .B1(_0490_),
    .B2(\cu.reg_file.reg_e[4] ),
    .X(_0673_));
 sky130_fd_sc_hd__a21o_1 _3603_ (.A1(\cu.reg_file.reg_l[4] ),
    .A2(_0620_),
    .B1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__a22o_1 _3604_ (.A1(\cu.reg_file.reg_h[4] ),
    .A2(_0496_),
    .B1(_0499_),
    .B2(\cu.alu_f[4] ),
    .X(_0675_));
 sky130_fd_sc_hd__a221o_1 _3605_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0503_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_mem[4] ),
    .C1(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__a221o_1 _3606_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_0502_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[4] ),
    .C1(_0505_),
    .X(_0677_));
 sky130_fd_sc_hd__a221o_1 _3607_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0540_),
    .B1(_0493_),
    .B2(\cu.reg_file.reg_d[4] ),
    .C1(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__or2_1 _3608_ (.A(_0676_),
    .B(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__o22a_2 _3609_ (.A1(_0652_),
    .A2(_0672_),
    .B1(_0674_),
    .B2(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__and2b_1 _3610_ (.A_N(_0670_),
    .B(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__and2b_1 _3611_ (.A_N(_0680_),
    .B(_0670_),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_2 _3612_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_1 _3613_ (.A(_0663_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__o211a_1 _3614_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .C1(\cu.reg_file.reg_l[3] ),
    .X(_0685_));
 sky130_fd_sc_hd__a221o_1 _3615_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_0486_),
    .B1(_0490_),
    .B2(\cu.reg_file.reg_e[3] ),
    .C1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a22o_1 _3616_ (.A1(\cu.reg_file.reg_h[3] ),
    .A2(_0496_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[3] ),
    .X(_0687_));
 sky130_fd_sc_hd__a221o_1 _3617_ (.A1(\cu.alu_f[3] ),
    .A2(_0499_),
    .B1(_0495_),
    .B2(\cu.reg_file.reg_mem[3] ),
    .C1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__a221o_1 _3618_ (.A1(\cu.pc.pc_o[3] ),
    .A2(_0502_),
    .B1(_0503_),
    .B2(\cu.reg_file.reg_b[3] ),
    .C1(_0537_),
    .X(_0689_));
 sky130_fd_sc_hd__a221o_1 _3619_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0540_),
    .B1(_0493_),
    .B2(\cu.reg_file.reg_d[3] ),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(\cu.id.cb_opcode_y[0] ),
    .Y(_0691_));
 sky130_fd_sc_hd__o21ai_1 _3621_ (.A1(_0294_),
    .A2(_0691_),
    .B1(_0537_),
    .Y(_0692_));
 sky130_fd_sc_hd__o31a_4 _3622_ (.A1(_0686_),
    .A2(_0688_),
    .A3(_0690_),
    .B1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__or3_1 _3623_ (.A(_0294_),
    .B(_0691_),
    .C(_0633_),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _3624_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[3] ),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _3625_ (.A1(\cu.reg_file.reg_mem[3] ),
    .A2(_0439_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[3] ),
    .X(_0696_));
 sky130_fd_sc_hd__a2111o_1 _3626_ (.A1(\cu.reg_file.reg_l[3] ),
    .A2(_0423_),
    .B1(_0695_),
    .C1(_0696_),
    .D1(_0407_),
    .X(_0697_));
 sky130_fd_sc_hd__a22o_1 _3627_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_0434_),
    .B1(_0435_),
    .B2(\cu.reg_file.reg_b[3] ),
    .X(_0698_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0433_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__o2bb2a_2 _3629_ (.A1_N(_0408_),
    .A2_N(_0694_),
    .B1(_0697_),
    .B2(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nor2_1 _3630_ (.A(_0693_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__o211a_1 _3631_ (.A1(_0466_),
    .A2(_0488_),
    .B1(_0483_),
    .C1(\cu.reg_file.reg_l[2] ),
    .X(_0702_));
 sky130_fd_sc_hd__a221o_1 _3632_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_0486_),
    .B1(_0490_),
    .B2(\cu.reg_file.reg_e[2] ),
    .C1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _3633_ (.A1(\cu.reg_file.reg_h[2] ),
    .A2(_0496_),
    .B1(_0500_),
    .B2(\cu.reg_file.reg_a[2] ),
    .X(_0704_));
 sky130_fd_sc_hd__a221o_1 _3634_ (.A1(\cu.alu_f[2] ),
    .A2(_0499_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[2] ),
    .C1(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__a221o_1 _3635_ (.A1(\cu.pc.pc_o[2] ),
    .A2(_0502_),
    .B1(_0503_),
    .B2(\cu.reg_file.reg_b[2] ),
    .C1(_0537_),
    .X(_0706_));
 sky130_fd_sc_hd__a221o_1 _3636_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0623_),
    .B1(_0493_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__a21o_1 _3637_ (.A1(_2954_),
    .A2(_0342_),
    .B1(_0508_),
    .X(_0708_));
 sky130_fd_sc_hd__o31ai_4 _3638_ (.A1(_0703_),
    .A2(_0705_),
    .A3(_0707_),
    .B1(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(_0584_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__xnor2_4 _3640_ (.A(_0546_),
    .B(_0595_),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _3641_ (.A(_0447_),
    .B(net142),
    .X(_0712_));
 sky130_fd_sc_hd__a2bb2o_1 _3642_ (.A1_N(_0711_),
    .A2_N(_0712_),
    .B1(_0546_),
    .B2(_0596_),
    .X(_0713_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(_0584_),
    .B(_0709_),
    .Y(_0714_));
 sky130_fd_sc_hd__a21oi_1 _3644_ (.A1(_0710_),
    .A2(_0713_),
    .B1(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(_0693_),
    .B(_0700_),
    .Y(_0716_));
 sky130_fd_sc_hd__o21ai_2 _3646_ (.A1(_0701_),
    .A2(_0715_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_1 _3647_ (.A(_0651_),
    .B(_0662_),
    .Y(_0718_));
 sky130_fd_sc_hd__and2_1 _3648_ (.A(_0670_),
    .B(_0680_),
    .X(_0719_));
 sky130_fd_sc_hd__and2b_1 _3649_ (.A_N(_0718_),
    .B(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__a221o_1 _3650_ (.A1(_0651_),
    .A2(_0662_),
    .B1(_0684_),
    .B2(_0717_),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__or3_1 _3651_ (.A(_0293_),
    .B(_0372_),
    .C(_0633_),
    .X(_0722_));
 sky130_fd_sc_hd__a22o_1 _3652_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\cu.reg_file.reg_e[7] ),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _3653_ (.A1(\cu.reg_file.reg_mem[7] ),
    .A2(_0439_),
    .B1(_0436_),
    .B2(\cu.reg_file.reg_a[7] ),
    .X(_0724_));
 sky130_fd_sc_hd__a2111o_1 _3654_ (.A1(\cu.reg_file.reg_l[7] ),
    .A2(_0423_),
    .B1(_0723_),
    .C1(_0724_),
    .D1(_0407_),
    .X(_0725_));
 sky130_fd_sc_hd__a22o_1 _3655_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_0434_),
    .B1(_0435_),
    .B2(\cu.reg_file.reg_b[7] ),
    .X(_0726_));
 sky130_fd_sc_hd__a221o_1 _3656_ (.A1(\cu.reg_file.reg_sp[7] ),
    .A2(_0433_),
    .B1(_0440_),
    .B2(\cu.reg_file.reg_h[7] ),
    .C1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__o2bb2a_2 _3657_ (.A1_N(_0407_),
    .A2_N(_0722_),
    .B1(_0725_),
    .B2(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(_0567_),
    .B(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _3659_ (.A(_0567_),
    .B(_0728_),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _3660_ (.A(_0729_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__buf_2 _3661_ (.A(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__inv_2 _3662_ (.A(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__and2_1 _3663_ (.A(_0631_),
    .B(_0642_),
    .X(_0734_));
 sky130_fd_sc_hd__and2b_1 _3664_ (.A_N(_0730_),
    .B(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__a311o_1 _3665_ (.A1(_0644_),
    .A2(_0721_),
    .A3(_0733_),
    .B1(_0735_),
    .C1(_0729_),
    .X(_0736_));
 sky130_fd_sc_hd__and3_1 _3666_ (.A(_2954_),
    .B(_2916_),
    .C(_0537_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_4 _3667_ (.A(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__buf_4 _3668_ (.A(_0502_),
    .X(_0739_));
 sky130_fd_sc_hd__and2_2 _3669_ (.A(_0466_),
    .B(_0483_),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _3670_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0741_));
 sky130_fd_sc_hd__and2_2 _3671_ (.A(_0466_),
    .B(_0481_),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _3672_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[8] ),
    .X(_0743_));
 sky130_fd_sc_hd__a211o_1 _3673_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_0739_),
    .B1(_0741_),
    .C1(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a221o_1 _3674_ (.A1(\cu.reg_file.reg_a[0] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[8] ),
    .C1(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__a22oi_4 _3675_ (.A1(\cu.id.imm_i[8] ),
    .A2(_0738_),
    .B1(_0745_),
    .B2(_0652_),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_4 _3676_ (.A(_0422_),
    .B(_0414_),
    .Y(_0747_));
 sky130_fd_sc_hd__a22o_1 _3677_ (.A1(\cu.reg_file.reg_sp[8] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[0] ),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _3678_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[0] ),
    .X(_0749_));
 sky130_fd_sc_hd__a211oi_4 _3679_ (.A1(\cu.reg_file.reg_mem[8] ),
    .A2(_0636_),
    .B1(_0748_),
    .C1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__xor2_2 _3680_ (.A(_0746_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__xor2_1 _3681_ (.A(_0736_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__xnor2_1 _3682_ (.A(_0644_),
    .B(_0721_),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_2 _3683_ (.A(_0683_),
    .Y(_0754_));
 sky130_fd_sc_hd__a21oi_1 _3684_ (.A1(_0717_),
    .A2(_0754_),
    .B1(_0719_),
    .Y(_0755_));
 sky130_fd_sc_hd__xnor2_1 _3685_ (.A(_0663_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _3686_ (.A(_0512_),
    .B(_0711_),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2b_2 _3687_ (.A_N(_0714_),
    .B(_0710_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _3688_ (.A(_0713_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _3689_ (.A(_0757_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__xor2_1 _3690_ (.A(_0693_),
    .B(_0700_),
    .X(_0761_));
 sky130_fd_sc_hd__inv_2 _3691_ (.A(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__xnor2_1 _3692_ (.A(_0715_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(_0760_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__xnor2_1 _3694_ (.A(_0717_),
    .B(_0683_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _3695_ (.A(_0764_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__or3_2 _3696_ (.A(_0753_),
    .B(_0756_),
    .C(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__a21o_1 _3697_ (.A1(_0644_),
    .A2(_0721_),
    .B1(_0734_),
    .X(_0768_));
 sky130_fd_sc_hd__xnor2_2 _3698_ (.A(_0768_),
    .B(_0733_),
    .Y(_0769_));
 sky130_fd_sc_hd__or3b_1 _3699_ (.A(_0767_),
    .B(_0769_),
    .C_N(_0752_),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _3700_ (.A(_0513_),
    .B(_0529_),
    .X(_0771_));
 sky130_fd_sc_hd__clkbuf_4 _3701_ (.A(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__or2_2 _3702_ (.A(_0515_),
    .B(_0603_),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_0619_),
    .B(_0548_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_4 _3704_ (.A(_0773_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__nor2_2 _3705_ (.A(_0513_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__a21o_1 _3706_ (.A1(_0770_),
    .A2(_0772_),
    .B1(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_2 _3707_ (.A(_0513_),
    .B(_0529_),
    .Y(_0778_));
 sky130_fd_sc_hd__nor4_1 _3708_ (.A(_0767_),
    .B(_0769_),
    .C(_0752_),
    .D(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__or2b_1 _3709_ (.A(_0447_),
    .B_N(net142),
    .X(_0780_));
 sky130_fd_sc_hd__and2b_1 _3710_ (.A_N(_0595_),
    .B(_0546_),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_1 _3711_ (.A1(_0780_),
    .A2(_0711_),
    .B1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__and2b_1 _3712_ (.A_N(_0709_),
    .B(_0584_),
    .X(_0783_));
 sky130_fd_sc_hd__and2b_1 _3713_ (.A_N(_0761_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__and2b_1 _3714_ (.A_N(_0700_),
    .B(_0693_),
    .X(_0785_));
 sky130_fd_sc_hd__a311o_2 _3715_ (.A1(_0758_),
    .A2(_0762_),
    .A3(_0782_),
    .B1(_0784_),
    .C1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__and2_1 _3716_ (.A(_0643_),
    .B(_0732_),
    .X(_0787_));
 sky130_fd_sc_hd__nand4_1 _3717_ (.A(_0663_),
    .B(_0683_),
    .C(_0786_),
    .D(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__and2b_1 _3718_ (.A_N(_0642_),
    .B(_0631_),
    .X(_0789_));
 sky130_fd_sc_hd__inv_2 _3719_ (.A(_0567_),
    .Y(_0790_));
 sky130_fd_sc_hd__o2bb2a_1 _3720_ (.A1_N(_0732_),
    .A2_N(_0789_),
    .B1(_0728_),
    .B2(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__and2b_1 _3721_ (.A_N(_0651_),
    .B(_0662_),
    .X(_0792_));
 sky130_fd_sc_hd__a21o_1 _3722_ (.A1(_0663_),
    .A2(_0681_),
    .B1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _3723_ (.A(_0787_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__a31o_1 _3724_ (.A1(_0788_),
    .A2(_0791_),
    .A3(_0794_),
    .B1(_0751_),
    .X(_0795_));
 sky130_fd_sc_hd__nand4_1 _3725_ (.A(_0751_),
    .B(_0788_),
    .C(_0791_),
    .D(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__and2_1 _3726_ (.A(_0795_),
    .B(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__a31o_1 _3727_ (.A1(_0663_),
    .A2(_0683_),
    .A3(_0786_),
    .B1(_0793_),
    .X(_0798_));
 sky130_fd_sc_hd__a21oi_1 _3728_ (.A1(_0643_),
    .A2(_0798_),
    .B1(_0789_),
    .Y(_0799_));
 sky130_fd_sc_hd__xnor2_2 _3729_ (.A(_0732_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_1 _3730_ (.A(_0644_),
    .B(_0798_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21oi_1 _3731_ (.A1(_0683_),
    .A2(_0786_),
    .B1(_0681_),
    .Y(_0802_));
 sky130_fd_sc_hd__xnor2_1 _3732_ (.A(_0663_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__xnor2_1 _3733_ (.A(_0754_),
    .B(_0786_),
    .Y(_0804_));
 sky130_fd_sc_hd__xor2_1 _3734_ (.A(_0758_),
    .B(_0782_),
    .X(_0805_));
 sky130_fd_sc_hd__or3b_1 _3735_ (.A(_0573_),
    .B(_0511_),
    .C_N(_0711_),
    .X(_0806_));
 sky130_fd_sc_hd__or2_1 _3736_ (.A(_0805_),
    .B(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__a21oi_1 _3737_ (.A1(_0758_),
    .A2(_0782_),
    .B1(_0783_),
    .Y(_0808_));
 sky130_fd_sc_hd__xnor2_2 _3738_ (.A(_0762_),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__or3_1 _3739_ (.A(_0804_),
    .B(_0807_),
    .C(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__or3_2 _3740_ (.A(_0801_),
    .B(_0803_),
    .C(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__or3_1 _3741_ (.A(_0800_),
    .B(_0811_),
    .C(_0797_),
    .X(_0812_));
 sky130_fd_sc_hd__o21ai_1 _3742_ (.A1(_0800_),
    .A2(_0811_),
    .B1(_0797_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand2_1 _3743_ (.A(_0812_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _3744_ (.A(_0401_),
    .B(_0529_),
    .Y(_0815_));
 sky130_fd_sc_hd__buf_2 _3745_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a22o_1 _3746_ (.A1(_0775_),
    .A2(_0797_),
    .B1(_0814_),
    .B2(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a211o_1 _3747_ (.A1(_0752_),
    .A2(_0777_),
    .B1(_0779_),
    .C1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(_0510_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _3749_ (.A(_0603_),
    .B(_0554_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_0613_),
    .B(_0574_),
    .Y(_0821_));
 sky130_fd_sc_hd__a21o_2 _3751_ (.A1(_0551_),
    .A2(_0820_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__a22o_1 _3752_ (.A1(_0819_),
    .A2(_0559_),
    .B1(_0822_),
    .B2(_0567_),
    .X(_0823_));
 sky130_fd_sc_hd__and3_2 _3753_ (.A(_0384_),
    .B(_0392_),
    .C(_0400_),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _3754_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[7] ),
    .X(_0825_));
 sky130_fd_sc_hd__a22o_1 _3755_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[15] ),
    .X(_0826_));
 sky130_fd_sc_hd__a211o_1 _3756_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_0739_),
    .B1(_0825_),
    .C1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__a221o_1 _3757_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[15] ),
    .C1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__a22oi_4 _3758_ (.A1(\cu.id.imm_i[15] ),
    .A2(_0738_),
    .B1(_0828_),
    .B2(_0652_),
    .Y(_0829_));
 sky130_fd_sc_hd__a22o_1 _3759_ (.A1(\cu.reg_file.reg_sp[15] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[7] ),
    .X(_0830_));
 sky130_fd_sc_hd__a22o_1 _3760_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[7] ),
    .X(_0831_));
 sky130_fd_sc_hd__a211oi_4 _3761_ (.A1(\cu.reg_file.reg_mem[15] ),
    .A2(_0636_),
    .B1(_0830_),
    .C1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__xnor2_4 _3762_ (.A(_0829_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a22o_1 _3763_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[6] ),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _3764_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[14] ),
    .X(_0835_));
 sky130_fd_sc_hd__a211o_1 _3765_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_0739_),
    .B1(_0834_),
    .C1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _3766_ (.A1(\cu.reg_file.reg_a[6] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[14] ),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__a22oi_4 _3767_ (.A1(\cu.id.imm_i[14] ),
    .A2(_0738_),
    .B1(_0837_),
    .B2(_0652_),
    .Y(_0838_));
 sky130_fd_sc_hd__a22o_1 _3768_ (.A1(\cu.reg_file.reg_sp[14] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[6] ),
    .X(_0839_));
 sky130_fd_sc_hd__a22o_1 _3769_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[6] ),
    .X(_0840_));
 sky130_fd_sc_hd__a211oi_2 _3770_ (.A1(\cu.reg_file.reg_mem[14] ),
    .A2(_0636_),
    .B1(_0839_),
    .C1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__and2b_1 _3771_ (.A_N(_0838_),
    .B(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__or2b_1 _3772_ (.A(_0841_),
    .B_N(_0838_),
    .X(_0843_));
 sky130_fd_sc_hd__and2b_1 _3773_ (.A_N(_0842_),
    .B(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__inv_2 _3774_ (.A(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__a22o_1 _3775_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[5] ),
    .X(_0846_));
 sky130_fd_sc_hd__a22o_1 _3776_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[13] ),
    .X(_0847_));
 sky130_fd_sc_hd__a211o_1 _3777_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_0739_),
    .B1(_0846_),
    .C1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__a221o_1 _3778_ (.A1(\cu.reg_file.reg_a[5] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[13] ),
    .C1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__a22oi_4 _3779_ (.A1(\cu.id.imm_i[13] ),
    .A2(_0738_),
    .B1(_0849_),
    .B2(_0652_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _3780_ (.A1(\cu.reg_file.reg_sp[13] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[5] ),
    .X(_0851_));
 sky130_fd_sc_hd__a22o_1 _3781_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[5] ),
    .X(_0852_));
 sky130_fd_sc_hd__a211oi_2 _3782_ (.A1(\cu.reg_file.reg_mem[13] ),
    .A2(_0636_),
    .B1(_0851_),
    .C1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__or2b_1 _3783_ (.A(_0850_),
    .B_N(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__or2b_1 _3784_ (.A(_0853_),
    .B_N(_0850_),
    .X(_0855_));
 sky130_fd_sc_hd__nand2_2 _3785_ (.A(_0854_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a22o_1 _3786_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[4] ),
    .X(_0857_));
 sky130_fd_sc_hd__a22o_1 _3787_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[12] ),
    .X(_0858_));
 sky130_fd_sc_hd__a211o_1 _3788_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_0739_),
    .B1(_0857_),
    .C1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__a221o_1 _3789_ (.A1(\cu.reg_file.reg_a[4] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[12] ),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a22oi_4 _3790_ (.A1(\cu.id.imm_i[12] ),
    .A2(_0738_),
    .B1(_0860_),
    .B2(_0652_),
    .Y(_0861_));
 sky130_fd_sc_hd__a22o_1 _3791_ (.A1(\cu.reg_file.reg_sp[12] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[4] ),
    .X(_0862_));
 sky130_fd_sc_hd__a22o_1 _3792_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[4] ),
    .X(_0863_));
 sky130_fd_sc_hd__a211oi_4 _3793_ (.A1(\cu.reg_file.reg_mem[12] ),
    .A2(_0636_),
    .B1(_0862_),
    .C1(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__xnor2_2 _3794_ (.A(_0861_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__inv_2 _3795_ (.A(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a22o_1 _3796_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[11] ),
    .X(_0867_));
 sky130_fd_sc_hd__a221o_1 _3797_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__a21o_1 _3798_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_0739_),
    .B1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a221o_1 _3799_ (.A1(\cu.reg_file.reg_a[3] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[11] ),
    .C1(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a22oi_2 _3800_ (.A1(\cu.id.imm_i[11] ),
    .A2(_0738_),
    .B1(_0870_),
    .B2(_0652_),
    .Y(_0871_));
 sky130_fd_sc_hd__a22o_1 _3801_ (.A1(\cu.reg_file.reg_sp[11] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[3] ),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _3802_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[3] ),
    .X(_0873_));
 sky130_fd_sc_hd__a211oi_1 _3803_ (.A1(\cu.reg_file.reg_mem[11] ),
    .A2(_0636_),
    .B1(_0872_),
    .C1(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__and2b_1 _3804_ (.A_N(_0871_),
    .B(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__and2b_1 _3805_ (.A_N(_0874_),
    .B(_0871_),
    .X(_0876_));
 sky130_fd_sc_hd__or2_1 _3806_ (.A(_0875_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _3807_ (.A1(\cu.reg_file.reg_d[2] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0878_));
 sky130_fd_sc_hd__a22o_1 _3808_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[10] ),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _3809_ (.A1(\cu.pc.pc_o[10] ),
    .A2(_0739_),
    .B1(_0878_),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a221o_1 _3810_ (.A1(\cu.reg_file.reg_a[2] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[10] ),
    .C1(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__a22o_1 _3811_ (.A1(\cu.id.imm_i[10] ),
    .A2(_0738_),
    .B1(_0881_),
    .B2(_0652_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _3812_ (.A1(\cu.reg_file.reg_sp[10] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[2] ),
    .X(_0883_));
 sky130_fd_sc_hd__a22o_1 _3813_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[2] ),
    .X(_0884_));
 sky130_fd_sc_hd__a211oi_2 _3814_ (.A1(\cu.reg_file.reg_mem[10] ),
    .A2(_0636_),
    .B1(_0883_),
    .C1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__xor2_1 _3815_ (.A(_0882_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__inv_2 _3816_ (.A(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a22o_1 _3817_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0742_),
    .B1(_0623_),
    .B2(\cu.reg_file.reg_sp[9] ),
    .X(_0888_));
 sky130_fd_sc_hd__a221o_1 _3818_ (.A1(\cu.reg_file.reg_d[1] ),
    .A2(_0489_),
    .B1(_0740_),
    .B2(\cu.reg_file.reg_h[1] ),
    .C1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__a21o_1 _3819_ (.A1(\cu.pc.pc_o[9] ),
    .A2(_0739_),
    .B1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _3820_ (.A1(\cu.reg_file.reg_a[1] ),
    .A2(_0624_),
    .B1(_0627_),
    .B2(\cu.reg_file.reg_mem[9] ),
    .C1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__a22oi_2 _3821_ (.A1(\cu.id.imm_i[9] ),
    .A2(_0738_),
    .B1(_0891_),
    .B2(_0652_),
    .Y(_0892_));
 sky130_fd_sc_hd__a22o_1 _3822_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_0639_),
    .B1(_0747_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_0893_));
 sky130_fd_sc_hd__a22o_1 _3823_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\cu.reg_file.reg_d[1] ),
    .X(_0894_));
 sky130_fd_sc_hd__a211oi_2 _3824_ (.A1(\cu.reg_file.reg_mem[9] ),
    .A2(_0636_),
    .B1(_0893_),
    .C1(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2b_1 _3825_ (.A(_0892_),
    .B_N(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or2b_1 _3826_ (.A(_0895_),
    .B_N(_0892_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_2 _3827_ (.A(_0896_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nor2_1 _3828_ (.A(_0746_),
    .B(_0750_),
    .Y(_0899_));
 sky130_fd_sc_hd__a2bb2o_1 _3829_ (.A1_N(_0892_),
    .A2_N(_0895_),
    .B1(_0898_),
    .B2(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__a31o_1 _3830_ (.A1(_0736_),
    .A2(_0751_),
    .A3(_0898_),
    .B1(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__inv_2 _3831_ (.A(_0882_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_1 _3832_ (.A(_0902_),
    .B(_0885_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21o_1 _3833_ (.A1(_0887_),
    .A2(_0901_),
    .B1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__nor2_1 _3834_ (.A(_0871_),
    .B(_0874_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21o_1 _3835_ (.A1(_0877_),
    .A2(_0904_),
    .B1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nor2_1 _3836_ (.A(_0861_),
    .B(_0864_),
    .Y(_0907_));
 sky130_fd_sc_hd__a21o_1 _3837_ (.A1(_0866_),
    .A2(_0906_),
    .B1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__nor2_1 _3838_ (.A(_0850_),
    .B(_0853_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _3839_ (.A1(_0856_),
    .A2(_0908_),
    .B1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_1 _3840_ (.A(_0838_),
    .B(_0841_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21oi_1 _3841_ (.A1(_0845_),
    .A2(_0910_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2_1 _3842_ (.A(_0829_),
    .B(_0832_),
    .X(_0913_));
 sky130_fd_sc_hd__o21a_1 _3843_ (.A1(_0833_),
    .A2(_0912_),
    .B1(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__nand2_1 _3844_ (.A(_0776_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__and2_2 _3845_ (.A(_0773_),
    .B(_0774_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _3846_ (.A(_0401_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__clkbuf_4 _3847_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__inv_2 _3848_ (.A(_0832_),
    .Y(_0919_));
 sky130_fd_sc_hd__or2b_1 _3849_ (.A(_0746_),
    .B_N(_0750_),
    .X(_0920_));
 sky130_fd_sc_hd__and2b_1 _3850_ (.A_N(_0895_),
    .B(_0892_),
    .X(_0921_));
 sky130_fd_sc_hd__a31o_1 _3851_ (.A1(_0920_),
    .A2(_0896_),
    .A3(_0795_),
    .B1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2_1 _3852_ (.A(_0887_),
    .B(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a21boi_1 _3853_ (.A1(_0882_),
    .A2(_0885_),
    .B1_N(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__o21ba_1 _3854_ (.A1(_0876_),
    .A2(_0924_),
    .B1_N(_0875_),
    .X(_0925_));
 sky130_fd_sc_hd__or2b_1 _3855_ (.A(_0861_),
    .B_N(_0864_),
    .X(_0926_));
 sky130_fd_sc_hd__o21a_1 _3856_ (.A1(_0866_),
    .A2(_0925_),
    .B1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__and2b_1 _3857_ (.A_N(_0853_),
    .B(_0850_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_1 _3858_ (.A1(_0854_),
    .A2(_0927_),
    .B1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__o21ai_2 _3859_ (.A1(_0842_),
    .A2(_0929_),
    .B1(_0843_),
    .Y(_0930_));
 sky130_fd_sc_hd__o21a_1 _3860_ (.A1(_0829_),
    .A2(_0919_),
    .B1(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__a21o_1 _3861_ (.A1(_0829_),
    .A2(_0919_),
    .B1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__xnor2_1 _3862_ (.A(_0865_),
    .B(_0925_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _3863_ (.A(_0920_),
    .B(_0795_),
    .Y(_0934_));
 sky130_fd_sc_hd__xor2_2 _3864_ (.A(_0898_),
    .B(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__or2b_1 _3865_ (.A(_0812_),
    .B_N(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2_1 _3866_ (.A(_0887_),
    .B(_0922_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _3867_ (.A(_0923_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__and2b_1 _3868_ (.A_N(_0936_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_1 _3869_ (.A(_0877_),
    .B(_0924_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_0939_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_1 _3871_ (.A(_0933_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__xnor2_2 _3872_ (.A(_0856_),
    .B(_0927_),
    .Y(_0943_));
 sky130_fd_sc_hd__xnor2_1 _3873_ (.A(_0844_),
    .B(_0929_),
    .Y(_0944_));
 sky130_fd_sc_hd__and3_1 _3874_ (.A(_0942_),
    .B(_0943_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_2 _3875_ (.A(_0833_),
    .B(_0930_),
    .X(_0946_));
 sky130_fd_sc_hd__and3_1 _3876_ (.A(_0816_),
    .B(_0945_),
    .C(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _3877_ (.A(_0833_),
    .B(_0912_),
    .X(_0948_));
 sky130_fd_sc_hd__xnor2_1 _3878_ (.A(_0845_),
    .B(_0910_),
    .Y(_0949_));
 sky130_fd_sc_hd__xnor2_1 _3879_ (.A(_0856_),
    .B(_0908_),
    .Y(_0950_));
 sky130_fd_sc_hd__xnor2_1 _3880_ (.A(_0877_),
    .B(_0904_),
    .Y(_0951_));
 sky130_fd_sc_hd__xnor2_1 _3881_ (.A(_0887_),
    .B(_0901_),
    .Y(_0952_));
 sky130_fd_sc_hd__a21oi_1 _3882_ (.A1(_0736_),
    .A2(_0751_),
    .B1(_0899_),
    .Y(_0953_));
 sky130_fd_sc_hd__xnor2_1 _3883_ (.A(_0898_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__or2b_1 _3884_ (.A(_0770_),
    .B_N(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__or3_1 _3885_ (.A(_0951_),
    .B(_0952_),
    .C(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__xnor2_1 _3886_ (.A(_0866_),
    .B(_0906_),
    .Y(_0957_));
 sky130_fd_sc_hd__or3_1 _3887_ (.A(_0950_),
    .B(_0956_),
    .C(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__nor2_1 _3888_ (.A(_0949_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(_0948_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__o2bb2a_1 _3890_ (.A1_N(_0914_),
    .A2_N(_0960_),
    .B1(_0772_),
    .B2(_0776_),
    .X(_0961_));
 sky130_fd_sc_hd__a311o_1 _3891_ (.A1(_0918_),
    .A2(_0778_),
    .A3(_0932_),
    .B1(_0947_),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_1 _3892_ (.A(_0824_),
    .B(_0915_),
    .C(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a211o_1 _3893_ (.A1(_0619_),
    .A2(_0818_),
    .B1(_0823_),
    .C1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nor2_1 _3894_ (.A(_2900_),
    .B(_2910_),
    .Y(_0965_));
 sky130_fd_sc_hd__a311o_1 _3895_ (.A1(_0455_),
    .A2(_2928_),
    .A3(_0965_),
    .B1(_2912_),
    .C1(_2925_),
    .X(_0966_));
 sky130_fd_sc_hd__or2_2 _3896_ (.A(_0379_),
    .B(net148),
    .X(_0967_));
 sky130_fd_sc_hd__a211o_1 _3897_ (.A1(_2896_),
    .A2(_0386_),
    .B1(_0306_),
    .C1(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__o21ba_1 _3898_ (.A1(_0966_),
    .A2(_0968_),
    .B1_N(_0326_),
    .X(_0969_));
 sky130_fd_sc_hd__o22a_1 _3899_ (.A1(_2915_),
    .A2(_0304_),
    .B1(_2914_),
    .B2(_2934_),
    .X(_0970_));
 sky130_fd_sc_hd__nand2_1 _3900_ (.A(_2946_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__and2_1 _3901_ (.A(_2888_),
    .B(_2889_),
    .X(_0972_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(_0521_),
    .Y(_0973_));
 sky130_fd_sc_hd__a221o_1 _3903_ (.A1(_0359_),
    .A2(_0972_),
    .B1(_0364_),
    .B2(_0973_),
    .C1(_0296_),
    .X(_0974_));
 sky130_fd_sc_hd__or4_4 _3904_ (.A(_0320_),
    .B(_0969_),
    .C(_0971_),
    .D(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_1 _3905_ (.A(_0361_),
    .B(_0330_),
    .Y(_0976_));
 sky130_fd_sc_hd__a22oi_1 _3906_ (.A1(_2889_),
    .A2(_0965_),
    .B1(_0522_),
    .B2(_0359_),
    .Y(_0977_));
 sky130_fd_sc_hd__and4b_1 _3907_ (.A_N(_0306_),
    .B(_0526_),
    .C(_0976_),
    .D(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__and4b_1 _3908_ (.A_N(_0449_),
    .B(_0970_),
    .C(_0978_),
    .D(_2946_),
    .X(_0979_));
 sky130_fd_sc_hd__nor2_1 _3909_ (.A(_0297_),
    .B(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_0975_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _3911_ (.A(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _3912_ (.A(_2928_),
    .B(_0965_),
    .Y(_0983_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_2929_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__nor4_1 _3914_ (.A(_0308_),
    .B(_0326_),
    .C(_0739_),
    .D(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand2_4 _3915_ (.A(_0527_),
    .B(net237),
    .Y(_0986_));
 sky130_fd_sc_hd__nor3_1 _3916_ (.A(_0972_),
    .B(_0327_),
    .C(_0379_),
    .Y(_0987_));
 sky130_fd_sc_hd__o21a_1 _3917_ (.A1(_2922_),
    .A2(_2884_),
    .B1(_0471_),
    .X(_0988_));
 sky130_fd_sc_hd__a41o_1 _3918_ (.A1(_0983_),
    .A2(_0970_),
    .A3(_0987_),
    .A4(_0988_),
    .B1(_0296_),
    .X(_0989_));
 sky130_fd_sc_hd__a2111o_1 _3919_ (.A1(_2922_),
    .A2(_0386_),
    .B1(_0310_),
    .C1(_0322_),
    .D1(_0984_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_1 _3920_ (.A(_0295_),
    .B(_0967_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_4 _3921_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_4 _3922_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__or4_2 _3923_ (.A(_0449_),
    .B(_0971_),
    .C(_0990_),
    .D(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand3b_1 _3924_ (.A_N(_0986_),
    .B(_0989_),
    .C(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__inv_2 _3925_ (.A(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__or2_1 _3926_ (.A(_0989_),
    .B(_0994_),
    .X(_0997_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(_0986_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_2 _3928_ (.A(_0979_),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _3929_ (.A(_0975_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _3930_ (.A(_0998_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_0980_),
    .B(_0998_),
    .Y(_1002_));
 sky130_fd_sc_hd__nand2_1 _3932_ (.A(_1001_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__or2b_1 _3933_ (.A(_0994_),
    .B_N(_0989_),
    .X(_1004_));
 sky130_fd_sc_hd__or3_1 _3934_ (.A(_0975_),
    .B(_0979_),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o21ai_1 _3935_ (.A1(_0999_),
    .A2(_0997_),
    .B1(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_2 _3936_ (.A(_0975_),
    .Y(_1007_));
 sky130_fd_sc_hd__and2b_1 _3937_ (.A_N(_1004_),
    .B(_0986_),
    .X(_1008_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_0998_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__or3_1 _3939_ (.A(_1007_),
    .B(_0980_),
    .C(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__a21bo_1 _3940_ (.A1(_0986_),
    .A2(_1006_),
    .B1_N(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_2 _3941_ (.A(_0296_),
    .B(_2929_),
    .Y(_1012_));
 sky130_fd_sc_hd__and3_1 _3942_ (.A(_0372_),
    .B(_2932_),
    .C(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__o21a_1 _3943_ (.A1(\alu.Cin ),
    .A2(_1013_),
    .B1(_1012_),
    .X(_1014_));
 sky130_fd_sc_hd__a2111o_1 _3944_ (.A1(_0982_),
    .A2(_0996_),
    .B1(_1003_),
    .C1(_1011_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and3_1 _3945_ (.A(_0975_),
    .B(_0980_),
    .C(_1008_),
    .X(_1016_));
 sky130_fd_sc_hd__and2b_1 _3946_ (.A_N(_1013_),
    .B(_1014_),
    .X(_1017_));
 sky130_fd_sc_hd__nand2_1 _3947_ (.A(_1000_),
    .B(_1008_),
    .Y(_1018_));
 sky130_fd_sc_hd__or2_1 _3948_ (.A(_0970_),
    .B(_0986_),
    .X(_1019_));
 sky130_fd_sc_hd__nand3_1 _3949_ (.A(_0532_),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__nor3b_1 _3950_ (.A(_0981_),
    .B(_0997_),
    .C_N(_0986_),
    .Y(_1021_));
 sky130_fd_sc_hd__or4_1 _3951_ (.A(_1012_),
    .B(_0996_),
    .C(_1016_),
    .D(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__o41a_2 _3952_ (.A1(_1003_),
    .A2(_1011_),
    .A3(_1020_),
    .A4(_1022_),
    .B1(_2952_),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_1 _3953_ (.A(_0573_),
    .B(_1020_),
    .Y(_1024_));
 sky130_fd_sc_hd__o2bb2a_1 _3954_ (.A1_N(_1023_),
    .A2_N(_1024_),
    .B1(\alu.Cin ),
    .B2(_1021_),
    .X(_1025_));
 sky130_fd_sc_hd__a2111o_1 _3955_ (.A1(_0964_),
    .A2(_1015_),
    .B1(_1016_),
    .C1(_1017_),
    .D1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__nand2_2 _3956_ (.A(_2955_),
    .B(_0368_),
    .Y(_1027_));
 sky130_fd_sc_hd__o21a_1 _3957_ (.A1(\alu.Cin ),
    .A2(_1023_),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__a22o_1 _3958_ (.A1(_0370_),
    .A2(_0618_),
    .B1(_1026_),
    .B2(_1028_),
    .X(_0007_));
 sky130_fd_sc_hd__xor2_1 _3959_ (.A(_0711_),
    .B(_0712_),
    .X(_1029_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(_0512_),
    .Y(_1030_));
 sky130_fd_sc_hd__o21ai_1 _3961_ (.A1(_1030_),
    .A2(_1029_),
    .B1(_0772_),
    .Y(_1031_));
 sky130_fd_sc_hd__or2_2 _3962_ (.A(_0401_),
    .B(_0529_),
    .X(_1032_));
 sky130_fd_sc_hd__or2_1 _3963_ (.A(_1032_),
    .B(_0806_),
    .X(_1033_));
 sky130_fd_sc_hd__o211ai_1 _3964_ (.A1(_0757_),
    .A2(_1031_),
    .B1(_1033_),
    .C1(_0918_),
    .Y(_1034_));
 sky130_fd_sc_hd__or2_1 _3965_ (.A(_0780_),
    .B(_0711_),
    .X(_1035_));
 sky130_fd_sc_hd__a21oi_1 _3966_ (.A1(_0780_),
    .A2(_0711_),
    .B1(_0772_),
    .Y(_1036_));
 sky130_fd_sc_hd__o311a_1 _3967_ (.A1(_0573_),
    .A2(_0511_),
    .A3(_0401_),
    .B1(_1035_),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o22a_1 _3968_ (.A1(_0918_),
    .A2(_1029_),
    .B1(_1034_),
    .B2(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _3969_ (.A(_0571_),
    .B(_0711_),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _3970_ (.A(_0709_),
    .Y(_1040_));
 sky130_fd_sc_hd__or2b_1 _3971_ (.A(_0447_),
    .B_N(_0585_),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_1 _3972_ (.A(_0596_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__o22a_1 _3973_ (.A1(_0596_),
    .A2(_0600_),
    .B1(_0604_),
    .B2(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__o221ai_1 _3974_ (.A1(_0597_),
    .A2(_0608_),
    .B1(_1042_),
    .B2(_0610_),
    .C1(_0605_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_0532_),
    .B(_0546_),
    .Y(_1045_));
 sky130_fd_sc_hd__a221o_1 _3976_ (.A1(_0819_),
    .A2(_0822_),
    .B1(_1044_),
    .B2(_0546_),
    .C1(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__a211o_1 _3977_ (.A1(_0559_),
    .A2(_1040_),
    .B1(_1043_),
    .C1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__a211o_4 _3978_ (.A1(_0518_),
    .A2(_1038_),
    .B1(_1039_),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__clkbuf_4 _3979_ (.A(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__buf_4 _3980_ (.A(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__inv_2 _3981_ (.A(_1021_),
    .Y(_1051_));
 sky130_fd_sc_hd__o2111a_1 _3982_ (.A1(_0372_),
    .A2(_0371_),
    .B1(_0773_),
    .C1(_1019_),
    .D1(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__nor2_1 _3983_ (.A(_0395_),
    .B(_1019_),
    .Y(_1053_));
 sky130_fd_sc_hd__o2bb2a_1 _3984_ (.A1_N(_1023_),
    .A2_N(_1052_),
    .B1(_1053_),
    .B2(\cu.alu_f[1] ),
    .X(_1054_));
 sky130_fd_sc_hd__o21ai_1 _3985_ (.A1(_0455_),
    .A2(_1001_),
    .B1(_1002_),
    .Y(_1055_));
 sky130_fd_sc_hd__o221a_1 _3986_ (.A1(\cu.alu_f[1] ),
    .A2(_1023_),
    .B1(_1054_),
    .B2(_1055_),
    .C1(_1027_),
    .X(_1056_));
 sky130_fd_sc_hd__a21o_1 _3987_ (.A1(_0370_),
    .A2(_1050_),
    .B1(_1056_),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _3988_ (.A(_0600_),
    .Y(_1057_));
 sky130_fd_sc_hd__and3_1 _3989_ (.A(_0447_),
    .B(_0585_),
    .C(_0596_),
    .X(_1058_));
 sky130_fd_sc_hd__o2bb2a_1 _3990_ (.A1_N(_0585_),
    .A2_N(_1057_),
    .B1(_0604_),
    .B2(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__a221o_1 _3991_ (.A1(_0559_),
    .A2(_0693_),
    .B1(_0822_),
    .B2(_0546_),
    .C1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__a21oi_1 _3992_ (.A1(_0760_),
    .A2(_0771_),
    .B1(_0776_),
    .Y(_1061_));
 sky130_fd_sc_hd__o21bai_1 _3993_ (.A1(_0757_),
    .A2(_0759_),
    .B1_N(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a21oi_1 _3994_ (.A1(_0815_),
    .A2(_0806_),
    .B1(_0775_),
    .Y(_1063_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(_1033_),
    .A1(_1063_),
    .S(_0805_),
    .X(_1064_));
 sky130_fd_sc_hd__a2bb2o_1 _3996_ (.A1_N(_0918_),
    .A2_N(_0759_),
    .B1(_1062_),
    .B2(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_0619_),
    .B(_0824_),
    .Y(_1066_));
 sky130_fd_sc_hd__o22a_1 _3998_ (.A1(_0571_),
    .A2(_0758_),
    .B1(_1065_),
    .B2(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__o221a_1 _3999_ (.A1(_0585_),
    .A2(_0608_),
    .B1(_1058_),
    .B2(_0610_),
    .C1(_0605_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(_0532_),
    .A1(_1068_),
    .S(_1040_),
    .X(_1069_));
 sky130_fd_sc_hd__nand3b_4 _4001_ (.A_N(_1060_),
    .B(_1067_),
    .C(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__buf_4 _4002_ (.A(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_8 _4003_ (.A(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__and3b_1 _4004_ (.A_N(_0760_),
    .B(_0763_),
    .C(_0771_),
    .X(_1073_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(_0763_),
    .B(_1061_),
    .Y(_1074_));
 sky130_fd_sc_hd__nor2_1 _4006_ (.A(_0807_),
    .B(_0809_),
    .Y(_1075_));
 sky130_fd_sc_hd__a21o_1 _4007_ (.A1(_0816_),
    .A2(_0807_),
    .B1(_0775_),
    .X(_1076_));
 sky130_fd_sc_hd__a22o_1 _4008_ (.A1(_0816_),
    .A2(_1075_),
    .B1(_1076_),
    .B2(_0809_),
    .X(_1077_));
 sky130_fd_sc_hd__o31a_1 _4009_ (.A1(_1073_),
    .A2(_1074_),
    .A3(_1077_),
    .B1(_0518_),
    .X(_1078_));
 sky130_fd_sc_hd__nor2_1 _4010_ (.A(_0571_),
    .B(_0762_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_1 _4011_ (.A(_0597_),
    .B(_1041_),
    .Y(_1080_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(_0532_),
    .B(_0693_),
    .Y(_1081_));
 sky130_fd_sc_hd__a221o_1 _4013_ (.A1(_0604_),
    .A2(_0700_),
    .B1(_1080_),
    .B2(_0600_),
    .C1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__or2_1 _4014_ (.A(_0600_),
    .B(_0604_),
    .X(_1083_));
 sky130_fd_sc_hd__a2bb2o_1 _4015_ (.A1_N(_0610_),
    .A2_N(_1080_),
    .B1(_0700_),
    .B2(_0607_),
    .X(_1084_));
 sky130_fd_sc_hd__o21a_1 _4016_ (.A1(_1083_),
    .A2(_1084_),
    .B1(_0693_),
    .X(_1085_));
 sky130_fd_sc_hd__a221o_1 _4017_ (.A1(_0559_),
    .A2(_0680_),
    .B1(_0822_),
    .B2(_1040_),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__or4_4 _4018_ (.A(_1078_),
    .B(_1079_),
    .C(_1082_),
    .D(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__xnor2_1 _4019_ (.A(_1070_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_0769_),
    .B(_0772_),
    .Y(_1089_));
 sky130_fd_sc_hd__o2bb2a_1 _4021_ (.A1_N(_0775_),
    .A2_N(_0800_),
    .B1(_1089_),
    .B2(_0767_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_1 _4022_ (.A(_0800_),
    .B(_0811_),
    .Y(_1091_));
 sky130_fd_sc_hd__and2_1 _4023_ (.A(_0800_),
    .B(_0811_),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_1 _4024_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(_0767_),
    .B(_0771_),
    .Y(_1094_));
 sky130_fd_sc_hd__and2_1 _4026_ (.A(_0918_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__o22a_1 _4027_ (.A1(_1032_),
    .A2(_1093_),
    .B1(_1095_),
    .B2(_0769_),
    .X(_1096_));
 sky130_fd_sc_hd__a21oi_1 _4028_ (.A1(_1090_),
    .A2(_1096_),
    .B1(_1066_),
    .Y(_1097_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(_0447_),
    .B(_0585_),
    .X(_1098_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__a21oi_1 _4031_ (.A1(_0596_),
    .A2(_1099_),
    .B1(_0610_),
    .Y(_1100_));
 sky130_fd_sc_hd__a211o_1 _4032_ (.A1(_0607_),
    .A2(_0728_),
    .B1(_1083_),
    .C1(_0553_),
    .X(_1101_));
 sky130_fd_sc_hd__a32o_1 _4033_ (.A1(_0596_),
    .A2(_0600_),
    .A3(_1099_),
    .B1(_0728_),
    .B2(_0604_),
    .X(_1102_));
 sky130_fd_sc_hd__o22a_1 _4034_ (.A1(_1100_),
    .A2(_1101_),
    .B1(_1102_),
    .B2(_0567_),
    .X(_1103_));
 sky130_fd_sc_hd__o2bb2a_1 _4035_ (.A1_N(\alu.Cin ),
    .A2_N(_0555_),
    .B1(_0557_),
    .B2(net142),
    .X(_1104_));
 sky130_fd_sc_hd__o2bb2a_1 _4036_ (.A1_N(_0822_),
    .A2_N(_0631_),
    .B1(_0567_),
    .B2(_0532_),
    .X(_1105_));
 sky130_fd_sc_hd__o211a_1 _4037_ (.A1(_0571_),
    .A2(_0732_),
    .B1(_1104_),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__or3b_1 _4038_ (.A(_1097_),
    .B(_1103_),
    .C_N(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__buf_4 _4039_ (.A(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nand2_1 _4040_ (.A(_0607_),
    .B(_0642_),
    .Y(_1109_));
 sky130_fd_sc_hd__or2_1 _4041_ (.A(_0585_),
    .B(_0610_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_4 _4042_ (.A(_0447_),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_1111_),
    .B(_0596_),
    .Y(_1112_));
 sky130_fd_sc_hd__o2bb2a_1 _4044_ (.A1_N(_0610_),
    .A2_N(_1109_),
    .B1(_1110_),
    .B2(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__o21a_1 _4045_ (.A1(_1083_),
    .A2(_1113_),
    .B1(_0631_),
    .X(_1114_));
 sky130_fd_sc_hd__a2bb2o_1 _4046_ (.A1_N(_0532_),
    .A2_N(_0631_),
    .B1(_0567_),
    .B2(_0559_),
    .X(_1115_));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(_0585_),
    .B(_1057_),
    .X(_1116_));
 sky130_fd_sc_hd__nor2_1 _4048_ (.A(_1112_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a221o_1 _4049_ (.A1(_0604_),
    .A2(_0642_),
    .B1(_0662_),
    .B2(_0822_),
    .C1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__or2_1 _4050_ (.A(_0756_),
    .B(_0766_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_1 _4051_ (.A(_0803_),
    .B(_0810_),
    .Y(_1120_));
 sky130_fd_sc_hd__o21ai_1 _4052_ (.A1(_1032_),
    .A2(_1120_),
    .B1(_0916_),
    .Y(_1121_));
 sky130_fd_sc_hd__o2bb2a_1 _4053_ (.A1_N(_0801_),
    .A2_N(_1121_),
    .B1(_0811_),
    .B2(_1032_),
    .X(_1122_));
 sky130_fd_sc_hd__o221a_1 _4054_ (.A1(_1119_),
    .A2(_1094_),
    .B1(_1095_),
    .B2(_0753_),
    .C1(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__o22a_1 _4055_ (.A1(_0571_),
    .A2(_0643_),
    .B1(_1123_),
    .B2(_1066_),
    .X(_1124_));
 sky130_fd_sc_hd__or4b_4 _4056_ (.A(_1114_),
    .B(_1115_),
    .C(_1118_),
    .D_N(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_1108_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__and2_1 _4058_ (.A(_1108_),
    .B(_1125_),
    .X(_1127_));
 sky130_fd_sc_hd__nor2_1 _4059_ (.A(_1126_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__and2_1 _4060_ (.A(_0803_),
    .B(_0810_),
    .X(_1129_));
 sky130_fd_sc_hd__o21a_1 _4061_ (.A1(_1120_),
    .A2(_1129_),
    .B1(_0816_),
    .X(_1130_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(_0756_),
    .B(_0766_),
    .Y(_1131_));
 sky130_fd_sc_hd__a2bb2o_1 _4063_ (.A1_N(_0917_),
    .A2_N(_0756_),
    .B1(_0803_),
    .B2(_0775_),
    .X(_1132_));
 sky130_fd_sc_hd__a31o_1 _4064_ (.A1(_1119_),
    .A2(_0772_),
    .A3(_1131_),
    .B1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__o21a_1 _4065_ (.A1(_1130_),
    .A2(_1133_),
    .B1(_0518_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(_0596_),
    .B(_1098_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _4067_ (.A(_0600_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__a21oi_1 _4068_ (.A1(_0718_),
    .A2(_1136_),
    .B1(_0605_),
    .Y(_1137_));
 sky130_fd_sc_hd__a2bb2o_1 _4069_ (.A1_N(_0610_),
    .A2_N(_1135_),
    .B1(_0651_),
    .B2(_0607_),
    .X(_1138_));
 sky130_fd_sc_hd__a2bb2o_1 _4070_ (.A1_N(_0532_),
    .A2_N(_0662_),
    .B1(_0680_),
    .B2(_0822_),
    .X(_1139_));
 sky130_fd_sc_hd__a221o_1 _4071_ (.A1(_0559_),
    .A2(_0631_),
    .B1(_0662_),
    .B2(_1138_),
    .C1(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(_0571_),
    .B(_0663_),
    .Y(_1141_));
 sky130_fd_sc_hd__or4_1 _4073_ (.A(_1134_),
    .B(_1137_),
    .C(_1140_),
    .D(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__buf_4 _4074_ (.A(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _4075_ (.A(_0764_),
    .B(_0765_),
    .X(_1144_));
 sky130_fd_sc_hd__o21ai_1 _4076_ (.A1(_0807_),
    .A2(_0809_),
    .B1(_0804_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand2_1 _4077_ (.A(_0810_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__a221o_1 _4078_ (.A1(_0775_),
    .A2(_0804_),
    .B1(_1146_),
    .B2(_0816_),
    .C1(_0776_),
    .X(_1147_));
 sky130_fd_sc_hd__a31o_1 _4079_ (.A1(_0766_),
    .A2(_0772_),
    .A3(_1144_),
    .B1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o211a_1 _4080_ (.A1(_0918_),
    .A2(_0765_),
    .B1(_1148_),
    .C1(_0518_),
    .X(_1149_));
 sky130_fd_sc_hd__nor2_1 _4081_ (.A(_0571_),
    .B(_0683_),
    .Y(_1150_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(_0559_),
    .A2(_0662_),
    .B1(_0822_),
    .B2(_0693_),
    .X(_1151_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_1111_),
    .B(_0597_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _4084_ (.A(_0607_),
    .B(_0670_),
    .Y(_1153_));
 sky130_fd_sc_hd__a2bb2o_1 _4085_ (.A1_N(_1152_),
    .A2_N(_1110_),
    .B1(_1153_),
    .B2(_0610_),
    .X(_1154_));
 sky130_fd_sc_hd__nor2_1 _4086_ (.A(_1152_),
    .B(_1116_),
    .Y(_1155_));
 sky130_fd_sc_hd__a211oi_1 _4087_ (.A1(_0604_),
    .A2(_0670_),
    .B1(_0680_),
    .C1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__a32o_1 _4088_ (.A1(_0605_),
    .A2(_0680_),
    .A3(_1154_),
    .B1(_1156_),
    .B2(_0532_),
    .X(_1157_));
 sky130_fd_sc_hd__or4b_1 _4089_ (.A(_1149_),
    .B(_1150_),
    .C(_1151_),
    .D_N(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__buf_4 _4090_ (.A(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__xor2_1 _4091_ (.A(_1143_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__xor2_1 _4092_ (.A(_0616_),
    .B(_1048_),
    .X(_1161_));
 sky130_fd_sc_hd__xnor2_1 _4093_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__xnor2_1 _4094_ (.A(_1128_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__inv_2 _4095_ (.A(_0820_),
    .Y(_1164_));
 sky130_fd_sc_hd__o211ai_1 _4096_ (.A1(_0520_),
    .A2(_1164_),
    .B1(_0613_),
    .C1(_0552_),
    .Y(_1165_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(_1088_),
    .B(_1163_),
    .Y(_1166_));
 sky130_fd_sc_hd__o221a_1 _4098_ (.A1(_1088_),
    .A2(_1163_),
    .B1(_1165_),
    .B2(_0607_),
    .C1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__xnor2_1 _4099_ (.A(_0567_),
    .B(_1108_),
    .Y(_1168_));
 sky130_fd_sc_hd__xor2_1 _4100_ (.A(_0547_),
    .B(_0732_),
    .X(_1169_));
 sky130_fd_sc_hd__xor2_1 _4101_ (.A(_0945_),
    .B(_0946_),
    .X(_1170_));
 sky130_fd_sc_hd__o221a_1 _4102_ (.A1(_0916_),
    .A2(_0946_),
    .B1(_1170_),
    .B2(_1032_),
    .C1(_0918_),
    .X(_1171_));
 sky130_fd_sc_hd__o21a_1 _4103_ (.A1(_0948_),
    .A2(_0959_),
    .B1(_0772_),
    .X(_1172_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_0960_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__a2bb2o_2 _4105_ (.A1_N(_0918_),
    .A2_N(_0948_),
    .B1(_1171_),
    .B2(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__xnor2_1 _4106_ (.A(_0829_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__o21ai_1 _4107_ (.A1(_0548_),
    .A2(_0833_),
    .B1(_0824_),
    .Y(_1176_));
 sky130_fd_sc_hd__a211o_1 _4108_ (.A1(_0548_),
    .A2(_0833_),
    .B1(_1175_),
    .C1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__o31ai_1 _4109_ (.A1(_0395_),
    .A2(_1168_),
    .A3(_1169_),
    .B1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__o21a_1 _4110_ (.A1(\cu.alu_f[2] ),
    .A2(_1013_),
    .B1(_1012_),
    .X(_1179_));
 sky130_fd_sc_hd__a21oi_1 _4111_ (.A1(_1018_),
    .A2(_1019_),
    .B1(_0395_),
    .Y(_1180_));
 sky130_fd_sc_hd__or4b_2 _4112_ (.A(_0996_),
    .B(_1003_),
    .C(_1180_),
    .D_N(_1010_),
    .X(_1181_));
 sky130_fd_sc_hd__o221a_1 _4113_ (.A1(_1167_),
    .A2(_1178_),
    .B1(_1179_),
    .B2(_1181_),
    .C1(_1023_),
    .X(_1182_));
 sky130_fd_sc_hd__o21ai_2 _4114_ (.A1(_1013_),
    .A2(_1181_),
    .B1(_1023_),
    .Y(_1183_));
 sky130_fd_sc_hd__a21o_1 _4115_ (.A1(\cu.alu_f[2] ),
    .A2(_1183_),
    .B1(_0370_),
    .X(_1184_));
 sky130_fd_sc_hd__o22a_1 _4116_ (.A1(_1027_),
    .A2(_1072_),
    .B1(_1182_),
    .B2(_1184_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_2 _4117_ (.A(_2950_),
    .B(_2951_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_4 _4118_ (.A(_1087_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_8 _4119_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a22o_1 _4120_ (.A1(net207),
    .A2(_1185_),
    .B1(_0370_),
    .B2(_1187_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_4 _4121_ (.A(_1159_),
    .X(_1188_));
 sky130_fd_sc_hd__buf_4 _4122_ (.A(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__a22o_1 _4123_ (.A1(net208),
    .A2(_1185_),
    .B1(_0370_),
    .B2(_1189_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _4124_ (.A(_1143_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_8 _4125_ (.A(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__a22o_1 _4126_ (.A1(net209),
    .A2(_1185_),
    .B1(_0370_),
    .B2(_1191_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_4 _4127_ (.A(_1125_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_8 _4128_ (.A(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__a21oi_1 _4129_ (.A1(_0942_),
    .A2(_0943_),
    .B1(_0944_),
    .Y(_1194_));
 sky130_fd_sc_hd__nor2_1 _4130_ (.A(_0945_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__o221a_1 _4131_ (.A1(_0916_),
    .A2(_0944_),
    .B1(_1195_),
    .B2(_1032_),
    .C1(_0918_),
    .X(_1196_));
 sky130_fd_sc_hd__a21o_1 _4132_ (.A1(_0949_),
    .A2(_0958_),
    .B1(_0778_),
    .X(_1197_));
 sky130_fd_sc_hd__or2_1 _4133_ (.A(_0959_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _4134_ (.A1(_0776_),
    .A2(_0949_),
    .B1(_1196_),
    .B2(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__nand2_1 _4135_ (.A(_0942_),
    .B(_0943_),
    .Y(_1200_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_0942_),
    .B(_0943_),
    .X(_1201_));
 sky130_fd_sc_hd__a21o_1 _4137_ (.A1(_1200_),
    .A2(_1201_),
    .B1(_1032_),
    .X(_1202_));
 sky130_fd_sc_hd__nor2_1 _4138_ (.A(_0956_),
    .B(_0957_),
    .Y(_1203_));
 sky130_fd_sc_hd__or2_1 _4139_ (.A(_1203_),
    .B(_0778_),
    .X(_1204_));
 sky130_fd_sc_hd__and2_1 _4140_ (.A(_0918_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__nand3_1 _4141_ (.A(_0950_),
    .B(_1203_),
    .C(_0772_),
    .Y(_1206_));
 sky130_fd_sc_hd__o221a_1 _4142_ (.A1(_0916_),
    .A2(_0943_),
    .B1(_1205_),
    .B2(_0950_),
    .C1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__a21oi_4 _4143_ (.A1(_1202_),
    .A2(_1207_),
    .B1(_0517_),
    .Y(_1208_));
 sky130_fd_sc_hd__a21o_1 _4144_ (.A1(_0816_),
    .A2(_0941_),
    .B1(_0775_),
    .X(_1209_));
 sky130_fd_sc_hd__a22oi_1 _4145_ (.A1(_0816_),
    .A2(_0942_),
    .B1(_1209_),
    .B2(_0933_),
    .Y(_1210_));
 sky130_fd_sc_hd__o221a_1 _4146_ (.A1(_0956_),
    .A2(_1204_),
    .B1(_1205_),
    .B2(_0957_),
    .C1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__nor2_4 _4147_ (.A(_0517_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__nor2_1 _4148_ (.A(_0952_),
    .B(_0955_),
    .Y(_1213_));
 sky130_fd_sc_hd__or2_1 _4149_ (.A(_1213_),
    .B(_0778_),
    .X(_1214_));
 sky130_fd_sc_hd__and2_1 _4150_ (.A(_0917_),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nor2_1 _4151_ (.A(_0951_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__or2_1 _4152_ (.A(_0939_),
    .B(_0940_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2_1 _4153_ (.A(_0941_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__a2bb2o_1 _4154_ (.A1_N(_0916_),
    .A2_N(_0940_),
    .B1(_1218_),
    .B2(_0816_),
    .X(_1219_));
 sky130_fd_sc_hd__a31o_1 _4155_ (.A1(_0951_),
    .A2(_1213_),
    .A3(_0772_),
    .B1(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__o21a_4 _4156_ (.A1(_1216_),
    .A2(_1220_),
    .B1(_0824_),
    .X(_1221_));
 sky130_fd_sc_hd__a21oi_1 _4157_ (.A1(_0815_),
    .A2(_0936_),
    .B1(_0775_),
    .Y(_1222_));
 sky130_fd_sc_hd__o2bb2a_1 _4158_ (.A1_N(_0816_),
    .A2_N(_0939_),
    .B1(_1222_),
    .B2(_0938_),
    .X(_1223_));
 sky130_fd_sc_hd__o221a_1 _4159_ (.A1(_0955_),
    .A2(_1214_),
    .B1(_1215_),
    .B2(_0952_),
    .C1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__nor2_4 _4160_ (.A(_0517_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__xnor2_1 _4161_ (.A(_0935_),
    .B(_0812_),
    .Y(_1226_));
 sky130_fd_sc_hd__o32a_1 _4162_ (.A1(_0770_),
    .A2(_0954_),
    .A3(_0778_),
    .B1(_0935_),
    .B2(_0916_),
    .X(_1227_));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(_0954_),
    .B(_0777_),
    .Y(_1228_));
 sky130_fd_sc_hd__o211a_1 _4164_ (.A1(_1032_),
    .A2(_1226_),
    .B1(_1227_),
    .C1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__or4b_1 _4165_ (.A(_0517_),
    .B(_0818_),
    .C(_1225_),
    .D_N(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__nor4_1 _4166_ (.A(_1208_),
    .B(_1212_),
    .C(_1221_),
    .D(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__clkbuf_8 _4167_ (.A(_2931_),
    .X(_1232_));
 sky130_fd_sc_hd__nor2_2 _4168_ (.A(_1232_),
    .B(_0371_),
    .Y(_1233_));
 sky130_fd_sc_hd__a21oi_1 _4169_ (.A1(_0387_),
    .A2(_1233_),
    .B1(_0824_),
    .Y(_1234_));
 sky130_fd_sc_hd__a31o_1 _4170_ (.A1(_1174_),
    .A2(_1199_),
    .A3(_1231_),
    .B1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__or4_1 _4171_ (.A(_0616_),
    .B(_1048_),
    .C(_1070_),
    .D(_1087_),
    .X(_1236_));
 sky130_fd_sc_hd__nor3_1 _4172_ (.A(_1143_),
    .B(_1159_),
    .C(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(_0829_),
    .A1(_0838_),
    .S(_1111_),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(_0850_),
    .A1(_0861_),
    .S(_1111_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(_1238_),
    .A1(_1239_),
    .S(_0597_),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(_0871_),
    .A1(_0902_),
    .S(_1111_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(_0892_),
    .A1(_0746_),
    .S(_1111_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(_1241_),
    .A1(_1242_),
    .S(_0597_),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(_1240_),
    .A1(_1243_),
    .S(_0585_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(_0567_),
    .A1(_0631_),
    .S(_1111_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(_0662_),
    .A1(_0680_),
    .S(_1111_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(_1245_),
    .A1(_1246_),
    .S(_0597_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(_0546_),
    .A1(_0819_),
    .S(_1111_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(_0693_),
    .A1(_1040_),
    .S(_1111_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(_1248_),
    .A1(_1249_),
    .S(_0596_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(_1247_),
    .A1(_1250_),
    .S(_0585_),
    .X(_1251_));
 sky130_fd_sc_hd__nor2_1 _4187_ (.A(_0700_),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21o_1 _4188_ (.A1(_0700_),
    .A2(_1244_),
    .B1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__and3_1 _4189_ (.A(_0387_),
    .B(_1233_),
    .C(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a31o_1 _4190_ (.A1(_1126_),
    .A2(_1235_),
    .A3(_1237_),
    .B1(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__o21a_1 _4191_ (.A1(_1233_),
    .A2(_1181_),
    .B1(_1023_),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(\cu.alu_f[6] ),
    .A1(_1255_),
    .S(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(_1193_),
    .A1(_1257_),
    .S(_1027_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _4194_ (.A(_1258_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_4 _4195_ (.A(_1108_),
    .X(_1259_));
 sky130_fd_sc_hd__buf_4 _4196_ (.A(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(_1183_),
    .Y(_1261_));
 sky130_fd_sc_hd__nor2_4 _4198_ (.A(_0517_),
    .B(_1174_),
    .Y(_1262_));
 sky130_fd_sc_hd__a22o_1 _4199_ (.A1(_0517_),
    .A2(_1259_),
    .B1(_1262_),
    .B2(_1027_),
    .X(_1263_));
 sky130_fd_sc_hd__and3_1 _4200_ (.A(\cu.alu_f[7] ),
    .B(_1027_),
    .C(_1183_),
    .X(_1264_));
 sky130_fd_sc_hd__a221o_1 _4201_ (.A1(_0370_),
    .A2(_1260_),
    .B1(_1261_),
    .B2(_1263_),
    .C1(_1264_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _4202_ (.A(_2880_),
    .B(_0403_),
    .C(_0471_),
    .X(_1265_));
 sky130_fd_sc_hd__o211a_1 _4203_ (.A1(_0322_),
    .A2(_1265_),
    .B1(_2914_),
    .C1(_2947_),
    .X(_1266_));
 sky130_fd_sc_hd__buf_2 _4204_ (.A(\cu.id.state[2] ),
    .X(_1267_));
 sky130_fd_sc_hd__and3b_2 _4205_ (.A_N(\cu.id.state[1] ),
    .B(\cu.id.state[0] ),
    .C(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__or3b_1 _4206_ (.A(_0294_),
    .B(_1266_),
    .C_N(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__buf_2 _4207_ (.A(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__o211ai_2 _4208_ (.A1(_2886_),
    .A2(_2947_),
    .B1(_0339_),
    .C1(_2914_),
    .Y(_1271_));
 sky130_fd_sc_hd__a31o_1 _4209_ (.A1(_2880_),
    .A2(_0334_),
    .A3(_0403_),
    .B1(_0293_),
    .X(_1272_));
 sky130_fd_sc_hd__inv_2 _4210_ (.A(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__or2_1 _4211_ (.A(_0359_),
    .B(_2947_),
    .X(_1274_));
 sky130_fd_sc_hd__a21o_1 _4212_ (.A1(_0334_),
    .A2(_1265_),
    .B1(_0293_),
    .X(_1275_));
 sky130_fd_sc_hd__a31o_1 _4213_ (.A1(_2914_),
    .A2(_0339_),
    .A3(_1274_),
    .B1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a31o_2 _4214_ (.A1(_2914_),
    .A2(_2947_),
    .A3(_0339_),
    .B1(_1275_),
    .X(_1277_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(_0471_),
    .Y(_1278_));
 sky130_fd_sc_hd__a2111oi_1 _4216_ (.A1(_1271_),
    .A2(_1273_),
    .B1(_1276_),
    .C1(_1277_),
    .D1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__buf_2 _4217_ (.A(net144),
    .X(_1280_));
 sky130_fd_sc_hd__and3_2 _4218_ (.A(_1271_),
    .B(_1273_),
    .C(_1276_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_4 _4219_ (.A(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__and3b_2 _4220_ (.A_N(_1276_),
    .B(_1271_),
    .C(_1273_),
    .X(_1283_));
 sky130_fd_sc_hd__buf_2 _4221_ (.A(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__nor2_4 _4222_ (.A(_0295_),
    .B(_0471_),
    .Y(_1285_));
 sky130_fd_sc_hd__clkbuf_4 _4223_ (.A(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a22o_1 _4224_ (.A1(\cu.reg_file.reg_a[0] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[0] ),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _4225_ (.A1(\cu.reg_file.reg_e[0] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[0] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a21oi_1 _4226_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_1280_),
    .B1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__nor2_1 _4227_ (.A(_1270_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(_2907_),
    .B(_2935_),
    .Y(_1291_));
 sky130_fd_sc_hd__and3_1 _4229_ (.A(_2954_),
    .B(_1291_),
    .C(_1268_),
    .X(_1292_));
 sky130_fd_sc_hd__buf_2 _4230_ (.A(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__buf_2 _4231_ (.A(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__inv_2 _4232_ (.A(_1270_),
    .Y(_1295_));
 sky130_fd_sc_hd__nor2_2 _4233_ (.A(_1295_),
    .B(_1293_),
    .Y(_1296_));
 sky130_fd_sc_hd__buf_2 _4234_ (.A(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_4 _4235_ (.A(\cu.pc.pc_o[0] ),
    .X(_1298_));
 sky130_fd_sc_hd__buf_2 _4236_ (.A(\cu.id.state[0] ),
    .X(_1299_));
 sky130_fd_sc_hd__buf_2 _4237_ (.A(\cu.id.state[1] ),
    .X(_1300_));
 sky130_fd_sc_hd__and2b_1 _4238_ (.A_N(_1299_),
    .B(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__inv_2 _4239_ (.A(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__nor2_2 _4240_ (.A(_2950_),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__clkbuf_8 _4241_ (.A(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__a221o_1 _4242_ (.A1(_0344_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(_1298_),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__a211oi_1 _4243_ (.A1(_0359_),
    .A2(_0319_),
    .B1(_0334_),
    .C1(_2917_),
    .Y(_1306_));
 sky130_fd_sc_hd__a211o_2 _4244_ (.A1(_0334_),
    .A2(_0403_),
    .B1(_1306_),
    .C1(_0295_),
    .X(_1307_));
 sky130_fd_sc_hd__o31a_1 _4245_ (.A1(_2912_),
    .A2(_0361_),
    .A3(_0967_),
    .B1(_0334_),
    .X(_1308_));
 sky130_fd_sc_hd__a2111o_2 _4246_ (.A1(_2886_),
    .A2(_0319_),
    .B1(_1308_),
    .C1(_0295_),
    .D1(_2917_),
    .X(_1309_));
 sky130_fd_sc_hd__and3b_2 _4247_ (.A_N(_0992_),
    .B(_1307_),
    .C(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_4 _4248_ (.A(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_2 _4249_ (.A(_1307_),
    .B(_1309_),
    .Y(_1312_));
 sky130_fd_sc_hd__buf_2 _4250_ (.A(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__nor2b_2 _4251_ (.A(_1307_),
    .B_N(_1309_),
    .Y(_1314_));
 sky130_fd_sc_hd__buf_2 _4252_ (.A(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__or4b_2 _4253_ (.A(_2896_),
    .B(_2904_),
    .C(_2934_),
    .D_N(_2922_),
    .X(_1316_));
 sky130_fd_sc_hd__inv_2 _4254_ (.A(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or4_2 _4255_ (.A(_0295_),
    .B(_2917_),
    .C(_0319_),
    .D(_1308_),
    .X(_1318_));
 sky130_fd_sc_hd__nor2_4 _4256_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__clkbuf_4 _4257_ (.A(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_2 _4258_ (.A(_1267_),
    .B(_1301_),
    .Y(_1321_));
 sky130_fd_sc_hd__clkbuf_4 _4259_ (.A(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a31o_1 _4260_ (.A1(_0344_),
    .A2(_2954_),
    .A3(_1317_),
    .B1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a221o_1 _4261_ (.A1(\cu.reg_file.reg_sp[0] ),
    .A2(_0993_),
    .B1(_1320_),
    .B2(_1298_),
    .C1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__a221o_1 _4262_ (.A1(\cu.reg_file.reg_e[0] ),
    .A2(_1313_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_l[0] ),
    .C1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__a21oi_2 _4263_ (.A1(\cu.reg_file.reg_c[0] ),
    .A2(_1311_),
    .B1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__o21bai_4 _4264_ (.A1(_1290_),
    .A2(_1305_),
    .B1_N(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__inv_2 _4265_ (.A(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__and2_1 _4266_ (.A(\mc.rw.state[2] ),
    .B(_2701_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_4 _4267_ (.A(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_4 _4268_ (.A(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__or2_1 _4269_ (.A(_2698_),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_2 _4270_ (.A(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_4 _4271_ (.A(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_4 _4272_ (.A(_1327_),
    .X(_1335_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(\mc.rw.state[2] ),
    .B(_2708_),
    .Y(_1336_));
 sky130_fd_sc_hd__or4_1 _4274_ (.A(_2703_),
    .B(_2709_),
    .C(_1335_),
    .D(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__o21a_1 _4275_ (.A1(_1328_),
    .A2(_1334_),
    .B1(_1337_),
    .X(net35));
 sky130_fd_sc_hd__nor2_2 _4276_ (.A(_0295_),
    .B(_1316_),
    .Y(_1338_));
 sky130_fd_sc_hd__clkbuf_4 _4277_ (.A(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__a221o_1 _4278_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(_0341_),
    .C1(_1322_),
    .X(_1340_));
 sky130_fd_sc_hd__a221o_1 _4279_ (.A1(\cu.pc.pc_o[1] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[1] ),
    .C1(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__a21oi_1 _4280_ (.A1(\cu.reg_file.reg_l[1] ),
    .A2(_1315_),
    .B1(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _4281_ (.A(\cu.reg_file.reg_c[1] ),
    .B(_1311_),
    .Y(_1343_));
 sky130_fd_sc_hd__a22o_1 _4282_ (.A1(\cu.reg_file.reg_a[1] ),
    .A2(_1277_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[1] ),
    .X(_1344_));
 sky130_fd_sc_hd__a221o_1 _4283_ (.A1(\cu.reg_file.reg_e[1] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[1] ),
    .C1(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__a21o_1 _4284_ (.A1(\cu.reg_file.reg_c[1] ),
    .A2(_1280_),
    .B1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a221o_1 _4285_ (.A1(_0341_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[1] ),
    .C1(_1303_),
    .X(_1347_));
 sky130_fd_sc_hd__a21oi_1 _4286_ (.A1(_1295_),
    .A2(_1346_),
    .B1(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__a21oi_4 _4287_ (.A1(_1342_),
    .A2(_1343_),
    .B1(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__xnor2_1 _4288_ (.A(_1330_),
    .B(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4289_ (.A(_1328_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__o21a_1 _4290_ (.A1(_1328_),
    .A2(_1350_),
    .B1(_1333_),
    .X(_1352_));
 sky130_fd_sc_hd__or2_2 _4291_ (.A(_2709_),
    .B(_1336_),
    .X(_1353_));
 sky130_fd_sc_hd__buf_4 _4292_ (.A(_1349_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_4 _4293_ (.A(_2706_),
    .X(_1355_));
 sky130_fd_sc_hd__nor2_1 _4294_ (.A(_1355_),
    .B(_1354_),
    .Y(_1356_));
 sky130_fd_sc_hd__a221o_4 _4295_ (.A1(_1351_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(_1354_),
    .C1(_1356_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 _4296_ (.A(_1304_),
    .X(_1357_));
 sky130_fd_sc_hd__a22o_1 _4297_ (.A1(\cu.reg_file.reg_a[2] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[2] ),
    .X(_1358_));
 sky130_fd_sc_hd__a221o_1 _4298_ (.A1(\cu.reg_file.reg_e[2] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[2] ),
    .C1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__a21oi_1 _4299_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_1280_),
    .B1(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(_1270_),
    .B(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__a221o_1 _4301_ (.A1(_0342_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[2] ),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _4302_ (.A(\cu.reg_file.reg_e[2] ),
    .B(_1313_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_8 _4303_ (.A(_1322_),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _4304_ (.A1(\cu.reg_file.reg_sp[2] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(_0342_),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__a221o_1 _4305_ (.A1(\cu.pc.pc_o[2] ),
    .A2(_1320_),
    .B1(_1315_),
    .B2(\cu.reg_file.reg_l[2] ),
    .C1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__a211o_1 _4306_ (.A1(\cu.reg_file.reg_c[2] ),
    .A2(_1311_),
    .B1(_1363_),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__o21ai_1 _4307_ (.A1(_1357_),
    .A2(_1362_),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__clkbuf_4 _4308_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a211o_1 _4309_ (.A1(_2703_),
    .A2(_1354_),
    .B1(_1353_),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_4 _4310_ (.A(_2703_),
    .X(_1371_));
 sky130_fd_sc_hd__inv_2 _4311_ (.A(_1349_),
    .Y(_1372_));
 sky130_fd_sc_hd__o21a_2 _4312_ (.A1(_1357_),
    .A2(_1362_),
    .B1(_1367_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_4 _4313_ (.A(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__a21o_1 _4314_ (.A1(_1371_),
    .A2(_1372_),
    .B1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(\mc.rw.state[2] ),
    .B(_2701_),
    .Y(_1376_));
 sky130_fd_sc_hd__a22o_1 _4316_ (.A1(_1376_),
    .A2(_1349_),
    .B1(_1350_),
    .B2(_1328_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_1376_),
    .B(_1373_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_1330_),
    .B(_1368_),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _4319_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__xnor2_1 _4320_ (.A(_1377_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__a22o_1 _4321_ (.A1(_1370_),
    .A2(_1375_),
    .B1(_1381_),
    .B2(_1334_),
    .X(net43));
 sky130_fd_sc_hd__a21bo_1 _4322_ (.A1(_1377_),
    .A2(_1379_),
    .B1_N(_1378_),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _4323_ (.A1(\cu.reg_file.reg_a[3] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[3] ),
    .X(_1383_));
 sky130_fd_sc_hd__a221o_1 _4324_ (.A1(\cu.reg_file.reg_e[3] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[3] ),
    .C1(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__a21oi_1 _4325_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_1280_),
    .B1(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__nor2_1 _4326_ (.A(_1270_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__a221o_1 _4327_ (.A1(\cu.id.cb_opcode_y[0] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[3] ),
    .C1(_1304_),
    .X(_1387_));
 sky130_fd_sc_hd__and2_1 _4328_ (.A(\cu.reg_file.reg_l[3] ),
    .B(_1315_),
    .X(_1388_));
 sky130_fd_sc_hd__a221o_1 _4329_ (.A1(\cu.reg_file.reg_sp[3] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(\cu.id.cb_opcode_y[0] ),
    .C1(_1322_),
    .X(_1389_));
 sky130_fd_sc_hd__a221o_1 _4330_ (.A1(\cu.pc.pc_o[3] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[3] ),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__a211o_1 _4331_ (.A1(\cu.reg_file.reg_c[3] ),
    .A2(_1311_),
    .B1(_1388_),
    .C1(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__o21a_2 _4332_ (.A1(_1386_),
    .A2(_1387_),
    .B1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__or2_1 _4333_ (.A(_1376_),
    .B(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_1382_),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__clkbuf_4 _4335_ (.A(_1376_),
    .X(_1395_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(_1395_),
    .B(_1392_),
    .Y(_1396_));
 sky130_fd_sc_hd__or2b_1 _4337_ (.A(_1394_),
    .B_N(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__a21o_1 _4338_ (.A1(_1396_),
    .A2(_1393_),
    .B1(_1382_),
    .X(_1398_));
 sky130_fd_sc_hd__buf_2 _4339_ (.A(_1392_),
    .X(_1399_));
 sky130_fd_sc_hd__nor2_4 _4340_ (.A(_1349_),
    .B(_1373_),
    .Y(_1400_));
 sky130_fd_sc_hd__nor2_2 _4341_ (.A(_2709_),
    .B(_1336_),
    .Y(_1401_));
 sky130_fd_sc_hd__o21ai_1 _4342_ (.A1(_1355_),
    .A2(_1400_),
    .B1(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__and2b_1 _4343_ (.A_N(_1392_),
    .B(_1400_),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(_1399_),
    .A2(_1402_),
    .B1(_1403_),
    .B2(_1371_),
    .X(_1404_));
 sky130_fd_sc_hd__a31o_2 _4345_ (.A1(_1334_),
    .A2(_1397_),
    .A3(_1398_),
    .B1(_1404_),
    .X(net44));
 sky130_fd_sc_hd__a22o_1 _4346_ (.A1(\cu.reg_file.reg_a[4] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[4] ),
    .X(_1405_));
 sky130_fd_sc_hd__a221o_1 _4347_ (.A1(\cu.reg_file.reg_e[4] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[4] ),
    .C1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__a21oi_1 _4348_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_1280_),
    .B1(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__nor2_1 _4349_ (.A(_1270_),
    .B(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__a221o_2 _4350_ (.A1(_0374_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[4] ),
    .C1(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__and2_1 _4351_ (.A(\cu.reg_file.reg_l[4] ),
    .B(_1315_),
    .X(_1410_));
 sky130_fd_sc_hd__a221o_1 _4352_ (.A1(\cu.reg_file.reg_sp[4] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(_0374_),
    .C1(_1364_),
    .X(_1411_));
 sky130_fd_sc_hd__a221o_1 _4353_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[4] ),
    .C1(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__a211o_2 _4354_ (.A1(\cu.reg_file.reg_c[4] ),
    .A2(_1311_),
    .B1(_1410_),
    .C1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__o21ai_4 _4355_ (.A1(_1357_),
    .A2(_1409_),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_1403_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__o21a_4 _4357_ (.A1(_1357_),
    .A2(_1409_),
    .B1(_1413_),
    .X(_1416_));
 sky130_fd_sc_hd__o21ai_1 _4358_ (.A1(_1355_),
    .A2(_1403_),
    .B1(_1401_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_1395_),
    .B(_1416_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(_1330_),
    .B(_1414_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _4362_ (.A(_1419_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__a21o_1 _4363_ (.A1(_1396_),
    .A2(_1394_),
    .B1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_1333_),
    .B(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__a31o_1 _4365_ (.A1(_1396_),
    .A2(_1394_),
    .A3(_1421_),
    .B1(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__o211ai_2 _4366_ (.A1(_1355_),
    .A2(_1415_),
    .B1(_1418_),
    .C1(_1424_),
    .Y(net45));
 sky130_fd_sc_hd__a22o_1 _4367_ (.A1(\cu.reg_file.reg_a[5] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[5] ),
    .X(_1425_));
 sky130_fd_sc_hd__a221o_1 _4368_ (.A1(\cu.reg_file.reg_e[5] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[5] ),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a21oi_1 _4369_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_1280_),
    .B1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nor2_1 _4370_ (.A(_1270_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__a221o_1 _4371_ (.A1(_0373_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[5] ),
    .C1(_1357_),
    .X(_1429_));
 sky130_fd_sc_hd__and2_1 _4372_ (.A(\cu.reg_file.reg_l[5] ),
    .B(_1315_),
    .X(_1430_));
 sky130_fd_sc_hd__a221o_1 _4373_ (.A1(\cu.reg_file.reg_sp[5] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(_0373_),
    .C1(_1364_),
    .X(_1431_));
 sky130_fd_sc_hd__a221o_1 _4374_ (.A1(\cu.pc.pc_o[5] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[5] ),
    .C1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a211o_1 _4375_ (.A1(\cu.reg_file.reg_c[5] ),
    .A2(_1311_),
    .B1(_1430_),
    .C1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__o21a_2 _4376_ (.A1(_1428_),
    .A2(_1429_),
    .B1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__nor2_1 _4377_ (.A(_1416_),
    .B(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(_1403_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__a21bo_1 _4379_ (.A1(_1415_),
    .A2(_1434_),
    .B1_N(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__or2_1 _4380_ (.A(_1395_),
    .B(_1434_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(_1395_),
    .B(_1434_),
    .Y(_1439_));
 sky130_fd_sc_hd__and2_1 _4382_ (.A(_1438_),
    .B(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand2_1 _4383_ (.A(_1419_),
    .B(_1422_),
    .Y(_1441_));
 sky130_fd_sc_hd__o21ai_1 _4384_ (.A1(_1440_),
    .A2(_1441_),
    .B1(_1333_),
    .Y(_1442_));
 sky130_fd_sc_hd__a21oi_1 _4385_ (.A1(_1440_),
    .A2(_1441_),
    .B1(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a221o_4 _4386_ (.A1(_1353_),
    .A2(_1434_),
    .B1(_1437_),
    .B2(_1371_),
    .C1(_1443_),
    .X(net46));
 sky130_fd_sc_hd__or2b_1 _4387_ (.A(_1422_),
    .B_N(_1440_),
    .X(_1444_));
 sky130_fd_sc_hd__a22o_1 _4388_ (.A1(\cu.reg_file.reg_a[6] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[6] ),
    .X(_1445_));
 sky130_fd_sc_hd__a221o_1 _4389_ (.A1(\cu.reg_file.reg_e[6] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[6] ),
    .C1(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__a21oi_1 _4390_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_1280_),
    .B1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(_1270_),
    .B(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a221o_1 _4392_ (.A1(_0387_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[6] ),
    .C1(_1357_),
    .X(_1449_));
 sky130_fd_sc_hd__and2_1 _4393_ (.A(\cu.reg_file.reg_l[6] ),
    .B(_1315_),
    .X(_1450_));
 sky130_fd_sc_hd__a221o_1 _4394_ (.A1(\cu.reg_file.reg_sp[6] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(_0387_),
    .C1(_1322_),
    .X(_1451_));
 sky130_fd_sc_hd__a221o_1 _4395_ (.A1(\cu.pc.pc_o[6] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[6] ),
    .C1(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__a211o_1 _4396_ (.A1(\cu.reg_file.reg_c[6] ),
    .A2(_1311_),
    .B1(_1450_),
    .C1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__o21a_2 _4397_ (.A1(_1448_),
    .A2(_1449_),
    .B1(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__xnor2_1 _4398_ (.A(_1395_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__a31o_1 _4399_ (.A1(_1419_),
    .A2(_1439_),
    .A3(_1444_),
    .B1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__nand4_1 _4400_ (.A(_1419_),
    .B(_1439_),
    .C(_1455_),
    .D(_1444_),
    .Y(_1457_));
 sky130_fd_sc_hd__a21o_1 _4401_ (.A1(_2703_),
    .A2(_1436_),
    .B1(_1353_),
    .X(_1458_));
 sky130_fd_sc_hd__nor2_1 _4402_ (.A(_1436_),
    .B(_1454_),
    .Y(_1459_));
 sky130_fd_sc_hd__a22o_1 _4403_ (.A1(_1454_),
    .A2(_1458_),
    .B1(_1459_),
    .B2(_1371_),
    .X(_1460_));
 sky130_fd_sc_hd__a31o_1 _4404_ (.A1(_1334_),
    .A2(_1456_),
    .A3(_1457_),
    .B1(_1460_),
    .X(net47));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(_1454_),
    .Y(_1461_));
 sky130_fd_sc_hd__o21a_1 _4406_ (.A1(_1331_),
    .A2(_1461_),
    .B1(_1456_),
    .X(_1462_));
 sky130_fd_sc_hd__a22o_1 _4407_ (.A1(\cu.reg_file.reg_a[7] ),
    .A2(_1277_),
    .B1(_1286_),
    .B2(\cu.reg_file.reg_sp[7] ),
    .X(_1463_));
 sky130_fd_sc_hd__a221o_1 _4408_ (.A1(\cu.reg_file.reg_e[7] ),
    .A2(_1282_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_l[7] ),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__a21oi_1 _4409_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_1280_),
    .B1(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _4410_ (.A(_1270_),
    .B(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__a221o_1 _4411_ (.A1(\cu.id.cb_opcode_x[1] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[7] ),
    .C1(_1304_),
    .X(_1467_));
 sky130_fd_sc_hd__and2_1 _4412_ (.A(\cu.reg_file.reg_l[7] ),
    .B(_1315_),
    .X(_1468_));
 sky130_fd_sc_hd__a221o_1 _4413_ (.A1(\cu.reg_file.reg_sp[7] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(\cu.id.cb_opcode_x[1] ),
    .C1(_1322_),
    .X(_1469_));
 sky130_fd_sc_hd__a221o_1 _4414_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_e[7] ),
    .C1(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__a211o_1 _4415_ (.A1(\cu.reg_file.reg_c[7] ),
    .A2(_1311_),
    .B1(_1468_),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__o21ai_4 _4416_ (.A1(_1466_),
    .A2(_1467_),
    .B1(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__xnor2_1 _4417_ (.A(_1330_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__or2_1 _4418_ (.A(_1462_),
    .B(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_1462_),
    .B(_1473_),
    .Y(_1475_));
 sky130_fd_sc_hd__o21a_1 _4420_ (.A1(_1355_),
    .A2(_1459_),
    .B1(_1401_),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(_1459_),
    .B(_1472_),
    .Y(_1477_));
 sky130_fd_sc_hd__o22ai_1 _4422_ (.A1(_1472_),
    .A2(_1476_),
    .B1(_1477_),
    .B2(_1355_),
    .Y(_1478_));
 sky130_fd_sc_hd__a31o_1 _4423_ (.A1(_1334_),
    .A2(_1474_),
    .A3(_1475_),
    .B1(_1478_),
    .X(net48));
 sky130_fd_sc_hd__a31o_1 _4424_ (.A1(_1435_),
    .A2(_1461_),
    .A3(_1472_),
    .B1(_1330_),
    .X(_1479_));
 sky130_fd_sc_hd__or3_1 _4425_ (.A(_1455_),
    .B(_1444_),
    .C(_1473_),
    .X(_1480_));
 sky130_fd_sc_hd__or2_1 _4426_ (.A(\cu.id.state[1] ),
    .B(\cu.id.state[0] ),
    .X(_1481_));
 sky130_fd_sc_hd__or2_2 _4427_ (.A(_1267_),
    .B(_2951_),
    .X(_1482_));
 sky130_fd_sc_hd__nand2_2 _4428_ (.A(_1481_),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__or2_4 _4429_ (.A(_1268_),
    .B(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__a22o_1 _4430_ (.A1(\cu.reg_file.reg_d[0] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[8] ),
    .X(_1485_));
 sky130_fd_sc_hd__a221o_1 _4431_ (.A1(\cu.reg_file.reg_b[0] ),
    .A2(net144),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[0] ),
    .C1(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__nor2_2 _4432_ (.A(_1268_),
    .B(_1483_),
    .Y(_1487_));
 sky130_fd_sc_hd__clkbuf_8 _4433_ (.A(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__a221o_1 _4434_ (.A1(\cu.id.imm_i[8] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\cu.pc.pc_o[8] ),
    .C1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__a21o_1 _4435_ (.A1(_1295_),
    .A2(_1486_),
    .B1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__o21a_1 _4436_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_1484_),
    .B1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a221o_1 _4437_ (.A1(\cu.reg_file.reg_sp[8] ),
    .A2(_0992_),
    .B1(_1338_),
    .B2(\cu.id.imm_i[8] ),
    .C1(_1321_),
    .X(_1492_));
 sky130_fd_sc_hd__a221o_1 _4438_ (.A1(\cu.pc.pc_o[8] ),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[0] ),
    .C1(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__a221o_1 _4439_ (.A1(\cu.reg_file.reg_h[0] ),
    .A2(_1314_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[0] ),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__o21a_1 _4440_ (.A1(_1304_),
    .A2(_1491_),
    .B1(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_1395_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__or2_1 _4442_ (.A(_1395_),
    .B(_1495_),
    .X(_1497_));
 sky130_fd_sc_hd__nand2_1 _4443_ (.A(_1496_),
    .B(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a21o_1 _4444_ (.A1(_1479_),
    .A2(_1480_),
    .B1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__nand3_1 _4445_ (.A(_1498_),
    .B(_1479_),
    .C(_1480_),
    .Y(_1500_));
 sky130_fd_sc_hd__a21o_1 _4446_ (.A1(_2703_),
    .A2(_1477_),
    .B1(_1353_),
    .X(_1501_));
 sky130_fd_sc_hd__nor2_1 _4447_ (.A(_1477_),
    .B(_1495_),
    .Y(_1502_));
 sky130_fd_sc_hd__a22o_1 _4448_ (.A1(_1495_),
    .A2(_1501_),
    .B1(_1502_),
    .B2(_1371_),
    .X(_1503_));
 sky130_fd_sc_hd__a31o_2 _4449_ (.A1(_1334_),
    .A2(_1499_),
    .A3(_1500_),
    .B1(_1503_),
    .X(net49));
 sky130_fd_sc_hd__a22o_1 _4450_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_1286_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[1] ),
    .X(_1504_));
 sky130_fd_sc_hd__a22o_1 _4451_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_1280_),
    .B1(_1282_),
    .B2(\cu.reg_file.reg_d[1] ),
    .X(_1505_));
 sky130_fd_sc_hd__o21a_1 _4452_ (.A1(_1504_),
    .A2(_1505_),
    .B1(_1295_),
    .X(_1506_));
 sky130_fd_sc_hd__a221o_1 _4453_ (.A1(\cu.id.imm_i[9] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[9] ),
    .C1(_1303_),
    .X(_1507_));
 sky130_fd_sc_hd__and2_1 _4454_ (.A(\cu.reg_file.reg_h[1] ),
    .B(_1314_),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_1 _4455_ (.A1(\cu.reg_file.reg_sp[9] ),
    .A2(_0993_),
    .B1(_1339_),
    .B2(\cu.id.imm_i[9] ),
    .C1(_1322_),
    .X(_1509_));
 sky130_fd_sc_hd__a221o_1 _4456_ (.A1(\cu.pc.pc_o[9] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_d[1] ),
    .C1(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__a211o_1 _4457_ (.A1(\cu.reg_file.reg_b[1] ),
    .A2(_1311_),
    .B1(_1508_),
    .C1(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__o21ai_2 _4458_ (.A1(_1506_),
    .A2(_1507_),
    .B1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__or2_1 _4459_ (.A(_1330_),
    .B(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_1330_),
    .B(_1512_),
    .Y(_1514_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_1513_),
    .B(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__nand3_1 _4462_ (.A(_1496_),
    .B(_1499_),
    .C(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a21o_1 _4463_ (.A1(_1496_),
    .A2(_1499_),
    .B1(_1515_),
    .X(_1517_));
 sky130_fd_sc_hd__o21a_1 _4464_ (.A1(_2706_),
    .A2(_1502_),
    .B1(_1401_),
    .X(_1518_));
 sky130_fd_sc_hd__and2_1 _4465_ (.A(_1502_),
    .B(_1512_),
    .X(_1519_));
 sky130_fd_sc_hd__a2bb2o_1 _4466_ (.A1_N(_1512_),
    .A2_N(_1518_),
    .B1(_1519_),
    .B2(_1371_),
    .X(_1520_));
 sky130_fd_sc_hd__a31o_1 _4467_ (.A1(_1334_),
    .A2(_1516_),
    .A3(_1517_),
    .B1(_1520_),
    .X(net50));
 sky130_fd_sc_hd__a21bo_1 _4468_ (.A1(_1496_),
    .A2(_1499_),
    .B1_N(_1514_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_4 _4469_ (.A(\cu.pc.pc_o[10] ),
    .X(_1522_));
 sky130_fd_sc_hd__a22o_1 _4470_ (.A1(\cu.reg_file.reg_d[2] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[10] ),
    .X(_1523_));
 sky130_fd_sc_hd__a221o_1 _4471_ (.A1(\cu.reg_file.reg_b[2] ),
    .A2(net143),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[2] ),
    .C1(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__a221o_1 _4472_ (.A1(\cu.id.imm_i[10] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(_1522_),
    .C1(_1488_),
    .X(_1525_));
 sky130_fd_sc_hd__a21o_1 _4473_ (.A1(_1295_),
    .A2(_1524_),
    .B1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__o21a_1 _4474_ (.A1(_1522_),
    .A2(_1484_),
    .B1(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_1 _4475_ (.A1(\cu.reg_file.reg_sp[10] ),
    .A2(_0992_),
    .B1(_1338_),
    .B2(\cu.id.imm_i[10] ),
    .C1(_1321_),
    .X(_1528_));
 sky130_fd_sc_hd__a221o_1 _4476_ (.A1(_1522_),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[2] ),
    .C1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__a221o_1 _4477_ (.A1(\cu.reg_file.reg_h[2] ),
    .A2(_1314_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[2] ),
    .C1(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__o21ai_4 _4478_ (.A1(_1304_),
    .A2(_1527_),
    .B1(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__xnor2_1 _4479_ (.A(_1330_),
    .B(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__a21o_1 _4480_ (.A1(_1513_),
    .A2(_1521_),
    .B1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__nand3_1 _4481_ (.A(_1513_),
    .B(_1532_),
    .C(_1521_),
    .Y(_1534_));
 sky130_fd_sc_hd__o21a_1 _4482_ (.A1(_1355_),
    .A2(_1519_),
    .B1(_1401_),
    .X(_1535_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_1519_),
    .B(_1531_),
    .Y(_1536_));
 sky130_fd_sc_hd__o22ai_1 _4484_ (.A1(_1531_),
    .A2(_1535_),
    .B1(_1536_),
    .B2(_1355_),
    .Y(_1537_));
 sky130_fd_sc_hd__a31o_2 _4485_ (.A1(_1334_),
    .A2(_1533_),
    .A3(_1534_),
    .B1(_1537_),
    .X(net36));
 sky130_fd_sc_hd__a22o_1 _4486_ (.A1(\cu.reg_file.reg_d[3] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[11] ),
    .X(_1538_));
 sky130_fd_sc_hd__a221o_1 _4487_ (.A1(\cu.reg_file.reg_b[3] ),
    .A2(net143),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[3] ),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__a221o_1 _4488_ (.A1(\cu.id.imm_i[11] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\cu.pc.pc_o[11] ),
    .C1(_1488_),
    .X(_1540_));
 sky130_fd_sc_hd__a21o_1 _4489_ (.A1(_1295_),
    .A2(_1539_),
    .B1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__o21a_1 _4490_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1484_),
    .B1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__a221o_1 _4491_ (.A1(\cu.reg_file.reg_sp[11] ),
    .A2(_0992_),
    .B1(_1339_),
    .B2(\cu.id.imm_i[11] ),
    .C1(_1322_),
    .X(_1543_));
 sky130_fd_sc_hd__a221o_1 _4492_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[3] ),
    .C1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__a221o_1 _4493_ (.A1(\cu.reg_file.reg_h[3] ),
    .A2(_1315_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[3] ),
    .C1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__o21ai_4 _4494_ (.A1(_1304_),
    .A2(_1542_),
    .B1(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__or2_1 _4495_ (.A(_1331_),
    .B(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__nand2_1 _4496_ (.A(_1331_),
    .B(_1546_),
    .Y(_1548_));
 sky130_fd_sc_hd__nand2_1 _4497_ (.A(_1547_),
    .B(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__o21a_1 _4498_ (.A1(_1330_),
    .A2(_1531_),
    .B1(_1533_),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_1549_),
    .B(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__or2_1 _4500_ (.A(_1549_),
    .B(_1550_),
    .X(_1552_));
 sky130_fd_sc_hd__xor2_1 _4501_ (.A(_1536_),
    .B(_1546_),
    .X(_1553_));
 sky130_fd_sc_hd__a2bb2o_1 _4502_ (.A1_N(_1401_),
    .A2_N(_1546_),
    .B1(_1553_),
    .B2(_1371_),
    .X(_1554_));
 sky130_fd_sc_hd__a31o_1 _4503_ (.A1(_1334_),
    .A2(_1551_),
    .A3(_1552_),
    .B1(_1554_),
    .X(net37));
 sky130_fd_sc_hd__a22o_1 _4504_ (.A1(\cu.reg_file.reg_d[4] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[12] ),
    .X(_1555_));
 sky130_fd_sc_hd__a221o_1 _4505_ (.A1(\cu.reg_file.reg_b[4] ),
    .A2(net143),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[4] ),
    .C1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__a221o_1 _4506_ (.A1(\cu.id.imm_i[12] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\cu.pc.pc_o[12] ),
    .C1(_1487_),
    .X(_1557_));
 sky130_fd_sc_hd__a21o_1 _4507_ (.A1(_1295_),
    .A2(_1556_),
    .B1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__o21a_1 _4508_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_1484_),
    .B1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__a221o_1 _4509_ (.A1(\cu.reg_file.reg_sp[12] ),
    .A2(_0992_),
    .B1(_1338_),
    .B2(\cu.id.imm_i[12] ),
    .C1(_1321_),
    .X(_1560_));
 sky130_fd_sc_hd__a221o_1 _4510_ (.A1(\cu.pc.pc_o[12] ),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[4] ),
    .C1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__a221o_1 _4511_ (.A1(\cu.reg_file.reg_h[4] ),
    .A2(_1314_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[4] ),
    .C1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__o21ai_4 _4512_ (.A1(_1304_),
    .A2(_1559_),
    .B1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__xnor2_1 _4513_ (.A(_1331_),
    .B(_1563_),
    .Y(_1564_));
 sky130_fd_sc_hd__a21o_1 _4514_ (.A1(_1331_),
    .A2(_1546_),
    .B1(_1550_),
    .X(_1565_));
 sky130_fd_sc_hd__nand3_1 _4515_ (.A(_1547_),
    .B(_1564_),
    .C(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__a21o_1 _4516_ (.A1(_1547_),
    .A2(_1565_),
    .B1(_1564_),
    .X(_1567_));
 sky130_fd_sc_hd__and3_1 _4517_ (.A(_1519_),
    .B(_1531_),
    .C(_1546_),
    .X(_1568_));
 sky130_fd_sc_hd__xnor2_1 _4518_ (.A(_1568_),
    .B(_1563_),
    .Y(_1569_));
 sky130_fd_sc_hd__a2bb2o_1 _4519_ (.A1_N(_1401_),
    .A2_N(_1563_),
    .B1(_1569_),
    .B2(_1371_),
    .X(_1570_));
 sky130_fd_sc_hd__a31o_1 _4520_ (.A1(_1334_),
    .A2(_1566_),
    .A3(_1567_),
    .B1(_1570_),
    .X(net38));
 sky130_fd_sc_hd__a22o_1 _4521_ (.A1(\cu.reg_file.reg_d[5] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[13] ),
    .X(_1571_));
 sky130_fd_sc_hd__a221o_1 _4522_ (.A1(\cu.reg_file.reg_b[5] ),
    .A2(net143),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[5] ),
    .C1(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__a221o_1 _4523_ (.A1(\cu.id.imm_i[13] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\cu.pc.pc_o[13] ),
    .C1(_1487_),
    .X(_1573_));
 sky130_fd_sc_hd__a21o_1 _4524_ (.A1(_1295_),
    .A2(_1572_),
    .B1(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__o21a_1 _4525_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1484_),
    .B1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__a221o_1 _4526_ (.A1(\cu.reg_file.reg_sp[13] ),
    .A2(_0992_),
    .B1(_1338_),
    .B2(\cu.id.imm_i[13] ),
    .C1(_1321_),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_1 _4527_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[5] ),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a221o_1 _4528_ (.A1(\cu.reg_file.reg_h[5] ),
    .A2(_1314_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[5] ),
    .C1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o21a_2 _4529_ (.A1(_1303_),
    .A2(_1575_),
    .B1(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__or2_1 _4530_ (.A(_1395_),
    .B(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_1395_),
    .B(_1579_),
    .Y(_1581_));
 sky130_fd_sc_hd__o21ai_2 _4532_ (.A1(_1331_),
    .A2(_1563_),
    .B1(_1567_),
    .Y(_1582_));
 sky130_fd_sc_hd__a21o_1 _4533_ (.A1(_1580_),
    .A2(_1581_),
    .B1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__nor2_1 _4534_ (.A(_2699_),
    .B(_1331_),
    .Y(_1584_));
 sky130_fd_sc_hd__a31oi_1 _4535_ (.A1(_1580_),
    .A2(_1581_),
    .A3(_1582_),
    .B1(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_1568_),
    .B(_1563_),
    .Y(_1586_));
 sky130_fd_sc_hd__or2_1 _4537_ (.A(_1586_),
    .B(_1579_),
    .X(_1587_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(_1586_),
    .B(_1579_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21oi_1 _4539_ (.A1(_1587_),
    .A2(_1588_),
    .B1(_1355_),
    .Y(_1589_));
 sky130_fd_sc_hd__a221o_1 _4540_ (.A1(_1353_),
    .A2(_1579_),
    .B1(_1583_),
    .B2(_1585_),
    .C1(_1589_),
    .X(net39));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(_1580_),
    .B(_1582_),
    .Y(_1590_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1285_),
    .Y(_1591_));
 sky130_fd_sc_hd__a21bo_1 _4543_ (.A1(\cu.reg_file.reg_d[6] ),
    .A2(_1282_),
    .B1_N(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__a221o_1 _4544_ (.A1(\cu.reg_file.reg_b[6] ),
    .A2(net143),
    .B1(_1283_),
    .B2(\cu.reg_file.reg_h[6] ),
    .C1(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__a221o_1 _4545_ (.A1(\cu.id.imm_i[14] ),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\cu.pc.pc_o[14] ),
    .C1(_1488_),
    .X(_1594_));
 sky130_fd_sc_hd__a21o_1 _4546_ (.A1(_1295_),
    .A2(_1593_),
    .B1(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__o21a_1 _4547_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1484_),
    .B1(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__a221o_1 _4548_ (.A1(\cu.reg_file.reg_sp[14] ),
    .A2(_0992_),
    .B1(_1338_),
    .B2(\cu.id.imm_i[14] ),
    .C1(_1322_),
    .X(_1597_));
 sky130_fd_sc_hd__a221o_1 _4549_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1319_),
    .B1(_1312_),
    .B2(\cu.reg_file.reg_d[6] ),
    .C1(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__a221o_1 _4550_ (.A1(\cu.reg_file.reg_h[6] ),
    .A2(_1314_),
    .B1(_1310_),
    .B2(\cu.reg_file.reg_b[6] ),
    .C1(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__o21ai_4 _4551_ (.A1(_1304_),
    .A2(_1596_),
    .B1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__nor2_1 _4552_ (.A(_1331_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__and2_1 _4553_ (.A(_1331_),
    .B(_1600_),
    .X(_1602_));
 sky130_fd_sc_hd__or2_1 _4554_ (.A(_1601_),
    .B(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__a21oi_2 _4555_ (.A1(_1581_),
    .A2(_1590_),
    .B1(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__a31o_1 _4556_ (.A1(_1581_),
    .A2(_1603_),
    .A3(_1590_),
    .B1(_1584_),
    .X(_1605_));
 sky130_fd_sc_hd__xnor2_1 _4557_ (.A(_1587_),
    .B(_1600_),
    .Y(_1606_));
 sky130_fd_sc_hd__o22a_1 _4558_ (.A1(_1401_),
    .A2(_1600_),
    .B1(_1606_),
    .B2(_1355_),
    .X(_1607_));
 sky130_fd_sc_hd__o21ai_4 _4559_ (.A1(_1604_),
    .A2(_1605_),
    .B1(_1607_),
    .Y(net40));
 sky130_fd_sc_hd__a22o_1 _4560_ (.A1(\cu.reg_file.reg_d[7] ),
    .A2(_1281_),
    .B1(_1285_),
    .B2(\cu.reg_file.reg_sp[15] ),
    .X(_1608_));
 sky130_fd_sc_hd__a221o_1 _4561_ (.A1(\cu.reg_file.reg_b[7] ),
    .A2(_1280_),
    .B1(_1284_),
    .B2(\cu.reg_file.reg_h[7] ),
    .C1(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__a221o_1 _4562_ (.A1(\cu.id.imm_i[15] ),
    .A2(_1294_),
    .B1(_1297_),
    .B2(\cu.pc.pc_o[15] ),
    .C1(_1488_),
    .X(_1610_));
 sky130_fd_sc_hd__a21o_1 _4563_ (.A1(_1295_),
    .A2(_1609_),
    .B1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__o21a_1 _4564_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_1484_),
    .B1(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__a221o_1 _4565_ (.A1(\cu.reg_file.reg_sp[15] ),
    .A2(_0992_),
    .B1(_1339_),
    .B2(\cu.id.imm_i[15] ),
    .C1(_1322_),
    .X(_1613_));
 sky130_fd_sc_hd__a221o_1 _4566_ (.A1(\cu.pc.pc_o[15] ),
    .A2(_1320_),
    .B1(_1313_),
    .B2(\cu.reg_file.reg_d[7] ),
    .C1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__a221o_1 _4567_ (.A1(\cu.reg_file.reg_h[7] ),
    .A2(_1315_),
    .B1(_1311_),
    .B2(\cu.reg_file.reg_b[7] ),
    .C1(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__o21ai_4 _4568_ (.A1(_1304_),
    .A2(_1612_),
    .B1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__xnor2_1 _4569_ (.A(_1395_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__o21ai_1 _4570_ (.A1(_1601_),
    .A2(_1604_),
    .B1(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__or3_1 _4571_ (.A(_1601_),
    .B(_1604_),
    .C(_1617_),
    .X(_1619_));
 sky130_fd_sc_hd__and2b_1 _4572_ (.A_N(_1587_),
    .B(_1600_),
    .X(_1620_));
 sky130_fd_sc_hd__o21a_1 _4573_ (.A1(_2706_),
    .A2(_1620_),
    .B1(_1401_),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_1 _4574_ (.A(_1616_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__a31o_1 _4575_ (.A1(_1371_),
    .A2(_1620_),
    .A3(_1616_),
    .B1(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__a31o_1 _4576_ (.A1(_1333_),
    .A2(_1618_),
    .A3(_1619_),
    .B1(_1623_),
    .X(net41));
 sky130_fd_sc_hd__and2_4 _4577_ (.A(_0824_),
    .B(_0818_),
    .X(_1624_));
 sky130_fd_sc_hd__a22o_1 _4578_ (.A1(_2704_),
    .A2(_0618_),
    .B1(_1624_),
    .B2(_2699_),
    .X(net51));
 sky130_fd_sc_hd__nor2_4 _4579_ (.A(_0517_),
    .B(_1229_),
    .Y(_1625_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(_2704_),
    .A2(_1050_),
    .B1(_1625_),
    .B2(_2699_),
    .X(net52));
 sky130_fd_sc_hd__a22o_1 _4581_ (.A1(_2704_),
    .A2(_1072_),
    .B1(_1225_),
    .B2(_2699_),
    .X(net53));
 sky130_fd_sc_hd__a22o_1 _4582_ (.A1(_2704_),
    .A2(_1187_),
    .B1(_1221_),
    .B2(_2699_),
    .X(net54));
 sky130_fd_sc_hd__a22o_1 _4583_ (.A1(_2704_),
    .A2(_1189_),
    .B1(_1212_),
    .B2(_2699_),
    .X(net55));
 sky130_fd_sc_hd__a22o_1 _4584_ (.A1(_2704_),
    .A2(_1191_),
    .B1(_1208_),
    .B2(_2699_),
    .X(net56));
 sky130_fd_sc_hd__nor2_2 _4585_ (.A(_0517_),
    .B(_1199_),
    .Y(_1626_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(_2704_),
    .A2(_1193_),
    .B1(_1626_),
    .B2(_2699_),
    .X(net57));
 sky130_fd_sc_hd__a22o_1 _4587_ (.A1(_2704_),
    .A2(_1260_),
    .B1(_1262_),
    .B2(_2699_),
    .X(net58));
 sky130_fd_sc_hd__nand2_4 _4588_ (.A(_1327_),
    .B(_1372_),
    .Y(_1627_));
 sky130_fd_sc_hd__inv_2 _4589_ (.A(_1579_),
    .Y(_1628_));
 sky130_fd_sc_hd__or4_1 _4590_ (.A(_1563_),
    .B(_1628_),
    .C(_1600_),
    .D(_1616_),
    .X(_1629_));
 sky130_fd_sc_hd__or4b_1 _4591_ (.A(_1512_),
    .B(_1531_),
    .C(_1546_),
    .D_N(_1495_),
    .X(_1630_));
 sky130_fd_sc_hd__or3_4 _4592_ (.A(_1392_),
    .B(_1629_),
    .C(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__or4_4 _4593_ (.A(_1434_),
    .B(_1461_),
    .C(_1472_),
    .D(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__a211oi_2 _4594_ (.A1(_1374_),
    .A2(_1627_),
    .B1(_1632_),
    .C1(_1414_),
    .Y(_1633_));
 sky130_fd_sc_hd__or2_2 _4595_ (.A(\mc.cl.cmp_o ),
    .B(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__nand2_4 _4596_ (.A(_1327_),
    .B(_1400_),
    .Y(_1635_));
 sky130_fd_sc_hd__or3_2 _4597_ (.A(_1416_),
    .B(_1632_),
    .C(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_1 _4598_ (.A(_1454_),
    .B(_1472_),
    .Y(_1637_));
 sky130_fd_sc_hd__or3b_2 _4599_ (.A(_1434_),
    .B(_1631_),
    .C_N(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_1434_),
    .B(_1637_),
    .Y(_1639_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_1327_),
    .B(_1372_),
    .Y(_1640_));
 sky130_fd_sc_hd__or4_1 _4602_ (.A(_1373_),
    .B(_1414_),
    .C(_1639_),
    .D(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__nor2_1 _4603_ (.A(_1631_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__clkinv_4 _4604_ (.A(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__or3_2 _4605_ (.A(_1416_),
    .B(_1631_),
    .C(_1639_),
    .X(_1644_));
 sky130_fd_sc_hd__nand4_4 _4606_ (.A(_1636_),
    .B(_1638_),
    .C(_1643_),
    .D(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__nor2_4 _4607_ (.A(_1634_),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__a21o_1 _4608_ (.A1(_1364_),
    .A2(_1488_),
    .B1(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__buf_2 _4609_ (.A(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__buf_2 _4610_ (.A(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__buf_2 _4611_ (.A(_1484_),
    .X(_1650_));
 sky130_fd_sc_hd__buf_2 _4612_ (.A(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_4 _4613_ (.A(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__nor3_1 _4614_ (.A(\mc.rw.state[2] ),
    .B(\mc.rw.state[1] ),
    .C(\mc.rw.state[0] ),
    .Y(_1653_));
 sky130_fd_sc_hd__nor4_1 _4615_ (.A(\mc.cc.count[2] ),
    .B(\mc.cc.count[1] ),
    .C(\mc.cc.count[3] ),
    .D(\mc.cc.count[0] ),
    .Y(_1654_));
 sky130_fd_sc_hd__nand2_2 _4616_ (.A(\mc.cc.enable_edge_detector.prev_data ),
    .B(net149),
    .Y(_1655_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(_2703_),
    .A1(_2709_),
    .S(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__a31o_1 _4618_ (.A1(_1652_),
    .A2(_1646_),
    .A3(_1653_),
    .B1(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__a21o_1 _4619_ (.A1(_2707_),
    .A2(_1649_),
    .B1(_1657_),
    .X(\mc.rw.next_state[0] ));
 sky130_fd_sc_hd__a21oi_4 _4620_ (.A1(_1364_),
    .A2(_1488_),
    .B1(_1646_),
    .Y(_1658_));
 sky130_fd_sc_hd__clkbuf_8 _4621_ (.A(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__or3_1 _4622_ (.A(\mc.cl.cmp_o ),
    .B(_1364_),
    .C(_1616_),
    .X(_1660_));
 sky130_fd_sc_hd__inv_2 _4623_ (.A(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__or3_2 _4624_ (.A(_0297_),
    .B(_2921_),
    .C(_0379_),
    .X(_1662_));
 sky130_fd_sc_hd__or2_1 _4625_ (.A(_2934_),
    .B(_2906_),
    .X(_1663_));
 sky130_fd_sc_hd__nor3b_4 _4626_ (.A(_0314_),
    .B(_1662_),
    .C_N(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__clkbuf_4 _4627_ (.A(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(_1652_),
    .A1(_1661_),
    .S(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__a21oi_1 _4629_ (.A1(_1653_),
    .A2(_1666_),
    .B1(_2701_),
    .Y(_1667_));
 sky130_fd_sc_hd__o21ai_1 _4630_ (.A1(_1659_),
    .A2(_1667_),
    .B1(_2710_),
    .Y(\mc.rw.next_state[1] ));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(_1655_),
    .Y(_1668_));
 sky130_fd_sc_hd__or3b_4 _4632_ (.A(_0314_),
    .B(_1662_),
    .C_N(_1663_),
    .X(_1669_));
 sky130_fd_sc_hd__buf_4 _4633_ (.A(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_8 _4634_ (.A(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__a31o_1 _4635_ (.A1(_1653_),
    .A2(_1671_),
    .A3(_1661_),
    .B1(_1333_),
    .X(_1672_));
 sky130_fd_sc_hd__a221o_1 _4636_ (.A1(_2709_),
    .A2(_1668_),
    .B1(_1672_),
    .B2(_1649_),
    .C1(_1371_),
    .X(\mc.rw.next_state[2] ));
 sky130_fd_sc_hd__and2_1 _4637_ (.A(\ih.t.enable ),
    .B(_2860_),
    .X(_1673_));
 sky130_fd_sc_hd__clkbuf_4 _4638_ (.A(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__and2b_1 _4639_ (.A_N(\ih.t.count[0] ),
    .B(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _4640_ (.A(_1675_),
    .X(\ih.t.next_count[0] ));
 sky130_fd_sc_hd__clkbuf_4 _4641_ (.A(_1673_),
    .X(_1676_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .Y(_1677_));
 sky130_fd_sc_hd__or2_1 _4643_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .X(_1678_));
 sky130_fd_sc_hd__and3_1 _4644_ (.A(_1676_),
    .B(_1677_),
    .C(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _4645_ (.A(_1679_),
    .X(\ih.t.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _4646_ (.A1(\ih.t.count[0] ),
    .A2(\ih.t.count[1] ),
    .B1(\ih.t.count[2] ),
    .X(_1680_));
 sky130_fd_sc_hd__nand3_1 _4647_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .C(\ih.t.count[2] ),
    .Y(_1681_));
 sky130_fd_sc_hd__and3_1 _4648_ (.A(_1676_),
    .B(_1680_),
    .C(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _4649_ (.A(_1682_),
    .X(\ih.t.next_count[2] ));
 sky130_fd_sc_hd__and4_1 _4650_ (.A(\ih.t.count[0] ),
    .B(\ih.t.count[1] ),
    .C(\ih.t.count[2] ),
    .D(\ih.t.count[3] ),
    .X(_1683_));
 sky130_fd_sc_hd__a31o_1 _4651_ (.A1(\ih.t.count[0] ),
    .A2(\ih.t.count[1] ),
    .A3(\ih.t.count[2] ),
    .B1(\ih.t.count[3] ),
    .X(_1684_));
 sky130_fd_sc_hd__and3b_1 _4652_ (.A_N(_1683_),
    .B(_1684_),
    .C(_1676_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _4653_ (.A(_1685_),
    .X(\ih.t.next_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _4654_ (.A1(\ih.t.count[4] ),
    .A2(_1683_),
    .B1(_1674_),
    .Y(_1686_));
 sky130_fd_sc_hd__a21oi_1 _4655_ (.A1(net220),
    .A2(_1683_),
    .B1(_1686_),
    .Y(\ih.t.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4656_ (.A(\ih.t.count[4] ),
    .B(\ih.t.count[5] ),
    .C(_1683_),
    .X(_1687_));
 sky130_fd_sc_hd__a21o_1 _4657_ (.A1(\ih.t.count[4] ),
    .A2(_1683_),
    .B1(\ih.t.count[5] ),
    .X(_1688_));
 sky130_fd_sc_hd__and3b_1 _4658_ (.A_N(_1687_),
    .B(_1688_),
    .C(_1676_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _4659_ (.A(_1689_),
    .X(\ih.t.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4660_ (.A(\ih.t.count[6] ),
    .B(_1687_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_4 _4661_ (.A(_1673_),
    .X(_1691_));
 sky130_fd_sc_hd__o21ai_1 _4662_ (.A1(net235),
    .A2(_1687_),
    .B1(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(_1690_),
    .B(_1692_),
    .Y(\ih.t.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _4664_ (.A(\ih.t.count[6] ),
    .B(\ih.t.count[7] ),
    .C(_1687_),
    .X(_1693_));
 sky130_fd_sc_hd__o21ai_1 _4665_ (.A1(net223),
    .A2(_1690_),
    .B1(_1691_),
    .Y(_1694_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(_1693_),
    .B(_1694_),
    .Y(\ih.t.next_count[7] ));
 sky130_fd_sc_hd__and2_1 _4667_ (.A(\ih.t.count[8] ),
    .B(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__o21ai_1 _4668_ (.A1(net234),
    .A2(_1693_),
    .B1(_1691_),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_1 _4669_ (.A(_1695_),
    .B(_1696_),
    .Y(\ih.t.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _4670_ (.A(\ih.t.count[8] ),
    .B(\ih.t.count[9] ),
    .C(_1693_),
    .X(_1697_));
 sky130_fd_sc_hd__o21ai_1 _4671_ (.A1(net224),
    .A2(_1695_),
    .B1(_1691_),
    .Y(_1698_));
 sky130_fd_sc_hd__nor2_1 _4672_ (.A(_1697_),
    .B(_1698_),
    .Y(\ih.t.next_count[9] ));
 sky130_fd_sc_hd__o21ai_1 _4673_ (.A1(\ih.t.count[10] ),
    .A2(_1697_),
    .B1(_1674_),
    .Y(_1699_));
 sky130_fd_sc_hd__a21oi_1 _4674_ (.A1(net213),
    .A2(_1697_),
    .B1(_1699_),
    .Y(\ih.t.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4675_ (.A(\ih.t.count[10] ),
    .B(\ih.t.count[11] ),
    .C(_1697_),
    .X(_1700_));
 sky130_fd_sc_hd__a21o_1 _4676_ (.A1(\ih.t.count[10] ),
    .A2(_1697_),
    .B1(\ih.t.count[11] ),
    .X(_1701_));
 sky130_fd_sc_hd__and3b_1 _4677_ (.A_N(_1700_),
    .B(_1701_),
    .C(_1676_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _4678_ (.A(_1702_),
    .X(\ih.t.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4679_ (.A(\ih.t.count[12] ),
    .B(_1700_),
    .X(_1703_));
 sky130_fd_sc_hd__o21ai_1 _4680_ (.A1(\ih.t.count[12] ),
    .A2(_1700_),
    .B1(_1691_),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _4681_ (.A(_1703_),
    .B(_1704_),
    .Y(\ih.t.next_count[12] ));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(\ih.t.count[13] ),
    .A2(_1703_),
    .B1(_1674_),
    .Y(_1705_));
 sky130_fd_sc_hd__a21oi_1 _4683_ (.A1(net218),
    .A2(_1703_),
    .B1(_1705_),
    .Y(\ih.t.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _4684_ (.A(\ih.t.count[13] ),
    .B(\ih.t.count[14] ),
    .C(_1703_),
    .X(_1706_));
 sky130_fd_sc_hd__a31o_1 _4685_ (.A1(\ih.t.count[12] ),
    .A2(\ih.t.count[13] ),
    .A3(_1700_),
    .B1(\ih.t.count[14] ),
    .X(_1707_));
 sky130_fd_sc_hd__and3b_1 _4686_ (.A_N(_1706_),
    .B(_1707_),
    .C(_1676_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _4687_ (.A(_1708_),
    .X(\ih.t.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _4688_ (.A(\ih.t.count[15] ),
    .B(_1706_),
    .X(_1709_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(net232),
    .A2(_1706_),
    .B1(_1691_),
    .Y(_1710_));
 sky130_fd_sc_hd__nor2_1 _4690_ (.A(_1709_),
    .B(_1710_),
    .Y(\ih.t.next_count[15] ));
 sky130_fd_sc_hd__o21ai_1 _4691_ (.A1(\ih.t.count[16] ),
    .A2(_1709_),
    .B1(_1674_),
    .Y(_1711_));
 sky130_fd_sc_hd__a21oi_1 _4692_ (.A1(net212),
    .A2(_1709_),
    .B1(_1711_),
    .Y(\ih.t.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _4693_ (.A(\ih.t.count[16] ),
    .B(\ih.t.count[17] ),
    .C(_1709_),
    .X(_1712_));
 sky130_fd_sc_hd__a31o_1 _4694_ (.A1(\ih.t.count[15] ),
    .A2(\ih.t.count[16] ),
    .A3(_1706_),
    .B1(\ih.t.count[17] ),
    .X(_1713_));
 sky130_fd_sc_hd__and3b_1 _4695_ (.A_N(_1712_),
    .B(_1713_),
    .C(_1676_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _4696_ (.A(_1714_),
    .X(\ih.t.next_count[17] ));
 sky130_fd_sc_hd__and2_1 _4697_ (.A(\ih.t.count[18] ),
    .B(_1712_),
    .X(_1715_));
 sky130_fd_sc_hd__o21ai_1 _4698_ (.A1(net228),
    .A2(_1712_),
    .B1(_1691_),
    .Y(_1716_));
 sky130_fd_sc_hd__nor2_1 _4699_ (.A(_1715_),
    .B(_1716_),
    .Y(\ih.t.next_count[18] ));
 sky130_fd_sc_hd__o21ai_1 _4700_ (.A1(\ih.t.count[19] ),
    .A2(_1715_),
    .B1(_1674_),
    .Y(_1717_));
 sky130_fd_sc_hd__a21oi_1 _4701_ (.A1(net221),
    .A2(_1715_),
    .B1(_1717_),
    .Y(\ih.t.next_count[19] ));
 sky130_fd_sc_hd__and3_1 _4702_ (.A(\ih.t.count[19] ),
    .B(\ih.t.count[20] ),
    .C(_1715_),
    .X(_1718_));
 sky130_fd_sc_hd__a31o_1 _4703_ (.A1(\ih.t.count[18] ),
    .A2(\ih.t.count[19] ),
    .A3(_1712_),
    .B1(\ih.t.count[20] ),
    .X(_1719_));
 sky130_fd_sc_hd__and3b_1 _4704_ (.A_N(_1718_),
    .B(_1719_),
    .C(_1676_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _4705_ (.A(_1720_),
    .X(\ih.t.next_count[20] ));
 sky130_fd_sc_hd__and2_1 _4706_ (.A(\ih.t.count[21] ),
    .B(_1718_),
    .X(_1721_));
 sky130_fd_sc_hd__o21ai_1 _4707_ (.A1(net231),
    .A2(_1718_),
    .B1(_1691_),
    .Y(_1722_));
 sky130_fd_sc_hd__nor2_1 _4708_ (.A(_1721_),
    .B(_1722_),
    .Y(\ih.t.next_count[21] ));
 sky130_fd_sc_hd__o21ai_1 _4709_ (.A1(\ih.t.count[22] ),
    .A2(_1721_),
    .B1(_1674_),
    .Y(_1723_));
 sky130_fd_sc_hd__a21oi_1 _4710_ (.A1(net216),
    .A2(_1721_),
    .B1(_1723_),
    .Y(\ih.t.next_count[22] ));
 sky130_fd_sc_hd__and3_1 _4711_ (.A(\ih.t.count[22] ),
    .B(\ih.t.count[23] ),
    .C(_1721_),
    .X(_1724_));
 sky130_fd_sc_hd__a31o_1 _4712_ (.A1(\ih.t.count[21] ),
    .A2(\ih.t.count[22] ),
    .A3(_1718_),
    .B1(\ih.t.count[23] ),
    .X(_1725_));
 sky130_fd_sc_hd__and3b_1 _4713_ (.A_N(_1724_),
    .B(_1725_),
    .C(_1676_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _4714_ (.A(_1726_),
    .X(\ih.t.next_count[23] ));
 sky130_fd_sc_hd__and2_1 _4715_ (.A(\ih.t.count[24] ),
    .B(_1724_),
    .X(_1727_));
 sky130_fd_sc_hd__o21ai_1 _4716_ (.A1(net229),
    .A2(_1724_),
    .B1(_1691_),
    .Y(_1728_));
 sky130_fd_sc_hd__nor2_1 _4717_ (.A(_1727_),
    .B(_1728_),
    .Y(\ih.t.next_count[24] ));
 sky130_fd_sc_hd__o21ai_1 _4718_ (.A1(\ih.t.count[25] ),
    .A2(_1727_),
    .B1(_1674_),
    .Y(_1729_));
 sky130_fd_sc_hd__a21oi_1 _4719_ (.A1(net217),
    .A2(_1727_),
    .B1(_1729_),
    .Y(\ih.t.next_count[25] ));
 sky130_fd_sc_hd__and3_1 _4720_ (.A(\ih.t.count[25] ),
    .B(\ih.t.count[26] ),
    .C(_1727_),
    .X(_1730_));
 sky130_fd_sc_hd__a31o_1 _4721_ (.A1(\ih.t.count[24] ),
    .A2(\ih.t.count[25] ),
    .A3(_1724_),
    .B1(\ih.t.count[26] ),
    .X(_1731_));
 sky130_fd_sc_hd__and3b_1 _4722_ (.A_N(_1730_),
    .B(_1731_),
    .C(_1673_),
    .X(_1732_));
 sky130_fd_sc_hd__clkbuf_1 _4723_ (.A(_1732_),
    .X(\ih.t.next_count[26] ));
 sky130_fd_sc_hd__and2_1 _4724_ (.A(\ih.t.count[27] ),
    .B(_1730_),
    .X(_1733_));
 sky130_fd_sc_hd__o21ai_1 _4725_ (.A1(net230),
    .A2(_1730_),
    .B1(_1691_),
    .Y(_1734_));
 sky130_fd_sc_hd__nor2_1 _4726_ (.A(_1733_),
    .B(_1734_),
    .Y(\ih.t.next_count[27] ));
 sky130_fd_sc_hd__o21ai_1 _4727_ (.A1(\ih.t.count[28] ),
    .A2(_1733_),
    .B1(_1674_),
    .Y(_1735_));
 sky130_fd_sc_hd__a21oi_1 _4728_ (.A1(net219),
    .A2(_1733_),
    .B1(_1735_),
    .Y(\ih.t.next_count[28] ));
 sky130_fd_sc_hd__and3_1 _4729_ (.A(\ih.t.count[28] ),
    .B(\ih.t.count[29] ),
    .C(_1733_),
    .X(_1736_));
 sky130_fd_sc_hd__a31o_1 _4730_ (.A1(\ih.t.count[27] ),
    .A2(\ih.t.count[28] ),
    .A3(_1730_),
    .B1(\ih.t.count[29] ),
    .X(_1737_));
 sky130_fd_sc_hd__and3b_1 _4731_ (.A_N(_1736_),
    .B(_1737_),
    .C(_1673_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _4732_ (.A(_1738_),
    .X(\ih.t.next_count[29] ));
 sky130_fd_sc_hd__o21ai_1 _4733_ (.A1(net206),
    .A2(_1736_),
    .B1(_1674_),
    .Y(_1739_));
 sky130_fd_sc_hd__a21oi_1 _4734_ (.A1(net206),
    .A2(_1736_),
    .B1(_1739_),
    .Y(\ih.t.next_count[30] ));
 sky130_fd_sc_hd__a21o_1 _4735_ (.A1(\ih.t.count[30] ),
    .A2(_1736_),
    .B1(\ih.t.count[31] ),
    .X(_1740_));
 sky130_fd_sc_hd__nand3_1 _4736_ (.A(\ih.t.count[30] ),
    .B(\ih.t.count[31] ),
    .C(_1736_),
    .Y(_1741_));
 sky130_fd_sc_hd__and3_1 _4737_ (.A(_1676_),
    .B(_1740_),
    .C(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__clkbuf_1 _4738_ (.A(_1742_),
    .X(\ih.t.next_count[31] ));
 sky130_fd_sc_hd__o32a_1 _4739_ (.A1(_2912_),
    .A2(_0361_),
    .A3(_0967_),
    .B1(_0312_),
    .B2(_0324_),
    .X(_1743_));
 sky130_fd_sc_hd__and2b_1 _4740_ (.A_N(_2933_),
    .B(_0302_),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(\cu.alu_f[6] ),
    .A1(\alu.Cin ),
    .S(_0359_),
    .X(_1745_));
 sky130_fd_sc_hd__nor2_1 _4742_ (.A(_0313_),
    .B(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__or4_1 _4743_ (.A(_2911_),
    .B(_0309_),
    .C(_0379_),
    .D(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__o22a_1 _4744_ (.A1(_0336_),
    .A2(_1743_),
    .B1(_1744_),
    .B2(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__or4_1 _4745_ (.A(_0296_),
    .B(_0319_),
    .C(_1317_),
    .D(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__xnor2_1 _4746_ (.A(_2896_),
    .B(_1745_),
    .Y(_1750_));
 sky130_fd_sc_hd__o21ai_1 _4747_ (.A1(_2920_),
    .A2(_2927_),
    .B1(_2881_),
    .Y(_1751_));
 sky130_fd_sc_hd__or3_1 _4748_ (.A(_0302_),
    .B(_0449_),
    .C(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a31o_1 _4749_ (.A1(_2900_),
    .A2(_2923_),
    .A3(_1750_),
    .B1(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__or3b_1 _4750_ (.A(_0301_),
    .B(_1265_),
    .C_N(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__a31o_1 _4751_ (.A1(_0456_),
    .A2(_0457_),
    .A3(_1754_),
    .B1(_0296_),
    .X(_1755_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_1749_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__or3b_1 _4753_ (.A(_1267_),
    .B(_1299_),
    .C_N(_1300_),
    .X(_1757_));
 sky130_fd_sc_hd__or3b_1 _4754_ (.A(net148),
    .B(_0317_),
    .C_N(_0305_),
    .X(_1758_));
 sky130_fd_sc_hd__o31a_1 _4755_ (.A1(_1291_),
    .A2(_1317_),
    .A3(_1758_),
    .B1(_2954_),
    .X(_1759_));
 sky130_fd_sc_hd__or4b_1 _4756_ (.A(_1267_),
    .B(_1300_),
    .C(_1759_),
    .D_N(_1299_),
    .X(_1760_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_1757_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a41o_1 _4758_ (.A1(_2883_),
    .A2(_2916_),
    .A3(_2946_),
    .A4(_0976_),
    .B1(_0297_),
    .X(_1762_));
 sky130_fd_sc_hd__and4bb_1 _4759_ (.A_N(_1762_),
    .B_N(_1300_),
    .C(_2950_),
    .D(_1299_),
    .X(_1763_));
 sky130_fd_sc_hd__a21oi_1 _4760_ (.A1(_2950_),
    .A2(_1300_),
    .B1(_1299_),
    .Y(_1764_));
 sky130_fd_sc_hd__or2_1 _4761_ (.A(_1012_),
    .B(_1755_),
    .X(_1765_));
 sky130_fd_sc_hd__o21ai_1 _4762_ (.A1(_1482_),
    .A2(_1765_),
    .B1(_1749_),
    .Y(_1766_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_0371_),
    .B(_1756_),
    .Y(_1767_));
 sky130_fd_sc_hd__a21oi_1 _4764_ (.A1(_1658_),
    .A2(_1767_),
    .B1(_1482_),
    .Y(_1768_));
 sky130_fd_sc_hd__o22a_1 _4765_ (.A1(_1647_),
    .A2(_1766_),
    .B1(_1768_),
    .B2(_1268_),
    .X(_1769_));
 sky130_fd_sc_hd__o22a_1 _4766_ (.A1(_1299_),
    .A2(_1658_),
    .B1(_1764_),
    .B2(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__a211o_1 _4767_ (.A1(_1756_),
    .A2(_1761_),
    .B1(_1763_),
    .C1(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__or2_1 _4768_ (.A(\cu.id.is_halted ),
    .B(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__clkbuf_1 _4769_ (.A(_1772_),
    .X(_0004_));
 sky130_fd_sc_hd__a31o_1 _4770_ (.A1(_1300_),
    .A2(_1299_),
    .A3(_1765_),
    .B1(_1267_),
    .X(_1773_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_1658_),
    .B(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__o21ai_1 _4772_ (.A1(_1267_),
    .A2(_1755_),
    .B1(_1301_),
    .Y(_1775_));
 sky130_fd_sc_hd__or2b_1 _4773_ (.A(_1760_),
    .B_N(_1755_),
    .X(_1776_));
 sky130_fd_sc_hd__and3b_1 _4774_ (.A_N(_1763_),
    .B(_1775_),
    .C(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__o311a_1 _4775_ (.A1(_1482_),
    .A2(_1634_),
    .A3(_1645_),
    .B1(_1774_),
    .C1(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__nor2_1 _4776_ (.A(net198),
    .B(_1778_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21a_1 _4777_ (.A1(_1299_),
    .A2(_1646_),
    .B1(_1267_),
    .X(_1779_));
 sky130_fd_sc_hd__a21oi_1 _4778_ (.A1(_1299_),
    .A2(_1762_),
    .B1(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__or4b_1 _4779_ (.A(_1267_),
    .B(_1012_),
    .C(_1648_),
    .D_N(_1300_),
    .X(_1781_));
 sky130_fd_sc_hd__o211a_1 _4780_ (.A1(_1300_),
    .A2(_1780_),
    .B1(_1781_),
    .C1(_1302_),
    .X(_1782_));
 sky130_fd_sc_hd__nor2_1 _4781_ (.A(net198),
    .B(_1782_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor2_1 _4782_ (.A(_2708_),
    .B(_1655_),
    .Y(\mc.rw.cmp_check ));
 sky130_fd_sc_hd__nand2_1 _4783_ (.A(_2952_),
    .B(_0986_),
    .Y(_1783_));
 sky130_fd_sc_hd__or4b_1 _4784_ (.A(_0975_),
    .B(_0989_),
    .C(_1783_),
    .D_N(_0994_),
    .X(_1784_));
 sky130_fd_sc_hd__or2_1 _4785_ (.A(_0979_),
    .B(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(net201),
    .B(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__a21boi_1 _4787_ (.A1(_2876_),
    .A2(_1786_),
    .B1_N(net202),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _4788_ (.A(_1778_),
    .B(_1782_),
    .Y(_1787_));
 sky130_fd_sc_hd__o21a_1 _4789_ (.A1(_1771_),
    .A2(_1787_),
    .B1(_0297_),
    .X(_1788_));
 sky130_fd_sc_hd__o21ba_1 _4790_ (.A1(net201),
    .A2(_1788_),
    .B1_N(net203),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _4791_ (.A1(_0297_),
    .A2(_2952_),
    .B1(_1785_),
    .B2(net203),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _4792_ (.A(_0986_),
    .B(_0989_),
    .C(_0994_),
    .X(_1789_));
 sky130_fd_sc_hd__a21oi_1 _4793_ (.A1(_1000_),
    .A2(_1789_),
    .B1(net198),
    .Y(_1790_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(net201),
    .B(_1790_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _4795_ (.A(_1298_),
    .Y(_1791_));
 sky130_fd_sc_hd__xor2_1 _4796_ (.A(_0344_),
    .B(_1298_),
    .X(_1792_));
 sky130_fd_sc_hd__nor2_1 _4797_ (.A(_0292_),
    .B(_0337_),
    .Y(_1793_));
 sky130_fd_sc_hd__nor2_1 _4798_ (.A(_0297_),
    .B(_0358_),
    .Y(_1794_));
 sky130_fd_sc_hd__or2_2 _4799_ (.A(_1794_),
    .B(_0366_),
    .X(_1795_));
 sky130_fd_sc_hd__or4_2 _4800_ (.A(_1185_),
    .B(_1793_),
    .C(_0352_),
    .D(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__clkbuf_4 _4801_ (.A(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__buf_4 _4802_ (.A(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(_0616_),
    .A1(_1791_),
    .S(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__a2bb2o_2 _4804_ (.A1_N(_0986_),
    .A2_N(_1005_),
    .B1(_1789_),
    .B2(_0982_),
    .X(_1800_));
 sky130_fd_sc_hd__nand2_8 _4805_ (.A(_2952_),
    .B(_1800_),
    .Y(_1801_));
 sky130_fd_sc_hd__clkbuf_4 _4806_ (.A(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(_1792_),
    .A1(_1799_),
    .S(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__nor2_1 _4808_ (.A(_0308_),
    .B(_0309_),
    .Y(_1804_));
 sky130_fd_sc_hd__or2_1 _4809_ (.A(_2943_),
    .B(_0328_),
    .X(_1805_));
 sky130_fd_sc_hd__o311a_1 _4810_ (.A1(_2934_),
    .A2(_2902_),
    .A3(_2882_),
    .B1(_0313_),
    .C1(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__or2b_1 _4811_ (.A(_1806_),
    .B_N(_1750_),
    .X(_1807_));
 sky130_fd_sc_hd__o22a_1 _4812_ (.A1(_2920_),
    .A2(_2927_),
    .B1(_2943_),
    .B2(_0329_),
    .X(_1808_));
 sky130_fd_sc_hd__o211a_1 _4813_ (.A1(_0304_),
    .A2(_0303_),
    .B1(_1808_),
    .C1(_2954_),
    .X(_1809_));
 sky130_fd_sc_hd__o2111a_1 _4814_ (.A1(_0359_),
    .A2(_2924_),
    .B1(_1804_),
    .C1(_1807_),
    .D1(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__o21ai_1 _4815_ (.A1(_2946_),
    .A2(_1255_),
    .B1(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__buf_4 _4816_ (.A(net140),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_1791_),
    .A1(_1803_),
    .S(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__o22ai_1 _4818_ (.A1(_1300_),
    .A2(_1778_),
    .B1(_1782_),
    .B2(_1267_),
    .Y(_1814_));
 sky130_fd_sc_hd__xor2_1 _4819_ (.A(_1299_),
    .B(_1771_),
    .X(_1815_));
 sky130_fd_sc_hd__a211o_1 _4820_ (.A1(_1300_),
    .A2(_1778_),
    .B1(_1814_),
    .C1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_4 _4821_ (.A1(_2952_),
    .A2(net140),
    .B1(_1816_),
    .B2(_1483_),
    .X(_1817_));
 sky130_fd_sc_hd__buf_4 _4822_ (.A(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(_1298_),
    .A1(_1813_),
    .S(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _4824_ (.A(_1819_),
    .X(_0016_));
 sky130_fd_sc_hd__xor2_1 _4825_ (.A(_1298_),
    .B(\cu.pc.pc_o[1] ),
    .X(_1820_));
 sky130_fd_sc_hd__xor2_1 _4826_ (.A(_0341_),
    .B(\cu.pc.pc_o[1] ),
    .X(_1821_));
 sky130_fd_sc_hd__and3_1 _4827_ (.A(_0344_),
    .B(_1298_),
    .C(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__a21oi_1 _4828_ (.A1(_0344_),
    .A2(_1298_),
    .B1(_1821_),
    .Y(_1823_));
 sky130_fd_sc_hd__nor2_1 _4829_ (.A(_1822_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(_1048_),
    .A1(_1820_),
    .S(_1798_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(_1824_),
    .A1(_1825_),
    .S(_1802_),
    .X(_1826_));
 sky130_fd_sc_hd__mux2_1 _4832_ (.A0(_1820_),
    .A1(_1826_),
    .S(_1812_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2_1 _4833_ (.A0(\cu.pc.pc_o[1] ),
    .A1(_1827_),
    .S(_1818_),
    .X(_1828_));
 sky130_fd_sc_hd__clkbuf_1 _4834_ (.A(_1828_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _4835_ (.A(_1298_),
    .B(\cu.pc.pc_o[1] ),
    .C(\cu.pc.pc_o[2] ),
    .X(_1829_));
 sky130_fd_sc_hd__a21oi_1 _4836_ (.A1(_1298_),
    .A2(\cu.pc.pc_o[1] ),
    .B1(\cu.pc.pc_o[2] ),
    .Y(_1830_));
 sky130_fd_sc_hd__nor2_1 _4837_ (.A(_1829_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__nor2_1 _4838_ (.A(_0342_),
    .B(\cu.pc.pc_o[2] ),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0342_),
    .B(\cu.pc.pc_o[2] ),
    .Y(_1833_));
 sky130_fd_sc_hd__and2b_1 _4840_ (.A_N(_1832_),
    .B(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__a21oi_1 _4841_ (.A1(_0341_),
    .A2(\cu.pc.pc_o[1] ),
    .B1(_1822_),
    .Y(_1835_));
 sky130_fd_sc_hd__xnor2_1 _4842_ (.A(_1834_),
    .B(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(_1070_),
    .A1(_1831_),
    .S(_1798_),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(_1836_),
    .A1(_1837_),
    .S(_1802_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(_1831_),
    .A1(_1838_),
    .S(_1812_),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _4846_ (.A0(\cu.pc.pc_o[2] ),
    .A1(_1839_),
    .S(_1818_),
    .X(_1840_));
 sky130_fd_sc_hd__clkbuf_1 _4847_ (.A(_1840_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _4848_ (.A(\cu.pc.pc_o[3] ),
    .B(_1829_),
    .X(_1841_));
 sky130_fd_sc_hd__nor2_1 _4849_ (.A(\cu.pc.pc_o[3] ),
    .B(_1829_),
    .Y(_1842_));
 sky130_fd_sc_hd__nor2_1 _4850_ (.A(_1841_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__nor2_1 _4851_ (.A(\cu.id.cb_opcode_y[0] ),
    .B(\cu.pc.pc_o[3] ),
    .Y(_1844_));
 sky130_fd_sc_hd__nand2_1 _4852_ (.A(\cu.id.cb_opcode_y[0] ),
    .B(\cu.pc.pc_o[3] ),
    .Y(_1845_));
 sky130_fd_sc_hd__and2b_1 _4853_ (.A_N(_1844_),
    .B(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__o21a_1 _4854_ (.A1(_1832_),
    .A2(_1835_),
    .B1(_1833_),
    .X(_1847_));
 sky130_fd_sc_hd__xnor2_1 _4855_ (.A(_1846_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__mux2_1 _4856_ (.A0(_1087_),
    .A1(_1843_),
    .S(_1798_),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(_1848_),
    .A1(_1849_),
    .S(_1802_),
    .X(_1850_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(_1843_),
    .A1(_1850_),
    .S(_1812_),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(\cu.pc.pc_o[3] ),
    .A1(_1851_),
    .S(_1818_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _4860_ (.A(_1852_),
    .X(_0019_));
 sky130_fd_sc_hd__xor2_1 _4861_ (.A(\cu.pc.pc_o[4] ),
    .B(_1841_),
    .X(_1853_));
 sky130_fd_sc_hd__nor2_1 _4862_ (.A(_0374_),
    .B(\cu.pc.pc_o[4] ),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_0374_),
    .B(\cu.pc.pc_o[4] ),
    .Y(_1855_));
 sky130_fd_sc_hd__and2b_1 _4864_ (.A_N(_1854_),
    .B(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__o21a_1 _4865_ (.A1(_1844_),
    .A2(_1847_),
    .B1(_1845_),
    .X(_1857_));
 sky130_fd_sc_hd__xnor2_1 _4866_ (.A(_1856_),
    .B(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(_1159_),
    .A1(_1853_),
    .S(_1798_),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(_1858_),
    .A1(_1859_),
    .S(_1802_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_1853_),
    .A1(_1860_),
    .S(_1812_),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(\cu.pc.pc_o[4] ),
    .A1(_1861_),
    .S(_1818_),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _4871_ (.A(_1862_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _4872_ (.A(\cu.pc.pc_o[5] ),
    .B(\cu.pc.pc_o[4] ),
    .C(_1841_),
    .X(_1863_));
 sky130_fd_sc_hd__a21oi_1 _4873_ (.A1(\cu.pc.pc_o[4] ),
    .A2(_1841_),
    .B1(\cu.pc.pc_o[5] ),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _4874_ (.A(_1863_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_1 _4875_ (.A(_0373_),
    .B(\cu.pc.pc_o[5] ),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_0373_),
    .B(\cu.pc.pc_o[5] ),
    .Y(_1867_));
 sky130_fd_sc_hd__and2b_1 _4877_ (.A_N(_1866_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__o21a_1 _4878_ (.A1(_1854_),
    .A2(_1857_),
    .B1(_1855_),
    .X(_1869_));
 sky130_fd_sc_hd__xnor2_1 _4879_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(_1143_),
    .A1(_1865_),
    .S(_1798_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_1 _4881_ (.A0(_1870_),
    .A1(_1871_),
    .S(_1802_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _4882_ (.A0(_1865_),
    .A1(_1872_),
    .S(_1812_),
    .X(_1873_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(\cu.pc.pc_o[5] ),
    .A1(_1873_),
    .S(_1818_),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _4884_ (.A(_1874_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _4885_ (.A(\cu.pc.pc_o[6] ),
    .B(_1863_),
    .X(_1875_));
 sky130_fd_sc_hd__nor2_1 _4886_ (.A(\cu.pc.pc_o[6] ),
    .B(_1863_),
    .Y(_1876_));
 sky130_fd_sc_hd__nor2_1 _4887_ (.A(_1875_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__nor2_1 _4888_ (.A(_0387_),
    .B(\cu.pc.pc_o[6] ),
    .Y(_1878_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_0387_),
    .B(\cu.pc.pc_o[6] ),
    .Y(_1879_));
 sky130_fd_sc_hd__or2b_1 _4890_ (.A(_1878_),
    .B_N(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__o21a_1 _4891_ (.A1(_1866_),
    .A2(_1869_),
    .B1(_1867_),
    .X(_1881_));
 sky130_fd_sc_hd__xor2_1 _4892_ (.A(_1880_),
    .B(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4893_ (.A0(_1125_),
    .A1(_1877_),
    .S(_1798_),
    .X(_1883_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(_1882_),
    .A1(_1883_),
    .S(_1802_),
    .X(_1884_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(_1877_),
    .A1(_1884_),
    .S(_1812_),
    .X(_1885_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(\cu.pc.pc_o[6] ),
    .A1(_1885_),
    .S(_1818_),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _4897_ (.A(_1886_),
    .X(_0022_));
 sky130_fd_sc_hd__xor2_1 _4898_ (.A(\cu.pc.pc_o[7] ),
    .B(_1875_),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_1 _4899_ (.A(_2931_),
    .B(\cu.pc.pc_o[7] ),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(_2931_),
    .B(\cu.pc.pc_o[7] ),
    .Y(_1889_));
 sky130_fd_sc_hd__and2b_1 _4901_ (.A_N(_1888_),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__o21a_1 _4902_ (.A1(_1878_),
    .A2(_1881_),
    .B1(_1879_),
    .X(_1891_));
 sky130_fd_sc_hd__xnor2_1 _4903_ (.A(_1890_),
    .B(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(_1108_),
    .A1(_1887_),
    .S(_1797_),
    .X(_1893_));
 sky130_fd_sc_hd__mux2_1 _4905_ (.A0(_1892_),
    .A1(_1893_),
    .S(_1801_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(_1887_),
    .A1(_1894_),
    .S(_1812_),
    .X(_1895_));
 sky130_fd_sc_hd__mux2_1 _4907_ (.A0(\cu.pc.pc_o[7] ),
    .A1(_1895_),
    .S(_1818_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _4908_ (.A(_1896_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _4909_ (.A(\cu.pc.pc_o[7] ),
    .B(\cu.pc.pc_o[8] ),
    .C(_1875_),
    .X(_1897_));
 sky130_fd_sc_hd__a21oi_1 _4910_ (.A1(\cu.pc.pc_o[7] ),
    .A2(_1875_),
    .B1(\cu.pc.pc_o[8] ),
    .Y(_1898_));
 sky130_fd_sc_hd__nor2_1 _4911_ (.A(_1897_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_1624_),
    .A1(_1899_),
    .S(_1798_),
    .X(_1900_));
 sky130_fd_sc_hd__nor2_1 _4913_ (.A(_2931_),
    .B(\cu.pc.pc_o[8] ),
    .Y(_1901_));
 sky130_fd_sc_hd__and2_1 _4914_ (.A(\cu.id.cb_opcode_x[1] ),
    .B(\cu.pc.pc_o[8] ),
    .X(_1902_));
 sky130_fd_sc_hd__or2_1 _4915_ (.A(_1901_),
    .B(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__o21a_1 _4916_ (.A1(_1888_),
    .A2(_1891_),
    .B1(_1889_),
    .X(_1904_));
 sky130_fd_sc_hd__or2_1 _4917_ (.A(_1903_),
    .B(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__a21oi_1 _4918_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1801_),
    .Y(_1906_));
 sky130_fd_sc_hd__a22o_1 _4919_ (.A1(_1802_),
    .A2(_1900_),
    .B1(_1905_),
    .B2(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_1 _4920_ (.A0(_1899_),
    .A1(_1907_),
    .S(_1812_),
    .X(_1908_));
 sky130_fd_sc_hd__mux2_1 _4921_ (.A0(\cu.pc.pc_o[8] ),
    .A1(_1908_),
    .S(_1818_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _4922_ (.A(_1909_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _4923_ (.A(\cu.pc.pc_o[9] ),
    .B(_1897_),
    .X(_1910_));
 sky130_fd_sc_hd__nor2_1 _4924_ (.A(\cu.pc.pc_o[9] ),
    .B(_1897_),
    .Y(_1911_));
 sky130_fd_sc_hd__nor2_1 _4925_ (.A(_1910_),
    .B(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__xor2_1 _4926_ (.A(_2931_),
    .B(\cu.pc.pc_o[9] ),
    .X(_1913_));
 sky130_fd_sc_hd__or2b_1 _4927_ (.A(_1902_),
    .B_N(_1905_),
    .X(_1914_));
 sky130_fd_sc_hd__xor2_1 _4928_ (.A(_1913_),
    .B(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _4929_ (.A0(_1625_),
    .A1(_1912_),
    .S(_1797_),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_1 _4930_ (.A0(_1915_),
    .A1(_1916_),
    .S(_1801_),
    .X(_1917_));
 sky130_fd_sc_hd__mux2_1 _4931_ (.A0(_1912_),
    .A1(_1917_),
    .S(_1812_),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(\cu.pc.pc_o[9] ),
    .A1(_1918_),
    .S(_1818_),
    .X(_1919_));
 sky130_fd_sc_hd__clkbuf_1 _4933_ (.A(_1919_),
    .X(_0025_));
 sky130_fd_sc_hd__xor2_1 _4934_ (.A(_1522_),
    .B(_1910_),
    .X(_1920_));
 sky130_fd_sc_hd__or2_1 _4935_ (.A(_2931_),
    .B(_1522_),
    .X(_1921_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(_2931_),
    .B(_1522_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_1921_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__o21ai_1 _4938_ (.A1(\cu.pc.pc_o[9] ),
    .A2(\cu.pc.pc_o[8] ),
    .B1(_1232_),
    .Y(_1924_));
 sky130_fd_sc_hd__or2b_1 _4939_ (.A(_1905_),
    .B_N(_1913_),
    .X(_1925_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_1924_),
    .B(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__xnor2_1 _4941_ (.A(_1923_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__mux2_1 _4942_ (.A0(_1225_),
    .A1(_1920_),
    .S(_1797_),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_1 _4943_ (.A0(_1927_),
    .A1(_1928_),
    .S(_1801_),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _4944_ (.A0(_1920_),
    .A1(_1929_),
    .S(net140),
    .X(_1930_));
 sky130_fd_sc_hd__mux2_1 _4945_ (.A0(_1522_),
    .A1(_1930_),
    .S(_1817_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _4946_ (.A(_1931_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _4947_ (.A(\cu.pc.pc_o[11] ),
    .B(_1522_),
    .C(_1910_),
    .X(_1932_));
 sky130_fd_sc_hd__a21oi_1 _4948_ (.A1(_1522_),
    .A2(_1910_),
    .B1(\cu.pc.pc_o[11] ),
    .Y(_1933_));
 sky130_fd_sc_hd__nor2_1 _4949_ (.A(_1932_),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__xnor2_1 _4950_ (.A(_2931_),
    .B(\cu.pc.pc_o[11] ),
    .Y(_1935_));
 sky130_fd_sc_hd__a21bo_1 _4951_ (.A1(_1921_),
    .A2(_1926_),
    .B1_N(_1922_),
    .X(_1936_));
 sky130_fd_sc_hd__xnor2_1 _4952_ (.A(_1935_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(_1221_),
    .A1(_1934_),
    .S(_1797_),
    .X(_1938_));
 sky130_fd_sc_hd__mux2_1 _4954_ (.A0(_1937_),
    .A1(_1938_),
    .S(_1801_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _4955_ (.A0(_1934_),
    .A1(_1939_),
    .S(net140),
    .X(_1940_));
 sky130_fd_sc_hd__mux2_1 _4956_ (.A0(\cu.pc.pc_o[11] ),
    .A1(_1940_),
    .S(_1817_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_1 _4957_ (.A(_1941_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _4958_ (.A(\cu.pc.pc_o[12] ),
    .B(_1932_),
    .X(_1942_));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(\cu.pc.pc_o[12] ),
    .B(_1932_),
    .Y(_1943_));
 sky130_fd_sc_hd__nor2_1 _4960_ (.A(_1942_),
    .B(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__mux2_1 _4961_ (.A0(_1212_),
    .A1(_1944_),
    .S(_1798_),
    .X(_1945_));
 sky130_fd_sc_hd__and2_1 _4962_ (.A(_2931_),
    .B(\cu.pc.pc_o[12] ),
    .X(_1946_));
 sky130_fd_sc_hd__nor2_1 _4963_ (.A(_1232_),
    .B(\cu.pc.pc_o[12] ),
    .Y(_1947_));
 sky130_fd_sc_hd__or2_1 _4964_ (.A(_1946_),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__o21ai_1 _4965_ (.A1(\cu.pc.pc_o[11] ),
    .A2(_1522_),
    .B1(_1232_),
    .Y(_1949_));
 sky130_fd_sc_hd__o311a_1 _4966_ (.A1(_1923_),
    .A2(_1925_),
    .A3(_1935_),
    .B1(_1949_),
    .C1(_1924_),
    .X(_1950_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(_1948_),
    .B(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__a21oi_1 _4968_ (.A1(_1948_),
    .A2(_1950_),
    .B1(_1801_),
    .Y(_1952_));
 sky130_fd_sc_hd__a22o_1 _4969_ (.A1(_1802_),
    .A2(_1945_),
    .B1(_1951_),
    .B2(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(_1944_),
    .A1(_1953_),
    .S(net140),
    .X(_1954_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(\cu.pc.pc_o[12] ),
    .A1(_1954_),
    .S(_1817_),
    .X(_1955_));
 sky130_fd_sc_hd__clkbuf_1 _4972_ (.A(_1955_),
    .X(_0028_));
 sky130_fd_sc_hd__xor2_1 _4973_ (.A(\cu.pc.pc_o[13] ),
    .B(_1942_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _4974_ (.A(_1232_),
    .B(\cu.pc.pc_o[13] ),
    .Y(_1957_));
 sky130_fd_sc_hd__and2_1 _4975_ (.A(_1232_),
    .B(\cu.pc.pc_o[13] ),
    .X(_1958_));
 sky130_fd_sc_hd__nor2_1 _4976_ (.A(_1957_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__and2b_1 _4977_ (.A_N(_1946_),
    .B(_1951_),
    .X(_1960_));
 sky130_fd_sc_hd__xnor2_1 _4978_ (.A(_1959_),
    .B(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__mux2_1 _4979_ (.A0(_1208_),
    .A1(_1956_),
    .S(_1797_),
    .X(_1962_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(_1961_),
    .A1(_1962_),
    .S(_1801_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _4981_ (.A0(_1956_),
    .A1(_1963_),
    .S(net140),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _4982_ (.A0(\cu.pc.pc_o[13] ),
    .A1(_1964_),
    .S(_1817_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_1 _4983_ (.A(_1965_),
    .X(_0029_));
 sky130_fd_sc_hd__and3_1 _4984_ (.A(\cu.pc.pc_o[14] ),
    .B(\cu.pc.pc_o[13] ),
    .C(_1942_),
    .X(_1966_));
 sky130_fd_sc_hd__a21oi_1 _4985_ (.A1(\cu.pc.pc_o[13] ),
    .A2(_1942_),
    .B1(\cu.pc.pc_o[14] ),
    .Y(_1967_));
 sky130_fd_sc_hd__nor2_1 _4986_ (.A(_1966_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__xor2_1 _4987_ (.A(_1232_),
    .B(\cu.pc.pc_o[14] ),
    .X(_1969_));
 sky130_fd_sc_hd__and2b_1 _4988_ (.A_N(_1951_),
    .B(_1959_),
    .X(_1970_));
 sky130_fd_sc_hd__or3_1 _4989_ (.A(_1946_),
    .B(_1958_),
    .C(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__and2_1 _4990_ (.A(_1969_),
    .B(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__o21bai_1 _4991_ (.A1(_1969_),
    .A2(_1971_),
    .B1_N(_1801_),
    .Y(_1973_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_1626_),
    .A1(_1968_),
    .S(_1798_),
    .X(_1974_));
 sky130_fd_sc_hd__a2bb2o_1 _4993_ (.A1_N(_1972_),
    .A2_N(_1973_),
    .B1(_1974_),
    .B2(_1802_),
    .X(_1975_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_1968_),
    .A1(_1975_),
    .S(net140),
    .X(_1976_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(\cu.pc.pc_o[14] ),
    .A1(_1976_),
    .S(_1817_),
    .X(_1977_));
 sky130_fd_sc_hd__clkbuf_1 _4996_ (.A(_1977_),
    .X(_0030_));
 sky130_fd_sc_hd__xor2_1 _4997_ (.A(\cu.pc.pc_o[15] ),
    .B(_1966_),
    .X(_1978_));
 sky130_fd_sc_hd__o21a_1 _4998_ (.A1(\cu.pc.pc_o[14] ),
    .A2(_1971_),
    .B1(_1232_),
    .X(_1979_));
 sky130_fd_sc_hd__o21ba_1 _4999_ (.A1(_1232_),
    .A2(_1972_),
    .B1_N(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__xor2_1 _5000_ (.A(\cu.pc.pc_o[15] ),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(_1262_),
    .A1(_1978_),
    .S(_1797_),
    .X(_1982_));
 sky130_fd_sc_hd__mux2_1 _5002_ (.A0(_1981_),
    .A1(_1982_),
    .S(_1801_),
    .X(_1983_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(_1978_),
    .A1(_1983_),
    .S(net140),
    .X(_1984_));
 sky130_fd_sc_hd__mux2_1 _5004_ (.A0(\cu.pc.pc_o[15] ),
    .A1(_1984_),
    .S(_1817_),
    .X(_1985_));
 sky130_fd_sc_hd__clkbuf_1 _5005_ (.A(_1985_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(_0617_),
    .A1(_1624_),
    .S(_0368_),
    .X(_1986_));
 sky130_fd_sc_hd__and3_1 _5007_ (.A(_2955_),
    .B(_0367_),
    .C(_0352_),
    .X(_1987_));
 sky130_fd_sc_hd__buf_4 _5008_ (.A(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__mux2_1 _5009_ (.A0(\cu.reg_file.reg_a[0] ),
    .A1(_1986_),
    .S(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__clkbuf_1 _5010_ (.A(_1989_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(_1049_),
    .A1(_1625_),
    .S(_0368_),
    .X(_1990_));
 sky130_fd_sc_hd__mux2_1 _5012_ (.A0(\cu.reg_file.reg_a[1] ),
    .A1(_1990_),
    .S(_1988_),
    .X(_1991_));
 sky130_fd_sc_hd__clkbuf_1 _5013_ (.A(_1991_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(_1071_),
    .A1(_1225_),
    .S(_0368_),
    .X(_1992_));
 sky130_fd_sc_hd__mux2_1 _5015_ (.A0(\cu.reg_file.reg_a[2] ),
    .A1(_1992_),
    .S(_1988_),
    .X(_1993_));
 sky130_fd_sc_hd__clkbuf_1 _5016_ (.A(_1993_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(_1186_),
    .A1(_1221_),
    .S(_0368_),
    .X(_1994_));
 sky130_fd_sc_hd__mux2_1 _5018_ (.A0(\cu.reg_file.reg_a[3] ),
    .A1(_1994_),
    .S(_1988_),
    .X(_1995_));
 sky130_fd_sc_hd__clkbuf_1 _5019_ (.A(_1995_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(_1188_),
    .A1(_1212_),
    .S(_0368_),
    .X(_1996_));
 sky130_fd_sc_hd__mux2_1 _5021_ (.A0(\cu.reg_file.reg_a[4] ),
    .A1(_1996_),
    .S(_1988_),
    .X(_1997_));
 sky130_fd_sc_hd__clkbuf_1 _5022_ (.A(_1997_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _5023_ (.A0(_1190_),
    .A1(_1208_),
    .S(_0368_),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_1 _5024_ (.A0(\cu.reg_file.reg_a[5] ),
    .A1(_1998_),
    .S(_1988_),
    .X(_1999_));
 sky130_fd_sc_hd__clkbuf_1 _5025_ (.A(_1999_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _5026_ (.A0(_1192_),
    .A1(_1626_),
    .S(_0368_),
    .X(_2000_));
 sky130_fd_sc_hd__mux2_1 _5027_ (.A0(\cu.reg_file.reg_a[6] ),
    .A1(_2000_),
    .S(_1988_),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_1 _5028_ (.A(_2001_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(_1259_),
    .A1(_1262_),
    .S(_0368_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(\cu.reg_file.reg_a[7] ),
    .A1(_2002_),
    .S(_1988_),
    .X(_2003_));
 sky130_fd_sc_hd__clkbuf_1 _5031_ (.A(_2003_),
    .X(_0039_));
 sky130_fd_sc_hd__and4b_1 _5032_ (.A_N(_1793_),
    .B(_0352_),
    .C(_1794_),
    .D(_0366_),
    .X(_2004_));
 sky130_fd_sc_hd__buf_4 _5033_ (.A(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _5034_ (.A0(_0617_),
    .A1(_1624_),
    .S(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_1793_),
    .B(_0352_),
    .Y(_2007_));
 sky130_fd_sc_hd__nor2_1 _5036_ (.A(_1795_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__o21a_4 _5037_ (.A1(_2005_),
    .A2(_2008_),
    .B1(_2955_),
    .X(_2009_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(\cu.reg_file.reg_b[0] ),
    .A1(_2006_),
    .S(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _5039_ (.A(_2010_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _5040_ (.A0(_1049_),
    .A1(_1625_),
    .S(_2005_),
    .X(_2011_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(\cu.reg_file.reg_b[1] ),
    .A1(_2011_),
    .S(_2009_),
    .X(_2012_));
 sky130_fd_sc_hd__clkbuf_1 _5042_ (.A(_2012_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(_1071_),
    .A1(_1225_),
    .S(_2005_),
    .X(_2013_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(\cu.reg_file.reg_b[2] ),
    .A1(_2013_),
    .S(_2009_),
    .X(_2014_));
 sky130_fd_sc_hd__clkbuf_1 _5045_ (.A(_2014_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(_1186_),
    .A1(_1221_),
    .S(_2005_),
    .X(_2015_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(\cu.reg_file.reg_b[3] ),
    .A1(_2015_),
    .S(_2009_),
    .X(_2016_));
 sky130_fd_sc_hd__clkbuf_1 _5048_ (.A(_2016_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(_1188_),
    .A1(_1212_),
    .S(_2005_),
    .X(_2017_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(\cu.reg_file.reg_b[4] ),
    .A1(_2017_),
    .S(_2009_),
    .X(_2018_));
 sky130_fd_sc_hd__clkbuf_1 _5051_ (.A(_2018_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _5052_ (.A0(_1190_),
    .A1(_1208_),
    .S(_2005_),
    .X(_2019_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(\cu.reg_file.reg_b[5] ),
    .A1(_2019_),
    .S(_2009_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_1 _5054_ (.A(_2020_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(_1192_),
    .A1(_1626_),
    .S(_2005_),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(\cu.reg_file.reg_b[6] ),
    .A1(_2021_),
    .S(_2009_),
    .X(_2022_));
 sky130_fd_sc_hd__clkbuf_1 _5057_ (.A(_2022_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(_1259_),
    .A1(_1262_),
    .S(_2005_),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_1 _5059_ (.A0(\cu.reg_file.reg_b[7] ),
    .A1(_2023_),
    .S(_2009_),
    .X(_2024_));
 sky130_fd_sc_hd__clkbuf_1 _5060_ (.A(_2024_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _5061_ (.A(_0617_),
    .X(_2025_));
 sky130_fd_sc_hd__or3_2 _5062_ (.A(_0297_),
    .B(_0358_),
    .C(_0366_),
    .X(_2026_));
 sky130_fd_sc_hd__nor2_1 _5063_ (.A(_2007_),
    .B(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__o21a_4 _5064_ (.A1(_2005_),
    .A2(_2027_),
    .B1(_2955_),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _5065_ (.A0(\cu.reg_file.reg_c[0] ),
    .A1(_2025_),
    .S(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _5066_ (.A(_2029_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(\cu.reg_file.reg_c[1] ),
    .A1(_1049_),
    .S(_2028_),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _5068_ (.A(_2030_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(\cu.reg_file.reg_c[2] ),
    .A1(_1071_),
    .S(_2028_),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _5070_ (.A(_2031_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(\cu.reg_file.reg_c[3] ),
    .A1(_1186_),
    .S(_2028_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _5072_ (.A(_2032_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(\cu.reg_file.reg_c[4] ),
    .A1(_1188_),
    .S(_2028_),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_1 _5074_ (.A(_2033_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _5075_ (.A0(\cu.reg_file.reg_c[5] ),
    .A1(_1190_),
    .S(_2028_),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _5076_ (.A(_2034_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _5077_ (.A0(\cu.reg_file.reg_c[6] ),
    .A1(_1192_),
    .S(_2028_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _5078_ (.A(_2035_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _5079_ (.A0(\cu.reg_file.reg_c[7] ),
    .A1(_1259_),
    .S(_2028_),
    .X(_2036_));
 sky130_fd_sc_hd__clkbuf_1 _5080_ (.A(_2036_),
    .X(_0055_));
 sky130_fd_sc_hd__o21ai_2 _5081_ (.A1(_0292_),
    .A2(_0337_),
    .B1(_0352_),
    .Y(_2037_));
 sky130_fd_sc_hd__nor2_4 _5082_ (.A(_2037_),
    .B(_1795_),
    .Y(_2038_));
 sky130_fd_sc_hd__mux2_1 _5083_ (.A0(_0616_),
    .A1(_1624_),
    .S(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__and2b_1 _5084_ (.A_N(_0352_),
    .B(_1793_),
    .X(_2040_));
 sky130_fd_sc_hd__a21o_1 _5085_ (.A1(_0367_),
    .A2(_2040_),
    .B1(_2038_),
    .X(_2041_));
 sky130_fd_sc_hd__and2_1 _5086_ (.A(_2955_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__buf_4 _5087_ (.A(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _5088_ (.A0(\cu.reg_file.reg_d[0] ),
    .A1(_2039_),
    .S(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _5089_ (.A(_2044_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _5090_ (.A0(_1049_),
    .A1(_1625_),
    .S(_2038_),
    .X(_2045_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(\cu.reg_file.reg_d[1] ),
    .A1(_2045_),
    .S(_2043_),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _5092_ (.A(_2046_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(_1071_),
    .A1(_1225_),
    .S(_2038_),
    .X(_2047_));
 sky130_fd_sc_hd__mux2_1 _5094_ (.A0(\cu.reg_file.reg_d[2] ),
    .A1(_2047_),
    .S(_2043_),
    .X(_2048_));
 sky130_fd_sc_hd__clkbuf_1 _5095_ (.A(_2048_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(_1186_),
    .A1(_1221_),
    .S(_2038_),
    .X(_2049_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(\cu.reg_file.reg_d[3] ),
    .A1(_2049_),
    .S(_2043_),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _5098_ (.A(_2050_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(_1188_),
    .A1(_1212_),
    .S(_2038_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _5100_ (.A0(\cu.reg_file.reg_d[4] ),
    .A1(_2051_),
    .S(_2043_),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _5101_ (.A(_2052_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _5102_ (.A0(_1190_),
    .A1(_1208_),
    .S(_2038_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _5103_ (.A0(\cu.reg_file.reg_d[5] ),
    .A1(_2053_),
    .S(_2043_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _5104_ (.A(_2054_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(_1192_),
    .A1(_1626_),
    .S(_2038_),
    .X(_2055_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(\cu.reg_file.reg_d[6] ),
    .A1(_2055_),
    .S(_2043_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _5107_ (.A(_2056_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(_1108_),
    .A1(_1262_),
    .S(_2038_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(\cu.reg_file.reg_d[7] ),
    .A1(_2057_),
    .S(_2043_),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _5110_ (.A(_2058_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_2 _5111_ (.A(_0617_),
    .X(_2059_));
 sky130_fd_sc_hd__a31o_1 _5112_ (.A1(_1794_),
    .A2(_0366_),
    .A3(_2040_),
    .B1(_2038_),
    .X(_2060_));
 sky130_fd_sc_hd__and2_1 _5113_ (.A(_2955_),
    .B(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_4 _5114_ (.A(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(\cu.reg_file.reg_e[0] ),
    .A1(_2059_),
    .S(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _5116_ (.A(_2063_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(\cu.reg_file.reg_e[1] ),
    .A1(_1049_),
    .S(_2062_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _5118_ (.A(_2064_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _5119_ (.A0(\cu.reg_file.reg_e[2] ),
    .A1(_1071_),
    .S(_2062_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _5120_ (.A(_2065_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(\cu.reg_file.reg_e[3] ),
    .A1(_1186_),
    .S(_2062_),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _5122_ (.A(_2066_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(\cu.reg_file.reg_e[4] ),
    .A1(_1188_),
    .S(_2062_),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_1 _5124_ (.A(_2067_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _5125_ (.A0(\cu.reg_file.reg_e[5] ),
    .A1(_1190_),
    .S(_2062_),
    .X(_2068_));
 sky130_fd_sc_hd__clkbuf_1 _5126_ (.A(_2068_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(\cu.reg_file.reg_e[6] ),
    .A1(_1192_),
    .S(_2062_),
    .X(_2069_));
 sky130_fd_sc_hd__clkbuf_1 _5128_ (.A(_2069_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(\cu.reg_file.reg_e[7] ),
    .A1(_1259_),
    .S(_2062_),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _5130_ (.A(_2070_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _5131_ (.A(_2037_),
    .B(_2026_),
    .X(_2071_));
 sky130_fd_sc_hd__buf_4 _5132_ (.A(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(_1624_),
    .A1(_0616_),
    .S(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__or3b_1 _5134_ (.A(_0352_),
    .B(_1795_),
    .C_N(_1793_),
    .X(_2074_));
 sky130_fd_sc_hd__a21bo_4 _5135_ (.A1(_2072_),
    .A2(_2074_),
    .B1_N(_2955_),
    .X(_2075_));
 sky130_fd_sc_hd__mux2_1 _5136_ (.A0(_2073_),
    .A1(\cu.reg_file.reg_h[0] ),
    .S(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__clkbuf_1 _5137_ (.A(_2076_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _5138_ (.A0(_1625_),
    .A1(_1048_),
    .S(_2072_),
    .X(_2077_));
 sky130_fd_sc_hd__mux2_1 _5139_ (.A0(_2077_),
    .A1(\cu.reg_file.reg_h[1] ),
    .S(_2075_),
    .X(_2078_));
 sky130_fd_sc_hd__clkbuf_1 _5140_ (.A(_2078_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(_1225_),
    .A1(_1070_),
    .S(_2072_),
    .X(_2079_));
 sky130_fd_sc_hd__mux2_1 _5142_ (.A0(_2079_),
    .A1(\cu.reg_file.reg_h[2] ),
    .S(_2075_),
    .X(_2080_));
 sky130_fd_sc_hd__clkbuf_1 _5143_ (.A(_2080_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(_1221_),
    .A1(_1087_),
    .S(_2072_),
    .X(_2081_));
 sky130_fd_sc_hd__mux2_1 _5145_ (.A0(_2081_),
    .A1(\cu.reg_file.reg_h[3] ),
    .S(_2075_),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _5146_ (.A(_2082_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(_1212_),
    .A1(_1159_),
    .S(_2072_),
    .X(_2083_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(_2083_),
    .A1(\cu.reg_file.reg_h[4] ),
    .S(_2075_),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_1 _5149_ (.A(_2084_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _5150_ (.A0(_1208_),
    .A1(_1143_),
    .S(_2072_),
    .X(_2085_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(_2085_),
    .A1(\cu.reg_file.reg_h[5] ),
    .S(_2075_),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _5152_ (.A(_2086_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(_1626_),
    .A1(_1125_),
    .S(_2072_),
    .X(_2087_));
 sky130_fd_sc_hd__mux2_1 _5154_ (.A0(_2087_),
    .A1(\cu.reg_file.reg_h[6] ),
    .S(_2075_),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_1 _5155_ (.A(_2088_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(_1262_),
    .A1(_1108_),
    .S(_2072_),
    .X(_2089_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(_2089_),
    .A1(\cu.reg_file.reg_h[7] ),
    .S(_2075_),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_1 _5158_ (.A(_2090_),
    .X(_0079_));
 sky130_fd_sc_hd__inv_2 _5159_ (.A(_2026_),
    .Y(_2091_));
 sky130_fd_sc_hd__and3_1 _5160_ (.A(_2955_),
    .B(_2007_),
    .C(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__clkbuf_4 _5161_ (.A(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__mux2_1 _5162_ (.A0(\cu.reg_file.reg_l[0] ),
    .A1(_2059_),
    .S(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__clkbuf_1 _5163_ (.A(_2094_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _5164_ (.A0(\cu.reg_file.reg_l[1] ),
    .A1(_1049_),
    .S(_2093_),
    .X(_2095_));
 sky130_fd_sc_hd__clkbuf_1 _5165_ (.A(_2095_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _5166_ (.A0(\cu.reg_file.reg_l[2] ),
    .A1(_1071_),
    .S(_2093_),
    .X(_2096_));
 sky130_fd_sc_hd__clkbuf_1 _5167_ (.A(_2096_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(\cu.reg_file.reg_l[3] ),
    .A1(_1186_),
    .S(_2093_),
    .X(_2097_));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(_2097_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _5170_ (.A0(\cu.reg_file.reg_l[4] ),
    .A1(_1188_),
    .S(_2093_),
    .X(_2098_));
 sky130_fd_sc_hd__clkbuf_1 _5171_ (.A(_2098_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(\cu.reg_file.reg_l[5] ),
    .A1(_1190_),
    .S(_2093_),
    .X(_2099_));
 sky130_fd_sc_hd__clkbuf_1 _5173_ (.A(_2099_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(\cu.reg_file.reg_l[6] ),
    .A1(_1192_),
    .S(_2093_),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_1 _5175_ (.A(_2100_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(\cu.reg_file.reg_l[7] ),
    .A1(_1259_),
    .S(_2093_),
    .X(_2101_));
 sky130_fd_sc_hd__clkbuf_1 _5177_ (.A(_2101_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _5178_ (.A0(\mc.cl.next_data[8] ),
    .A1(net18),
    .S(\mc.count ),
    .X(_2102_));
 sky130_fd_sc_hd__and2_1 _5179_ (.A(_1649_),
    .B(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(_2103_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(\mc.cl.next_data[9] ),
    .A1(net19),
    .S(\mc.count ),
    .X(_2104_));
 sky130_fd_sc_hd__and2_1 _5182_ (.A(_1649_),
    .B(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__clkbuf_1 _5183_ (.A(_2105_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _5184_ (.A0(\mc.cl.next_data[10] ),
    .A1(net20),
    .S(\mc.count ),
    .X(_2106_));
 sky130_fd_sc_hd__and2_1 _5185_ (.A(_1649_),
    .B(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__clkbuf_1 _5186_ (.A(_2107_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(\mc.cl.next_data[11] ),
    .A1(net21),
    .S(\mc.count ),
    .X(_2108_));
 sky130_fd_sc_hd__and2_1 _5188_ (.A(_1649_),
    .B(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__clkbuf_1 _5189_ (.A(_2109_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(\mc.cl.next_data[12] ),
    .A1(net22),
    .S(\mc.count ),
    .X(_2110_));
 sky130_fd_sc_hd__and2_1 _5191_ (.A(_1649_),
    .B(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__clkbuf_1 _5192_ (.A(_2111_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(\mc.cl.next_data[13] ),
    .A1(net23),
    .S(\mc.count ),
    .X(_2112_));
 sky130_fd_sc_hd__and2_1 _5194_ (.A(_1649_),
    .B(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_1 _5195_ (.A(_2113_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _5196_ (.A0(\mc.cl.next_data[14] ),
    .A1(net24),
    .S(\mc.count ),
    .X(_2114_));
 sky130_fd_sc_hd__and2_1 _5197_ (.A(_1649_),
    .B(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _5198_ (.A(_2115_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(\mc.cl.next_data[15] ),
    .A1(net25),
    .S(\mc.count ),
    .X(_2116_));
 sky130_fd_sc_hd__and2_1 _5200_ (.A(_1649_),
    .B(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _5201_ (.A(_2117_),
    .X(_0095_));
 sky130_fd_sc_hd__or3b_1 _5202_ (.A(_1793_),
    .B(_0352_),
    .C_N(_2955_),
    .X(_2118_));
 sky130_fd_sc_hd__clkbuf_4 _5203_ (.A(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__inv_2 _5204_ (.A(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__mux2_1 _5205_ (.A0(\cu.reg_file.reg_sp[0] ),
    .A1(_2059_),
    .S(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__clkbuf_1 _5206_ (.A(_2121_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_4 _5207_ (.A(_1636_),
    .X(_2122_));
 sky130_fd_sc_hd__or2_1 _5208_ (.A(_1364_),
    .B(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__buf_2 _5209_ (.A(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(_0618_),
    .A1(\ih.gpio_interrupt_mask[0] ),
    .S(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_1 _5211_ (.A(_2125_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(_1050_),
    .A1(\ih.gpio_interrupt_mask[1] ),
    .S(_2124_),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_1 _5213_ (.A(_2126_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(_1072_),
    .A1(\ih.gpio_interrupt_mask[2] ),
    .S(_2124_),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_1 _5215_ (.A(_2127_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(_1187_),
    .A1(\ih.gpio_interrupt_mask[3] ),
    .S(_2124_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _5217_ (.A(_2128_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(_1189_),
    .A1(\ih.gpio_interrupt_mask[4] ),
    .S(_2124_),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _5219_ (.A(_2129_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(_1191_),
    .A1(\ih.gpio_interrupt_mask[5] ),
    .S(_2124_),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _5221_ (.A(_2130_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(_1193_),
    .A1(\ih.gpio_interrupt_mask[6] ),
    .S(_2124_),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(_2131_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(_1260_),
    .A1(\ih.gpio_interrupt_mask[7] ),
    .S(_2124_),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _5225_ (.A(_2132_),
    .X(_0104_));
 sky130_fd_sc_hd__a211o_1 _5226_ (.A1(_1374_),
    .A2(_1627_),
    .B1(_1632_),
    .C1(_1414_),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_4 _5227_ (.A(_1638_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_4 _5228_ (.A(_1416_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__and2_1 _5229_ (.A(_1357_),
    .B(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__buf_2 _5230_ (.A(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__or3_2 _5231_ (.A(_1367_),
    .B(_1627_),
    .C(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__or3_1 _5232_ (.A(_1364_),
    .B(_2133_),
    .C(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(_0618_),
    .A1(\ih.t.enable ),
    .S(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_1 _5234_ (.A(_2140_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(_0616_),
    .A1(_1624_),
    .S(_1671_),
    .X(_2141_));
 sky130_fd_sc_hd__nor2_1 _5236_ (.A(_1369_),
    .B(_1627_),
    .Y(_2142_));
 sky130_fd_sc_hd__clkbuf_4 _5237_ (.A(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_8 _5238_ (.A(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__or2_2 _5239_ (.A(_1327_),
    .B(_1372_),
    .X(_2145_));
 sky130_fd_sc_hd__nor2_1 _5240_ (.A(_1374_),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__or2_2 _5241_ (.A(_2142_),
    .B(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_4 _5242_ (.A(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__o211a_1 _5243_ (.A1(_1665_),
    .A2(_2148_),
    .B1(_1357_),
    .C1(_1633_),
    .X(_2149_));
 sky130_fd_sc_hd__o21a_4 _5244_ (.A1(_1671_),
    .A2(_2144_),
    .B1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(\ih.t.timer_max[24] ),
    .A1(_2141_),
    .S(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__clkbuf_1 _5246_ (.A(_2151_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(_1048_),
    .A1(_1625_),
    .S(_1671_),
    .X(_2152_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(\ih.t.timer_max[25] ),
    .A1(_2152_),
    .S(_2150_),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_1 _5249_ (.A(_2153_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5250_ (.A0(_1070_),
    .A1(_1225_),
    .S(_1671_),
    .X(_2154_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(\ih.t.timer_max[26] ),
    .A1(_2154_),
    .S(_2150_),
    .X(_2155_));
 sky130_fd_sc_hd__clkbuf_1 _5252_ (.A(_2155_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(_1087_),
    .A1(_1221_),
    .S(_1671_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(\ih.t.timer_max[27] ),
    .A1(_2156_),
    .S(_2150_),
    .X(_2157_));
 sky130_fd_sc_hd__clkbuf_1 _5255_ (.A(_2157_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(_1159_),
    .A1(_1212_),
    .S(_1671_),
    .X(_2158_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(\ih.t.timer_max[28] ),
    .A1(_2158_),
    .S(_2150_),
    .X(_2159_));
 sky130_fd_sc_hd__clkbuf_1 _5258_ (.A(_2159_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5259_ (.A0(_1143_),
    .A1(_1208_),
    .S(_1670_),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(\ih.t.timer_max[29] ),
    .A1(_2160_),
    .S(_2150_),
    .X(_2161_));
 sky130_fd_sc_hd__clkbuf_1 _5261_ (.A(_2161_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(_1125_),
    .A1(_1626_),
    .S(_1670_),
    .X(_2162_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(\ih.t.timer_max[30] ),
    .A1(_2162_),
    .S(_2150_),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_1 _5264_ (.A(_2163_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(_1108_),
    .A1(_1262_),
    .S(_1670_),
    .X(_2164_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(\ih.t.timer_max[31] ),
    .A1(_2164_),
    .S(_2150_),
    .X(_2165_));
 sky130_fd_sc_hd__clkbuf_1 _5267_ (.A(_2165_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_8 _5268_ (.A(_1644_),
    .X(_2166_));
 sky130_fd_sc_hd__nor2_8 _5269_ (.A(_2166_),
    .B(_2138_),
    .Y(_2167_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(net76),
    .A1(_2059_),
    .S(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_1 _5271_ (.A(_2168_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net77),
    .A1(_1049_),
    .S(_2167_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _5273_ (.A(_2169_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(net78),
    .A1(_1071_),
    .S(_2167_),
    .X(_2170_));
 sky130_fd_sc_hd__clkbuf_1 _5275_ (.A(_2170_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(net79),
    .A1(_1186_),
    .S(_2167_),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_1 _5277_ (.A(_2171_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(net80),
    .A1(_1188_),
    .S(_2167_),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _5279_ (.A(_2172_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(net81),
    .A1(_1190_),
    .S(_2167_),
    .X(_2173_));
 sky130_fd_sc_hd__clkbuf_1 _5281_ (.A(_2173_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(net82),
    .A1(_1192_),
    .S(_2167_),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _5283_ (.A(_2174_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net83),
    .A1(_1259_),
    .S(_2167_),
    .X(_2175_));
 sky130_fd_sc_hd__clkbuf_1 _5285_ (.A(_2175_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_2 _5286_ (.A(_1327_),
    .B(_1354_),
    .Y(_2176_));
 sky130_fd_sc_hd__and2_4 _5287_ (.A(_1369_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nor2_8 _5288_ (.A(_1364_),
    .B(_2166_),
    .Y(_2178_));
 sky130_fd_sc_hd__nand2_8 _5289_ (.A(_2177_),
    .B(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(_0618_),
    .A1(net84),
    .S(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__clkbuf_1 _5291_ (.A(_2180_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(_1050_),
    .A1(net85),
    .S(_2179_),
    .X(_2181_));
 sky130_fd_sc_hd__clkbuf_1 _5293_ (.A(_2181_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(_1072_),
    .A1(net86),
    .S(_2179_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_1 _5295_ (.A(_2182_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(_1187_),
    .A1(net87),
    .S(_2179_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _5297_ (.A(_2183_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(_1189_),
    .A1(net88),
    .S(_2179_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_1 _5299_ (.A(_2184_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(_1191_),
    .A1(net89),
    .S(_2179_),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _5301_ (.A(_2185_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(_1193_),
    .A1(net90),
    .S(_2179_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _5303_ (.A(_2186_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(_1260_),
    .A1(net91),
    .S(_2179_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_1 _5305_ (.A(_2187_),
    .X(_0129_));
 sky130_fd_sc_hd__nand2_2 _5306_ (.A(_1327_),
    .B(_1354_),
    .Y(_2188_));
 sky130_fd_sc_hd__nor2_1 _5307_ (.A(_1374_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__clkbuf_4 _5308_ (.A(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_8 _5309_ (.A(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__nand2_8 _5310_ (.A(_2178_),
    .B(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(_0618_),
    .A1(net92),
    .S(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_1 _5312_ (.A(_2193_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(_1050_),
    .A1(net93),
    .S(_2192_),
    .X(_2194_));
 sky130_fd_sc_hd__clkbuf_1 _5314_ (.A(_2194_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(_1072_),
    .A1(net94),
    .S(_2192_),
    .X(_2195_));
 sky130_fd_sc_hd__clkbuf_1 _5316_ (.A(_2195_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _5317_ (.A0(_1187_),
    .A1(net95),
    .S(_2192_),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _5318_ (.A(_2196_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(_1189_),
    .A1(net96),
    .S(_2192_),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _5320_ (.A(_2197_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(_1191_),
    .A1(net97),
    .S(_2192_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _5322_ (.A(_2198_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(_1193_),
    .A1(net98),
    .S(_2192_),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _5324_ (.A(_2199_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(_1260_),
    .A1(net99),
    .S(_2192_),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _5326_ (.A(_2200_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_4 _5327_ (.A(_2146_),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_8 _5328_ (.A(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__nand2_8 _5329_ (.A(_2202_),
    .B(_2178_),
    .Y(_2203_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(_0618_),
    .A1(net100),
    .S(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _5331_ (.A(_2204_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(_1050_),
    .A1(net101),
    .S(_2203_),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_1 _5333_ (.A(_2205_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(_1072_),
    .A1(net102),
    .S(_2203_),
    .X(_2206_));
 sky130_fd_sc_hd__clkbuf_1 _5335_ (.A(_2206_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(_1187_),
    .A1(net103),
    .S(_2203_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_1 _5337_ (.A(_2207_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(_1189_),
    .A1(net104),
    .S(_2203_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_1 _5339_ (.A(_2208_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5340_ (.A0(_1191_),
    .A1(net105),
    .S(_2203_),
    .X(_2209_));
 sky130_fd_sc_hd__clkbuf_1 _5341_ (.A(_2209_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(_1193_),
    .A1(net106),
    .S(_2203_),
    .X(_2210_));
 sky130_fd_sc_hd__clkbuf_1 _5343_ (.A(_2210_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(_1260_),
    .A1(net107),
    .S(_2203_),
    .X(_2211_));
 sky130_fd_sc_hd__clkbuf_1 _5345_ (.A(_2211_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_8 _5346_ (.A(_2144_),
    .B(_2178_),
    .Y(_2212_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(_0618_),
    .A1(net108),
    .S(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__clkbuf_1 _5348_ (.A(_2213_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(_1050_),
    .A1(net109),
    .S(_2212_),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_1 _5350_ (.A(_2214_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(_1072_),
    .A1(net110),
    .S(_2212_),
    .X(_2215_));
 sky130_fd_sc_hd__clkbuf_1 _5352_ (.A(_2215_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(_1187_),
    .A1(net111),
    .S(_2212_),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_1 _5354_ (.A(_2216_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(_1189_),
    .A1(net112),
    .S(_2212_),
    .X(_2217_));
 sky130_fd_sc_hd__clkbuf_1 _5356_ (.A(_2217_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(_1191_),
    .A1(net113),
    .S(_2212_),
    .X(_2218_));
 sky130_fd_sc_hd__clkbuf_1 _5358_ (.A(_2218_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(_1193_),
    .A1(net114),
    .S(_2212_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _5360_ (.A(_2219_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(_1260_),
    .A1(net115),
    .S(_2212_),
    .X(_2220_));
 sky130_fd_sc_hd__clkbuf_1 _5362_ (.A(_2220_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(_1374_),
    .B(_2176_),
    .X(_2221_));
 sky130_fd_sc_hd__buf_4 _5364_ (.A(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__nand2_4 _5365_ (.A(_2178_),
    .B(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(_0618_),
    .A1(net116),
    .S(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__clkbuf_1 _5367_ (.A(_2224_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(_1050_),
    .A1(net117),
    .S(_2223_),
    .X(_2225_));
 sky130_fd_sc_hd__clkbuf_1 _5369_ (.A(_2225_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(_1072_),
    .A1(net118),
    .S(_2223_),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_1 _5371_ (.A(_2226_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(_1187_),
    .A1(net119),
    .S(_2223_),
    .X(_2227_));
 sky130_fd_sc_hd__clkbuf_1 _5373_ (.A(_2227_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(_1189_),
    .A1(net120),
    .S(_2223_),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_1 _5375_ (.A(_2228_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(_1191_),
    .A1(net121),
    .S(_2223_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_1 _5377_ (.A(_2229_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(_1193_),
    .A1(net122),
    .S(_2223_),
    .X(_2230_));
 sky130_fd_sc_hd__clkbuf_1 _5379_ (.A(_2230_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(_1260_),
    .A1(net123),
    .S(_2223_),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_1 _5381_ (.A(_2231_),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _5382_ (.A(_1369_),
    .B(_2188_),
    .Y(_2232_));
 sky130_fd_sc_hd__clkbuf_8 _5383_ (.A(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__nand2_8 _5384_ (.A(_2178_),
    .B(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(_0618_),
    .A1(net124),
    .S(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_2235_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(_1050_),
    .A1(net125),
    .S(_2234_),
    .X(_2236_));
 sky130_fd_sc_hd__clkbuf_1 _5388_ (.A(_2236_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(_1072_),
    .A1(net126),
    .S(_2234_),
    .X(_2237_));
 sky130_fd_sc_hd__clkbuf_1 _5390_ (.A(_2237_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(_1187_),
    .A1(net127),
    .S(_2234_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _5392_ (.A(_2238_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(_1189_),
    .A1(net128),
    .S(_2234_),
    .X(_2239_));
 sky130_fd_sc_hd__clkbuf_1 _5394_ (.A(_2239_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(_1191_),
    .A1(net129),
    .S(_2234_),
    .X(_2240_));
 sky130_fd_sc_hd__clkbuf_1 _5396_ (.A(_2240_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(_1193_),
    .A1(net130),
    .S(_2234_),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_1 _5398_ (.A(_2241_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(_1260_),
    .A1(net131),
    .S(_2234_),
    .X(_2242_));
 sky130_fd_sc_hd__clkbuf_1 _5400_ (.A(_2242_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _5401_ (.A(_1369_),
    .B(_2145_),
    .Y(_2243_));
 sky130_fd_sc_hd__buf_4 _5402_ (.A(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__nand2_4 _5403_ (.A(_2178_),
    .B(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(_2025_),
    .A1(net132),
    .S(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__clkbuf_1 _5405_ (.A(_2246_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(_1050_),
    .A1(net133),
    .S(_2245_),
    .X(_2247_));
 sky130_fd_sc_hd__clkbuf_1 _5407_ (.A(_2247_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(_1072_),
    .A1(net134),
    .S(_2245_),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_1 _5409_ (.A(_2248_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(_1187_),
    .A1(net135),
    .S(_2245_),
    .X(_2249_));
 sky130_fd_sc_hd__clkbuf_1 _5411_ (.A(_2249_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5412_ (.A0(_1189_),
    .A1(net136),
    .S(_2245_),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_1 _5413_ (.A(_2250_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(_1191_),
    .A1(net137),
    .S(_2245_),
    .X(_2251_));
 sky130_fd_sc_hd__clkbuf_1 _5415_ (.A(_2251_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(_1193_),
    .A1(net138),
    .S(_2245_),
    .X(_2252_));
 sky130_fd_sc_hd__clkbuf_1 _5417_ (.A(_2252_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(_1260_),
    .A1(net139),
    .S(_2245_),
    .X(_2253_));
 sky130_fd_sc_hd__clkbuf_1 _5419_ (.A(_2253_),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _5420_ (.A(_1327_),
    .B(_1372_),
    .C(_1369_),
    .X(_2254_));
 sky130_fd_sc_hd__and3_1 _5421_ (.A(_1357_),
    .B(_2254_),
    .C(_2135_),
    .X(_2255_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(net68),
    .A1(_2059_),
    .S(_2255_),
    .X(_2256_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(_2256_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_2137_),
    .B(_2177_),
    .Y(_2257_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(_2025_),
    .A1(net69),
    .S(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__clkbuf_1 _5426_ (.A(_2258_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_2137_),
    .B(_2191_),
    .Y(_2259_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(_2025_),
    .A1(net70),
    .S(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__clkbuf_1 _5429_ (.A(_2260_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_2137_),
    .B(_2202_),
    .Y(_2261_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(_2025_),
    .A1(net71),
    .S(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_1 _5432_ (.A(_2262_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _5433_ (.A(_2137_),
    .B(_2144_),
    .Y(_2263_));
 sky130_fd_sc_hd__mux2_1 _5434_ (.A0(_2025_),
    .A1(net72),
    .S(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__clkbuf_1 _5435_ (.A(_2264_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_2137_),
    .B(_2222_),
    .Y(_2265_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(_2025_),
    .A1(net73),
    .S(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__clkbuf_1 _5438_ (.A(_2266_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _5439_ (.A(_2137_),
    .B(_2233_),
    .Y(_2267_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_2025_),
    .A1(net74),
    .S(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2268_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_2137_),
    .B(_2244_),
    .Y(_2269_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(_2025_),
    .A1(net75),
    .S(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__clkbuf_1 _5444_ (.A(_2270_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_2 _5445_ (.A(_1642_),
    .X(_2271_));
 sky130_fd_sc_hd__or2_1 _5446_ (.A(_1414_),
    .B(_2134_),
    .X(_2272_));
 sky130_fd_sc_hd__mux4_1 _5447_ (.A0(net73),
    .A1(net75),
    .A2(net72),
    .A3(net74),
    .S0(_1354_),
    .S1(_1335_),
    .X(_2273_));
 sky130_fd_sc_hd__nor2_1 _5448_ (.A(_1328_),
    .B(_1354_),
    .Y(_2274_));
 sky130_fd_sc_hd__a22o_1 _5449_ (.A1(net68),
    .A2(_2274_),
    .B1(_2176_),
    .B2(net69),
    .X(_2275_));
 sky130_fd_sc_hd__nor2_2 _5450_ (.A(_1328_),
    .B(_1372_),
    .Y(_2276_));
 sky130_fd_sc_hd__a22o_1 _5451_ (.A1(net71),
    .A2(_1640_),
    .B1(_2276_),
    .B2(net70),
    .X(_2277_));
 sky130_fd_sc_hd__or3_1 _5452_ (.A(_1374_),
    .B(_2275_),
    .C(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__o21ai_1 _5453_ (.A1(_1369_),
    .A2(_2273_),
    .B1(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__or4_1 _5454_ (.A(_1364_),
    .B(_2271_),
    .C(_2272_),
    .D(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__buf_2 _5455_ (.A(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__nor2_1 _5456_ (.A(_1635_),
    .B(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__mux2_1 _5457_ (.A0(net60),
    .A1(_2059_),
    .S(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _5458_ (.A(_2283_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_1369_),
    .B(_2176_),
    .Y(_2284_));
 sky130_fd_sc_hd__nor2_1 _5460_ (.A(_2284_),
    .B(_2281_),
    .Y(_2285_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(net61),
    .A1(_2059_),
    .S(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _5462_ (.A(_2286_),
    .X(_0187_));
 sky130_fd_sc_hd__inv_2 _5463_ (.A(_2191_),
    .Y(_2287_));
 sky130_fd_sc_hd__nor2_1 _5464_ (.A(_2287_),
    .B(_2281_),
    .Y(_2288_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(net62),
    .A1(_2059_),
    .S(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__clkbuf_1 _5466_ (.A(_2289_),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _5467_ (.A(_2202_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _5468_ (.A(_2290_),
    .B(_2281_),
    .Y(_2291_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net63),
    .A1(_2059_),
    .S(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _5470_ (.A(_2292_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _5471_ (.A(_2144_),
    .Y(_2293_));
 sky130_fd_sc_hd__nor2_1 _5472_ (.A(_2293_),
    .B(_2281_),
    .Y(_2294_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(net64),
    .A1(_2059_),
    .S(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(_2295_),
    .X(_0190_));
 sky130_fd_sc_hd__inv_2 _5475_ (.A(_2222_),
    .Y(_2296_));
 sky130_fd_sc_hd__nor2_1 _5476_ (.A(_2296_),
    .B(_2281_),
    .Y(_2297_));
 sky130_fd_sc_hd__mux2_1 _5477_ (.A0(net65),
    .A1(_0617_),
    .S(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _5478_ (.A(_2298_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _5479_ (.A(_2233_),
    .Y(_2299_));
 sky130_fd_sc_hd__nor2_1 _5480_ (.A(_2299_),
    .B(_2281_),
    .Y(_2300_));
 sky130_fd_sc_hd__mux2_1 _5481_ (.A0(net66),
    .A1(_0617_),
    .S(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5482_ (.A(_2301_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _5483_ (.A(_2244_),
    .Y(_2302_));
 sky130_fd_sc_hd__nor2_1 _5484_ (.A(_2302_),
    .B(_2281_),
    .Y(_2303_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(net67),
    .A1(_0617_),
    .S(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__clkbuf_1 _5486_ (.A(_2304_),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _5487_ (.A1(net84),
    .A2(_2177_),
    .B1(_2221_),
    .B2(net116),
    .X(_2305_));
 sky130_fd_sc_hd__a221o_1 _5488_ (.A1(net124),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net132),
    .C1(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__a22o_1 _5489_ (.A1(net108),
    .A2(_2143_),
    .B1(_2190_),
    .B2(net92),
    .X(_2307_));
 sky130_fd_sc_hd__a211o_1 _5490_ (.A1(net100),
    .A2(_2202_),
    .B1(_2307_),
    .C1(_2254_),
    .X(_2308_));
 sky130_fd_sc_hd__o22a_1 _5491_ (.A1(net76),
    .A2(_1635_),
    .B1(_2306_),
    .B2(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__and3_2 _5492_ (.A(\mc.cl.cmp_o ),
    .B(_1650_),
    .C(_2133_),
    .X(_2310_));
 sky130_fd_sc_hd__nor2_2 _5493_ (.A(_1399_),
    .B(_2284_),
    .Y(_2311_));
 sky130_fd_sc_hd__a22o_1 _5494_ (.A1(\ih.t.enable ),
    .A2(_2254_),
    .B1(_2189_),
    .B2(\ih.t.timer_max[8] ),
    .X(_2312_));
 sky130_fd_sc_hd__a22o_1 _5495_ (.A1(\ih.t.timer_max[24] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[16] ),
    .X(_2313_));
 sky130_fd_sc_hd__nor2_1 _5496_ (.A(_2312_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__o2bb2a_1 _5497_ (.A1_N(\ih.t.timer_max[0] ),
    .A2_N(_2311_),
    .B1(_2314_),
    .B2(_1399_),
    .X(_2315_));
 sky130_fd_sc_hd__or2_2 _5498_ (.A(_2177_),
    .B(_2190_),
    .X(_2316_));
 sky130_fd_sc_hd__clkbuf_4 _5499_ (.A(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__a221o_1 _5500_ (.A1(\ih.t.enable ),
    .A2(_2254_),
    .B1(_2147_),
    .B2(\ih.t.timer_max[16] ),
    .C1(_1664_),
    .X(_2318_));
 sky130_fd_sc_hd__a21oi_1 _5501_ (.A1(\ih.t.timer_max[0] ),
    .A2(_2317_),
    .B1(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__a21oi_1 _5502_ (.A1(_1665_),
    .A2(_2315_),
    .B1(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__a2111oi_4 _5503_ (.A1(_1374_),
    .A2(_1627_),
    .B1(_1632_),
    .C1(_1488_),
    .D1(_1414_),
    .Y(_2321_));
 sky130_fd_sc_hd__a22o_1 _5504_ (.A1(\mc.cl.next_data[0] ),
    .A2(_2310_),
    .B1(_2320_),
    .B2(net141),
    .X(_2322_));
 sky130_fd_sc_hd__nor2_2 _5505_ (.A(_1488_),
    .B(_2122_),
    .Y(_2323_));
 sky130_fd_sc_hd__nor3_4 _5506_ (.A(_1416_),
    .B(_1631_),
    .C(_1639_),
    .Y(_2324_));
 sky130_fd_sc_hd__a221o_1 _5507_ (.A1(_2122_),
    .A2(_2322_),
    .B1(_2323_),
    .B2(\ih.gpio_interrupt_mask[0] ),
    .C1(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__o211a_1 _5508_ (.A1(_2166_),
    .A2(_2309_),
    .B1(_2325_),
    .C1(_2134_),
    .X(_2326_));
 sky130_fd_sc_hd__a31o_1 _5509_ (.A1(net68),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2327_));
 sky130_fd_sc_hd__a22o_1 _5510_ (.A1(net64),
    .A2(_2274_),
    .B1(_2176_),
    .B2(net65),
    .X(_2328_));
 sky130_fd_sc_hd__a22o_1 _5511_ (.A1(net67),
    .A2(_1640_),
    .B1(_2276_),
    .B2(net66),
    .X(_2329_));
 sky130_fd_sc_hd__a22o_1 _5512_ (.A1(net60),
    .A2(_2274_),
    .B1(_2176_),
    .B2(net61),
    .X(_2330_));
 sky130_fd_sc_hd__a22o_1 _5513_ (.A1(net63),
    .A2(_1640_),
    .B1(_2276_),
    .B2(net62),
    .X(_2331_));
 sky130_fd_sc_hd__or3_1 _5514_ (.A(_1374_),
    .B(_2330_),
    .C(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__o31a_1 _5515_ (.A1(_1369_),
    .A2(_2328_),
    .A3(_2329_),
    .B1(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__or3_1 _5516_ (.A(net32),
    .B(_1335_),
    .C(_1354_),
    .X(_2334_));
 sky130_fd_sc_hd__o21a_1 _5517_ (.A1(net33),
    .A2(_2188_),
    .B1(_1374_),
    .X(_2335_));
 sky130_fd_sc_hd__o22a_1 _5518_ (.A1(net31),
    .A2(_1627_),
    .B1(_2145_),
    .B2(net34),
    .X(_2336_));
 sky130_fd_sc_hd__mux4_1 _5519_ (.A0(net28),
    .A1(net30),
    .A2(net27),
    .A3(net29),
    .S0(_1354_),
    .S1(_1335_),
    .X(_2337_));
 sky130_fd_sc_hd__a32o_1 _5520_ (.A1(_2334_),
    .A2(_2335_),
    .A3(_2336_),
    .B1(_2337_),
    .B2(_1369_),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(_2333_),
    .A1(_2338_),
    .S(_2279_),
    .X(_2339_));
 sky130_fd_sc_hd__and3b_1 _5522_ (.A_N(_2272_),
    .B(_2339_),
    .C(_1650_),
    .X(_2340_));
 sky130_fd_sc_hd__nand2_2 _5523_ (.A(_1670_),
    .B(_2188_),
    .Y(_2341_));
 sky130_fd_sc_hd__nand2_2 _5524_ (.A(_1627_),
    .B(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__a22o_1 _5525_ (.A1(net16),
    .A2(_2176_),
    .B1(_2276_),
    .B2(\ih.input_handler_enable ),
    .X(_2343_));
 sky130_fd_sc_hd__a21o_1 _5526_ (.A1(net2),
    .A2(_2342_),
    .B1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(net2),
    .A1(_2145_),
    .S(_2341_),
    .X(_2345_));
 sky130_fd_sc_hd__a31o_1 _5528_ (.A1(_1651_),
    .A2(_2344_),
    .A3(_2345_),
    .B1(_1643_),
    .X(_2346_));
 sky130_fd_sc_hd__o31a_2 _5529_ (.A1(_2326_),
    .A2(_2327_),
    .A3(_2340_),
    .B1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(\cu.reg_file.reg_mem[0] ),
    .A1(_2347_),
    .S(_1659_),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_1 _5531_ (.A(_2348_),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _5532_ (.A1(net125),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net133),
    .X(_2349_));
 sky130_fd_sc_hd__a21o_1 _5533_ (.A1(net93),
    .A2(_2191_),
    .B1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__or2_1 _5534_ (.A(net85),
    .B(_1335_),
    .X(_2351_));
 sky130_fd_sc_hd__a22o_1 _5535_ (.A1(net101),
    .A2(_2202_),
    .B1(_2351_),
    .B2(_1400_),
    .X(_2352_));
 sky130_fd_sc_hd__a221o_1 _5536_ (.A1(net109),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net117),
    .C1(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__o22a_1 _5537_ (.A1(net77),
    .A2(_1635_),
    .B1(_2350_),
    .B2(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__buf_2 _5538_ (.A(_2310_),
    .X(_2355_));
 sky130_fd_sc_hd__a22o_1 _5539_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[17] ),
    .X(_2356_));
 sky130_fd_sc_hd__a221o_1 _5540_ (.A1(\ih.t.timer_max[9] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[1] ),
    .C1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__and2b_1 _5541_ (.A_N(_1399_),
    .B(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__a221o_1 _5542_ (.A1(\ih.t.timer_max[17] ),
    .A2(_2148_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[1] ),
    .C1(_1665_),
    .X(_2359_));
 sky130_fd_sc_hd__o21a_1 _5543_ (.A1(_1670_),
    .A2(_2358_),
    .B1(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__a22o_1 _5544_ (.A1(\mc.cl.next_data[1] ),
    .A2(_2355_),
    .B1(net141),
    .B2(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__a221o_1 _5545_ (.A1(\ih.gpio_interrupt_mask[1] ),
    .A2(_2323_),
    .B1(_2361_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2362_));
 sky130_fd_sc_hd__o211a_1 _5546_ (.A1(_2166_),
    .A2(_2354_),
    .B1(_2362_),
    .C1(_2134_),
    .X(_2363_));
 sky130_fd_sc_hd__a31o_1 _5547_ (.A1(net69),
    .A2(_1651_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2364_));
 sky130_fd_sc_hd__and3_2 _5548_ (.A(_1328_),
    .B(_1372_),
    .C(_1665_),
    .X(_2365_));
 sky130_fd_sc_hd__a22o_1 _5549_ (.A1(net9),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net17),
    .X(_2366_));
 sky130_fd_sc_hd__and2_1 _5550_ (.A(_1651_),
    .B(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__o22a_2 _5551_ (.A1(_2363_),
    .A2(_2364_),
    .B1(_2367_),
    .B2(_1643_),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(\cu.reg_file.reg_mem[1] ),
    .A1(_2368_),
    .S(_1659_),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _5553_ (.A(_2369_),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _5554_ (.A1(net126),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net134),
    .X(_2370_));
 sky130_fd_sc_hd__a21o_1 _5555_ (.A1(net94),
    .A2(_2191_),
    .B1(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__or2_1 _5556_ (.A(net86),
    .B(_1335_),
    .X(_2372_));
 sky130_fd_sc_hd__a22o_1 _5557_ (.A1(net102),
    .A2(_2202_),
    .B1(_2372_),
    .B2(_1400_),
    .X(_2373_));
 sky130_fd_sc_hd__a221o_1 _5558_ (.A1(net110),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net118),
    .C1(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__o22a_1 _5559_ (.A1(net78),
    .A2(_1635_),
    .B1(_2371_),
    .B2(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__a22o_1 _5560_ (.A1(\ih.t.timer_max[26] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[18] ),
    .X(_2376_));
 sky130_fd_sc_hd__a221o_1 _5561_ (.A1(\ih.t.timer_max[10] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[2] ),
    .C1(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__and2b_1 _5562_ (.A_N(_1399_),
    .B(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__a221o_1 _5563_ (.A1(\ih.t.timer_max[18] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[2] ),
    .C1(_1665_),
    .X(_2379_));
 sky130_fd_sc_hd__o21a_1 _5564_ (.A1(_1670_),
    .A2(_2378_),
    .B1(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__a22o_1 _5565_ (.A1(\mc.cl.next_data[2] ),
    .A2(_2355_),
    .B1(net141),
    .B2(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__a221o_1 _5566_ (.A1(\ih.gpio_interrupt_mask[2] ),
    .A2(_2323_),
    .B1(_2381_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2382_));
 sky130_fd_sc_hd__o211a_1 _5567_ (.A1(_2166_),
    .A2(_2375_),
    .B1(_2382_),
    .C1(_2134_),
    .X(_2383_));
 sky130_fd_sc_hd__a31o_1 _5568_ (.A1(net70),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2384_));
 sky130_fd_sc_hd__a22o_1 _5569_ (.A1(net10),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net3),
    .X(_2385_));
 sky130_fd_sc_hd__and2_1 _5570_ (.A(_1651_),
    .B(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__o22a_2 _5571_ (.A1(_2383_),
    .A2(_2384_),
    .B1(_2386_),
    .B2(_1643_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(\cu.reg_file.reg_mem[2] ),
    .A1(_2387_),
    .S(_1659_),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _5573_ (.A(_2388_),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _5574_ (.A1(net127),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net135),
    .X(_2389_));
 sky130_fd_sc_hd__a21o_1 _5575_ (.A1(net95),
    .A2(_2191_),
    .B1(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__or2_1 _5576_ (.A(net87),
    .B(_1335_),
    .X(_2391_));
 sky130_fd_sc_hd__a22o_1 _5577_ (.A1(net103),
    .A2(_2202_),
    .B1(_2391_),
    .B2(_1400_),
    .X(_2392_));
 sky130_fd_sc_hd__a221o_1 _5578_ (.A1(net111),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net119),
    .C1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__o22a_1 _5579_ (.A1(net79),
    .A2(_1635_),
    .B1(_2390_),
    .B2(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__a22o_1 _5580_ (.A1(\ih.t.timer_max[27] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[19] ),
    .X(_2395_));
 sky130_fd_sc_hd__a221o_1 _5581_ (.A1(\ih.t.timer_max[11] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[3] ),
    .C1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__and2b_1 _5582_ (.A_N(_1399_),
    .B(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__a221o_1 _5583_ (.A1(\ih.t.timer_max[19] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[3] ),
    .C1(_1665_),
    .X(_2398_));
 sky130_fd_sc_hd__o21a_1 _5584_ (.A1(_1670_),
    .A2(_2397_),
    .B1(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__a22o_1 _5585_ (.A1(\mc.cl.next_data[3] ),
    .A2(_2310_),
    .B1(_2321_),
    .B2(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__a221o_1 _5586_ (.A1(\ih.gpio_interrupt_mask[3] ),
    .A2(_2323_),
    .B1(_2400_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2401_));
 sky130_fd_sc_hd__o211a_1 _5587_ (.A1(_2166_),
    .A2(_2394_),
    .B1(_2401_),
    .C1(_2134_),
    .X(_2402_));
 sky130_fd_sc_hd__a31o_1 _5588_ (.A1(net71),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2403_));
 sky130_fd_sc_hd__a22o_1 _5589_ (.A1(net11),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net4),
    .X(_2404_));
 sky130_fd_sc_hd__and2_1 _5590_ (.A(_1651_),
    .B(_2404_),
    .X(_2405_));
 sky130_fd_sc_hd__o22a_2 _5591_ (.A1(_2402_),
    .A2(_2403_),
    .B1(_2405_),
    .B2(_1643_),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(\cu.reg_file.reg_mem[3] ),
    .A1(_2406_),
    .S(_1659_),
    .X(_2407_));
 sky130_fd_sc_hd__clkbuf_1 _5593_ (.A(_2407_),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _5594_ (.A1(net128),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net136),
    .X(_2408_));
 sky130_fd_sc_hd__a21o_1 _5595_ (.A1(net96),
    .A2(_2191_),
    .B1(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__or2_1 _5596_ (.A(net88),
    .B(_1335_),
    .X(_2410_));
 sky130_fd_sc_hd__a22o_1 _5597_ (.A1(net104),
    .A2(_2202_),
    .B1(_2410_),
    .B2(_1400_),
    .X(_2411_));
 sky130_fd_sc_hd__a221o_1 _5598_ (.A1(net112),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net120),
    .C1(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__o22a_1 _5599_ (.A1(net80),
    .A2(_1635_),
    .B1(_2409_),
    .B2(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__a22o_1 _5600_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[20] ),
    .X(_2414_));
 sky130_fd_sc_hd__a221o_1 _5601_ (.A1(\ih.t.timer_max[12] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[4] ),
    .C1(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__and2b_1 _5602_ (.A_N(_1399_),
    .B(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__a221o_1 _5603_ (.A1(\ih.t.timer_max[20] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[4] ),
    .C1(_1665_),
    .X(_2417_));
 sky130_fd_sc_hd__o21a_1 _5604_ (.A1(_1670_),
    .A2(_2416_),
    .B1(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__a22o_1 _5605_ (.A1(\mc.cl.next_data[4] ),
    .A2(_2310_),
    .B1(_2321_),
    .B2(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__a221o_1 _5606_ (.A1(\ih.gpio_interrupt_mask[4] ),
    .A2(_2323_),
    .B1(_2419_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2420_));
 sky130_fd_sc_hd__o211a_1 _5607_ (.A1(_2166_),
    .A2(_2413_),
    .B1(_2420_),
    .C1(_2134_),
    .X(_2421_));
 sky130_fd_sc_hd__a31o_1 _5608_ (.A1(net72),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2422_));
 sky130_fd_sc_hd__a22o_1 _5609_ (.A1(net12),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net5),
    .X(_2423_));
 sky130_fd_sc_hd__and2_1 _5610_ (.A(_1651_),
    .B(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__o22a_2 _5611_ (.A1(_2421_),
    .A2(_2422_),
    .B1(_2424_),
    .B2(_1643_),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(\cu.reg_file.reg_mem[4] ),
    .A1(_2425_),
    .S(_1659_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5613_ (.A(_2426_),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_1 _5614_ (.A1(net129),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net137),
    .X(_2427_));
 sky130_fd_sc_hd__a21o_1 _5615_ (.A1(net97),
    .A2(_2191_),
    .B1(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__or2_1 _5616_ (.A(net89),
    .B(_1335_),
    .X(_2429_));
 sky130_fd_sc_hd__a22o_1 _5617_ (.A1(net105),
    .A2(_2202_),
    .B1(_2429_),
    .B2(_1400_),
    .X(_2430_));
 sky130_fd_sc_hd__a221o_1 _5618_ (.A1(net113),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net121),
    .C1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__o22a_1 _5619_ (.A1(net81),
    .A2(_1635_),
    .B1(_2428_),
    .B2(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__a22o_1 _5620_ (.A1(\ih.t.timer_max[29] ),
    .A2(_2143_),
    .B1(_2201_),
    .B2(\ih.t.timer_max[21] ),
    .X(_2433_));
 sky130_fd_sc_hd__a221o_1 _5621_ (.A1(\ih.t.timer_max[13] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[5] ),
    .C1(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__and2b_1 _5622_ (.A_N(_1399_),
    .B(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__a221o_1 _5623_ (.A1(\ih.t.timer_max[21] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[5] ),
    .C1(_1665_),
    .X(_2436_));
 sky130_fd_sc_hd__o21a_1 _5624_ (.A1(_1670_),
    .A2(_2435_),
    .B1(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__a22o_1 _5625_ (.A1(\mc.cl.next_data[5] ),
    .A2(_2310_),
    .B1(net141),
    .B2(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__a221o_1 _5626_ (.A1(\ih.gpio_interrupt_mask[5] ),
    .A2(_2323_),
    .B1(_2438_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2439_));
 sky130_fd_sc_hd__o211a_1 _5627_ (.A1(_2166_),
    .A2(_2432_),
    .B1(_2439_),
    .C1(_2134_),
    .X(_2440_));
 sky130_fd_sc_hd__a31o_1 _5628_ (.A1(net73),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2441_));
 sky130_fd_sc_hd__a22o_1 _5629_ (.A1(net13),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net6),
    .X(_2442_));
 sky130_fd_sc_hd__and2_1 _5630_ (.A(_1651_),
    .B(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__o22a_2 _5631_ (.A1(_2440_),
    .A2(_2441_),
    .B1(_2443_),
    .B2(_1643_),
    .X(_2444_));
 sky130_fd_sc_hd__mux2_1 _5632_ (.A0(\cu.reg_file.reg_mem[5] ),
    .A1(_2444_),
    .S(_1659_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_1 _5633_ (.A(_2445_),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _5634_ (.A1(net130),
    .A2(_2233_),
    .B1(_2244_),
    .B2(net138),
    .X(_2446_));
 sky130_fd_sc_hd__a21o_1 _5635_ (.A1(net98),
    .A2(_2191_),
    .B1(_2446_),
    .X(_2447_));
 sky130_fd_sc_hd__or2_1 _5636_ (.A(net90),
    .B(_1335_),
    .X(_2448_));
 sky130_fd_sc_hd__a22o_1 _5637_ (.A1(net106),
    .A2(_2201_),
    .B1(_2448_),
    .B2(_1400_),
    .X(_2449_));
 sky130_fd_sc_hd__a221o_1 _5638_ (.A1(net114),
    .A2(_2144_),
    .B1(_2222_),
    .B2(net122),
    .C1(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__o22a_1 _5639_ (.A1(net82),
    .A2(_1635_),
    .B1(_2447_),
    .B2(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__a22o_1 _5640_ (.A1(\ih.t.timer_max[30] ),
    .A2(_2143_),
    .B1(_2146_),
    .B2(\ih.t.timer_max[22] ),
    .X(_2452_));
 sky130_fd_sc_hd__a221o_1 _5641_ (.A1(\ih.t.timer_max[14] ),
    .A2(_2190_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[6] ),
    .C1(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__and2b_1 _5642_ (.A_N(_1399_),
    .B(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__a221o_1 _5643_ (.A1(\ih.t.timer_max[22] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[6] ),
    .C1(_1664_),
    .X(_2455_));
 sky130_fd_sc_hd__o21a_1 _5644_ (.A1(_1669_),
    .A2(_2454_),
    .B1(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__a22o_1 _5645_ (.A1(\mc.cl.next_data[6] ),
    .A2(_2310_),
    .B1(_2321_),
    .B2(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__a221o_1 _5646_ (.A1(\ih.gpio_interrupt_mask[6] ),
    .A2(_2323_),
    .B1(_2457_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2458_));
 sky130_fd_sc_hd__o211a_1 _5647_ (.A1(_2166_),
    .A2(_2451_),
    .B1(_2458_),
    .C1(_2134_),
    .X(_2459_));
 sky130_fd_sc_hd__a31o_1 _5648_ (.A1(net74),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2460_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(net14),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net7),
    .X(_2461_));
 sky130_fd_sc_hd__and2_1 _5650_ (.A(_1651_),
    .B(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__o22a_2 _5651_ (.A1(_2459_),
    .A2(_2460_),
    .B1(_2462_),
    .B2(_1643_),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _5652_ (.A0(\cu.reg_file.reg_mem[6] ),
    .A1(_2463_),
    .S(_1658_),
    .X(_2464_));
 sky130_fd_sc_hd__clkbuf_1 _5653_ (.A(_2464_),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _5654_ (.A1(net131),
    .A2(_2232_),
    .B1(_2243_),
    .B2(net139),
    .X(_2465_));
 sky130_fd_sc_hd__a21o_1 _5655_ (.A1(net99),
    .A2(_2190_),
    .B1(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__or2_1 _5656_ (.A(net91),
    .B(_1327_),
    .X(_2467_));
 sky130_fd_sc_hd__a22o_1 _5657_ (.A1(net107),
    .A2(_2201_),
    .B1(_2467_),
    .B2(_1400_),
    .X(_2468_));
 sky130_fd_sc_hd__a221o_1 _5658_ (.A1(net115),
    .A2(_2143_),
    .B1(_2222_),
    .B2(net123),
    .C1(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__o22a_1 _5659_ (.A1(net83),
    .A2(_1635_),
    .B1(_2466_),
    .B2(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__a22o_1 _5660_ (.A1(\ih.t.timer_max[31] ),
    .A2(_2142_),
    .B1(_2189_),
    .B2(\ih.t.timer_max[15] ),
    .X(_2471_));
 sky130_fd_sc_hd__a221o_1 _5661_ (.A1(\ih.t.timer_max[23] ),
    .A2(_2201_),
    .B1(_2311_),
    .B2(\ih.t.timer_max[7] ),
    .C1(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__and2b_1 _5662_ (.A_N(_1399_),
    .B(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__a221o_1 _5663_ (.A1(\ih.t.timer_max[23] ),
    .A2(_2147_),
    .B1(_2316_),
    .B2(\ih.t.timer_max[7] ),
    .C1(_1664_),
    .X(_2474_));
 sky130_fd_sc_hd__o21a_1 _5664_ (.A1(_1669_),
    .A2(_2473_),
    .B1(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__a22o_1 _5665_ (.A1(\mc.cl.next_data[7] ),
    .A2(_2310_),
    .B1(_2321_),
    .B2(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__a221o_1 _5666_ (.A1(\ih.gpio_interrupt_mask[7] ),
    .A2(_2323_),
    .B1(_2476_),
    .B2(_2122_),
    .C1(_2324_),
    .X(_2477_));
 sky130_fd_sc_hd__o211a_1 _5667_ (.A1(_2166_),
    .A2(_2470_),
    .B1(_2477_),
    .C1(_2134_),
    .X(_2478_));
 sky130_fd_sc_hd__a31o_1 _5668_ (.A1(net75),
    .A2(_1650_),
    .A3(_2135_),
    .B1(_2271_),
    .X(_2479_));
 sky130_fd_sc_hd__a22o_1 _5669_ (.A1(net15),
    .A2(_2342_),
    .B1(_2365_),
    .B2(net8),
    .X(_2480_));
 sky130_fd_sc_hd__and2_1 _5670_ (.A(_1651_),
    .B(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__o22a_2 _5671_ (.A1(_2478_),
    .A2(_2479_),
    .B1(_2481_),
    .B2(_1643_),
    .X(_2482_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(\cu.reg_file.reg_mem[7] ),
    .A1(_2482_),
    .S(_1658_),
    .X(_2483_));
 sky130_fd_sc_hd__clkbuf_1 _5673_ (.A(_2483_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_4 _5674_ (.A(_1643_),
    .B(_2341_),
    .Y(_2484_));
 sky130_fd_sc_hd__a22oi_1 _5675_ (.A1(\ih.t.timer_max[24] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[8] ),
    .Y(_2485_));
 sky130_fd_sc_hd__or3_2 _5676_ (.A(_1488_),
    .B(_2133_),
    .C(_1665_),
    .X(_2486_));
 sky130_fd_sc_hd__o2bb2a_1 _5677_ (.A1_N(\mc.cl.next_data[8] ),
    .A2_N(_2355_),
    .B1(_2485_),
    .B2(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__buf_2 _5678_ (.A(_1648_),
    .X(_2488_));
 sky130_fd_sc_hd__a2bb2o_1 _5679_ (.A1_N(_2487_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[8] ),
    .B2(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__a31o_1 _5680_ (.A1(net16),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2489_),
    .X(_0202_));
 sky130_fd_sc_hd__a22oi_1 _5681_ (.A1(\ih.t.timer_max[25] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[9] ),
    .Y(_2490_));
 sky130_fd_sc_hd__o2bb2a_1 _5682_ (.A1_N(\mc.cl.next_data[9] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__a2bb2o_1 _5683_ (.A1_N(_2491_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[9] ),
    .B2(_1648_),
    .X(_2492_));
 sky130_fd_sc_hd__a31o_1 _5684_ (.A1(net17),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2492_),
    .X(_0203_));
 sky130_fd_sc_hd__a22oi_1 _5685_ (.A1(\ih.t.timer_max[26] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[10] ),
    .Y(_2493_));
 sky130_fd_sc_hd__o2bb2a_1 _5686_ (.A1_N(\mc.cl.next_data[10] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__a2bb2o_1 _5687_ (.A1_N(_2494_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[10] ),
    .B2(_1648_),
    .X(_2495_));
 sky130_fd_sc_hd__a31o_1 _5688_ (.A1(net3),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2495_),
    .X(_0204_));
 sky130_fd_sc_hd__a22oi_1 _5689_ (.A1(\ih.t.timer_max[27] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[11] ),
    .Y(_2496_));
 sky130_fd_sc_hd__o2bb2a_1 _5690_ (.A1_N(\mc.cl.next_data[11] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__a2bb2o_1 _5691_ (.A1_N(_2497_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[11] ),
    .B2(_1648_),
    .X(_2498_));
 sky130_fd_sc_hd__a31o_1 _5692_ (.A1(net4),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2498_),
    .X(_0205_));
 sky130_fd_sc_hd__a22oi_1 _5693_ (.A1(\ih.t.timer_max[28] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[12] ),
    .Y(_2499_));
 sky130_fd_sc_hd__o2bb2a_1 _5694_ (.A1_N(\mc.cl.next_data[12] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__a2bb2o_1 _5695_ (.A1_N(_2500_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[12] ),
    .B2(_1648_),
    .X(_2501_));
 sky130_fd_sc_hd__a31o_1 _5696_ (.A1(net5),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2501_),
    .X(_0206_));
 sky130_fd_sc_hd__a22oi_1 _5697_ (.A1(\ih.t.timer_max[29] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[13] ),
    .Y(_2502_));
 sky130_fd_sc_hd__o2bb2a_1 _5698_ (.A1_N(\mc.cl.next_data[13] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__a2bb2o_1 _5699_ (.A1_N(_2503_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[13] ),
    .B2(_1648_),
    .X(_2504_));
 sky130_fd_sc_hd__a31o_1 _5700_ (.A1(net6),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2504_),
    .X(_0207_));
 sky130_fd_sc_hd__a22oi_1 _5701_ (.A1(\ih.t.timer_max[30] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[14] ),
    .Y(_2505_));
 sky130_fd_sc_hd__o2bb2a_1 _5702_ (.A1_N(\mc.cl.next_data[14] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__a2bb2o_1 _5703_ (.A1_N(_2506_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[14] ),
    .B2(_1648_),
    .X(_2507_));
 sky130_fd_sc_hd__a31o_1 _5704_ (.A1(net7),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2507_),
    .X(_0208_));
 sky130_fd_sc_hd__a22oi_1 _5705_ (.A1(\ih.t.timer_max[31] ),
    .A2(_2148_),
    .B1(_2317_),
    .B2(\ih.t.timer_max[15] ),
    .Y(_2508_));
 sky130_fd_sc_hd__o2bb2a_1 _5706_ (.A1_N(\mc.cl.next_data[15] ),
    .A2_N(_2355_),
    .B1(_2486_),
    .B2(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__a2bb2o_1 _5707_ (.A1_N(_2509_),
    .A2_N(_1645_),
    .B1(\cu.reg_file.reg_mem[15] ),
    .B2(_1648_),
    .X(_2510_));
 sky130_fd_sc_hd__a31o_1 _5708_ (.A1(net8),
    .A2(_1652_),
    .A3(_2484_),
    .B1(_2510_),
    .X(_0209_));
 sky130_fd_sc_hd__and3_1 _5709_ (.A(_1326_),
    .B(_1354_),
    .C(_2271_),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(net233),
    .A1(_0617_),
    .S(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _5711_ (.A(_2512_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_4 _5712_ (.A(\mc.count ),
    .X(_2513_));
 sky130_fd_sc_hd__nor2_4 _5713_ (.A(_2513_),
    .B(_1659_),
    .Y(_2514_));
 sky130_fd_sc_hd__o211a_1 _5714_ (.A1(_2711_),
    .A2(_1655_),
    .B1(_2488_),
    .C1(_2513_),
    .X(_2515_));
 sky130_fd_sc_hd__a31o_1 _5715_ (.A1(\mc.cc.enable ),
    .A2(_1668_),
    .A3(_2514_),
    .B1(_2515_),
    .X(_0211_));
 sky130_fd_sc_hd__nor2_1 _5716_ (.A(net1),
    .B(\ih.interrupt_source[3] ),
    .Y(_2516_));
 sky130_fd_sc_hd__a2111oi_1 _5717_ (.A1(net1),
    .A2(net199),
    .B1(_2873_),
    .C1(_2875_),
    .D1(_2516_),
    .Y(_0212_));
 sky130_fd_sc_hd__a22o_1 _5718_ (.A1(_2860_),
    .A2(_2873_),
    .B1(_2876_),
    .B2(net205),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _5719_ (.A(_2513_),
    .B(\mc.cl.next_data[0] ),
    .C(_2488_),
    .X(_2517_));
 sky130_fd_sc_hd__a21o_1 _5720_ (.A1(net18),
    .A2(_2514_),
    .B1(_2517_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _5721_ (.A(_2513_),
    .B(\mc.cl.next_data[1] ),
    .C(_2488_),
    .X(_2518_));
 sky130_fd_sc_hd__a21o_1 _5722_ (.A1(net19),
    .A2(_2514_),
    .B1(_2518_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _5723_ (.A(_2513_),
    .B(\mc.cl.next_data[2] ),
    .C(_2488_),
    .X(_2519_));
 sky130_fd_sc_hd__a21o_1 _5724_ (.A1(net20),
    .A2(_2514_),
    .B1(_2519_),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _5725_ (.A(_2513_),
    .B(\mc.cl.next_data[3] ),
    .C(_2488_),
    .X(_2520_));
 sky130_fd_sc_hd__a21o_1 _5726_ (.A1(net21),
    .A2(_2514_),
    .B1(_2520_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _5727_ (.A(_2513_),
    .B(\mc.cl.next_data[4] ),
    .C(_2488_),
    .X(_2521_));
 sky130_fd_sc_hd__a21o_1 _5728_ (.A1(net22),
    .A2(_2514_),
    .B1(_2521_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _5729_ (.A(_2513_),
    .B(\mc.cl.next_data[5] ),
    .C(_2488_),
    .X(_2522_));
 sky130_fd_sc_hd__a21o_1 _5730_ (.A1(net23),
    .A2(_2514_),
    .B1(_2522_),
    .X(_0219_));
 sky130_fd_sc_hd__and3_1 _5731_ (.A(_2513_),
    .B(\mc.cl.next_data[6] ),
    .C(_2488_),
    .X(_2523_));
 sky130_fd_sc_hd__a21o_1 _5732_ (.A1(net24),
    .A2(_2514_),
    .B1(_2523_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _5733_ (.A(_2513_),
    .B(\mc.cl.next_data[7] ),
    .C(_2488_),
    .X(_2524_));
 sky130_fd_sc_hd__a21o_1 _5734_ (.A1(net25),
    .A2(_2514_),
    .B1(_2524_),
    .X(_0221_));
 sky130_fd_sc_hd__or2_2 _5735_ (.A(\mc.cc.count[0] ),
    .B(_2711_),
    .X(_2525_));
 sky130_fd_sc_hd__nor2_1 _5736_ (.A(_1654_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__a22o_1 _5737_ (.A1(net214),
    .A2(_2711_),
    .B1(_2526_),
    .B2(\mc.cc.enable_edge_detector.prev_data ),
    .X(_0222_));
 sky130_fd_sc_hd__or2_1 _5738_ (.A(\mc.cc.enable_edge_detector.prev_data ),
    .B(_2711_),
    .X(_2527_));
 sky130_fd_sc_hd__o21ai_1 _5739_ (.A1(\mc.cc.count[1] ),
    .A2(_2525_),
    .B1(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__a21o_1 _5740_ (.A1(net227),
    .A2(_2525_),
    .B1(_2528_),
    .X(_0223_));
 sky130_fd_sc_hd__nor3_1 _5741_ (.A(\mc.cc.count[2] ),
    .B(\mc.cc.count[1] ),
    .C(_2525_),
    .Y(_2529_));
 sky130_fd_sc_hd__o211a_1 _5742_ (.A1(\mc.cc.count[1] ),
    .A2(_2525_),
    .B1(_2527_),
    .C1(\mc.cc.count[2] ),
    .X(_2530_));
 sky130_fd_sc_hd__a31o_1 _5743_ (.A1(net210),
    .A2(\mc.cc.enable_edge_detector.prev_data ),
    .A3(_2529_),
    .B1(_2530_),
    .X(_0224_));
 sky130_fd_sc_hd__and3b_1 _5744_ (.A_N(_2529_),
    .B(\mc.cc.count[3] ),
    .C(_2527_),
    .X(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _5745_ (.A(_2531_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _5746_ (.A(\cu.reg_file.reg_sp[1] ),
    .Y(_2532_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(_2532_),
    .A1(_1048_),
    .S(_2120_),
    .X(_2533_));
 sky130_fd_sc_hd__or4b_2 _5748_ (.A(_1007_),
    .B(_0980_),
    .C(_0989_),
    .D_N(_0994_),
    .X(_2534_));
 sky130_fd_sc_hd__or2_1 _5749_ (.A(_0296_),
    .B(_0471_),
    .X(_2535_));
 sky130_fd_sc_hd__clkbuf_2 _5750_ (.A(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__buf_2 _5751_ (.A(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__buf_4 _5752_ (.A(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__o21ai_2 _5753_ (.A1(_0986_),
    .A2(_2534_),
    .B1(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__o31a_4 _5754_ (.A1(_0739_),
    .A2(_2120_),
    .A3(_2539_),
    .B1(_2952_),
    .X(_2540_));
 sky130_fd_sc_hd__buf_4 _5755_ (.A(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(\cu.reg_file.reg_sp[1] ),
    .A1(_2533_),
    .S(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__clkbuf_1 _5757_ (.A(_2542_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(\cu.reg_file.reg_sp[2] ),
    .B(_2536_),
    .Y(_2543_));
 sky130_fd_sc_hd__or2_1 _5759_ (.A(\cu.reg_file.reg_sp[2] ),
    .B(_2536_),
    .X(_2544_));
 sky130_fd_sc_hd__and2_1 _5760_ (.A(_2543_),
    .B(_2544_),
    .X(_2545_));
 sky130_fd_sc_hd__xnor2_1 _5761_ (.A(_2532_),
    .B(_2545_),
    .Y(_2546_));
 sky130_fd_sc_hd__buf_4 _5762_ (.A(_2119_),
    .X(_2547_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(_1070_),
    .A1(_2546_),
    .S(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(\cu.reg_file.reg_sp[2] ),
    .A1(_2548_),
    .S(_2541_),
    .X(_2549_));
 sky130_fd_sc_hd__clkbuf_1 _5765_ (.A(_2549_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _5766_ (.A(\cu.reg_file.reg_sp[3] ),
    .B(_2536_),
    .Y(_2550_));
 sky130_fd_sc_hd__and2_1 _5767_ (.A(\cu.reg_file.reg_sp[3] ),
    .B(_2536_),
    .X(_2551_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(_2550_),
    .B(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__a21bo_1 _5769_ (.A1(\cu.reg_file.reg_sp[1] ),
    .A2(_2545_),
    .B1_N(_2543_),
    .X(_2553_));
 sky130_fd_sc_hd__xor2_1 _5770_ (.A(_2552_),
    .B(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(_1087_),
    .A1(_2554_),
    .S(_2547_),
    .X(_2555_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(\cu.reg_file.reg_sp[3] ),
    .A1(_2555_),
    .S(_2541_),
    .X(_2556_));
 sky130_fd_sc_hd__clkbuf_1 _5773_ (.A(_2556_),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _5774_ (.A(\cu.reg_file.reg_sp[4] ),
    .B(_2536_),
    .Y(_2557_));
 sky130_fd_sc_hd__and2_1 _5775_ (.A(\cu.reg_file.reg_sp[4] ),
    .B(_2536_),
    .X(_2558_));
 sky130_fd_sc_hd__nor2_1 _5776_ (.A(_2557_),
    .B(_2558_),
    .Y(_2559_));
 sky130_fd_sc_hd__a21o_1 _5777_ (.A1(_2552_),
    .A2(_2553_),
    .B1(_2551_),
    .X(_2560_));
 sky130_fd_sc_hd__xor2_1 _5778_ (.A(_2559_),
    .B(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(_1159_),
    .A1(_2561_),
    .S(_2547_),
    .X(_2562_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(\cu.reg_file.reg_sp[4] ),
    .A1(_2562_),
    .S(_2541_),
    .X(_2563_));
 sky130_fd_sc_hd__clkbuf_1 _5781_ (.A(_2563_),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _5782_ (.A(\cu.reg_file.reg_sp[5] ),
    .B(_2537_),
    .X(_2564_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(\cu.reg_file.reg_sp[5] ),
    .B(_2537_),
    .Y(_2565_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(_2564_),
    .B(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__a311o_1 _5785_ (.A1(_2552_),
    .A2(_2553_),
    .A3(_2559_),
    .B1(_2558_),
    .C1(_2551_),
    .X(_2567_));
 sky130_fd_sc_hd__xnor2_1 _5786_ (.A(_2566_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(_1143_),
    .A1(_2568_),
    .S(_2547_),
    .X(_2569_));
 sky130_fd_sc_hd__mux2_1 _5788_ (.A0(\cu.reg_file.reg_sp[5] ),
    .A1(_2569_),
    .S(_2541_),
    .X(_2570_));
 sky130_fd_sc_hd__clkbuf_1 _5789_ (.A(_2570_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _5790_ (.A(\cu.reg_file.reg_sp[6] ),
    .B(_2537_),
    .X(_2571_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(\cu.reg_file.reg_sp[6] ),
    .B(_2537_),
    .Y(_2572_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(_2571_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__a21bo_1 _5793_ (.A1(_2564_),
    .A2(_2567_),
    .B1_N(_2565_),
    .X(_2574_));
 sky130_fd_sc_hd__xnor2_1 _5794_ (.A(_2573_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(_1125_),
    .A1(_2575_),
    .S(_2547_),
    .X(_2576_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(\cu.reg_file.reg_sp[6] ),
    .A1(_2576_),
    .S(_2541_),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _5797_ (.A(_2577_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _5798_ (.A(\cu.reg_file.reg_sp[7] ),
    .B(_2537_),
    .X(_2578_));
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(\cu.reg_file.reg_sp[7] ),
    .B(_2537_),
    .Y(_2579_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_2578_),
    .B(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__a21bo_1 _5801_ (.A1(_2571_),
    .A2(_2574_),
    .B1_N(_2572_),
    .X(_2581_));
 sky130_fd_sc_hd__xnor2_1 _5802_ (.A(_2580_),
    .B(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__mux2_1 _5803_ (.A0(_1108_),
    .A1(_2582_),
    .S(_2547_),
    .X(_2583_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(\cu.reg_file.reg_sp[7] ),
    .A1(_2583_),
    .S(_2541_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _5805_ (.A(_2584_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _5806_ (.A(\cu.reg_file.reg_sp[8] ),
    .B(_2537_),
    .X(_2585_));
 sky130_fd_sc_hd__nand2_1 _5807_ (.A(\cu.reg_file.reg_sp[8] ),
    .B(_2537_),
    .Y(_2586_));
 sky130_fd_sc_hd__nand2_1 _5808_ (.A(_2585_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__a21bo_1 _5809_ (.A1(_2578_),
    .A2(_2581_),
    .B1_N(_2579_),
    .X(_2588_));
 sky130_fd_sc_hd__xnor2_1 _5810_ (.A(_2587_),
    .B(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(_1624_),
    .A1(_2589_),
    .S(_2547_),
    .X(_2590_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(\cu.reg_file.reg_sp[8] ),
    .A1(_2590_),
    .S(_2541_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _5813_ (.A(_2591_),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _5814_ (.A(\cu.reg_file.reg_sp[9] ),
    .B(_2537_),
    .X(_2592_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(\cu.reg_file.reg_sp[9] ),
    .B(_2538_),
    .Y(_2593_));
 sky130_fd_sc_hd__nand2_1 _5816_ (.A(_2592_),
    .B(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__a21bo_1 _5817_ (.A1(_2585_),
    .A2(_2588_),
    .B1_N(_2586_),
    .X(_2595_));
 sky130_fd_sc_hd__xnor2_1 _5818_ (.A(_2594_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(_1625_),
    .A1(_2596_),
    .S(_2547_),
    .X(_2597_));
 sky130_fd_sc_hd__mux2_1 _5820_ (.A0(\cu.reg_file.reg_sp[9] ),
    .A1(_2597_),
    .S(_2541_),
    .X(_2598_));
 sky130_fd_sc_hd__clkbuf_1 _5821_ (.A(_2598_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _5822_ (.A(\cu.reg_file.reg_sp[10] ),
    .B(_2538_),
    .X(_2599_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(\cu.reg_file.reg_sp[10] ),
    .B(_2538_),
    .Y(_2600_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_2599_),
    .B(_2600_),
    .Y(_2601_));
 sky130_fd_sc_hd__a21bo_1 _5825_ (.A1(_2592_),
    .A2(_2595_),
    .B1_N(_2593_),
    .X(_2602_));
 sky130_fd_sc_hd__xnor2_1 _5826_ (.A(_2601_),
    .B(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(_1225_),
    .A1(_2603_),
    .S(_2547_),
    .X(_2604_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(\cu.reg_file.reg_sp[10] ),
    .A1(_2604_),
    .S(_2541_),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _5829_ (.A(_2605_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _5830_ (.A(\cu.reg_file.reg_sp[11] ),
    .B(_2538_),
    .X(_2606_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(\cu.reg_file.reg_sp[11] ),
    .B(_2538_),
    .Y(_2607_));
 sky130_fd_sc_hd__nand2_1 _5832_ (.A(_2606_),
    .B(_2607_),
    .Y(_2608_));
 sky130_fd_sc_hd__a21bo_1 _5833_ (.A1(_2599_),
    .A2(_2602_),
    .B1_N(_2600_),
    .X(_2609_));
 sky130_fd_sc_hd__xnor2_1 _5834_ (.A(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(_1221_),
    .A1(_2610_),
    .S(_2547_),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(\cu.reg_file.reg_sp[11] ),
    .A1(_2611_),
    .S(_2540_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _5837_ (.A(_2612_),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _5838_ (.A(\cu.reg_file.reg_sp[12] ),
    .B(_2538_),
    .X(_2613_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(\cu.reg_file.reg_sp[12] ),
    .B(_2538_),
    .Y(_2614_));
 sky130_fd_sc_hd__nand2_1 _5840_ (.A(_2613_),
    .B(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__a21bo_1 _5841_ (.A1(_2606_),
    .A2(_2609_),
    .B1_N(_2607_),
    .X(_2616_));
 sky130_fd_sc_hd__xnor2_1 _5842_ (.A(_2615_),
    .B(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(_1212_),
    .A1(_2617_),
    .S(_2119_),
    .X(_2618_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(\cu.reg_file.reg_sp[12] ),
    .A1(_2618_),
    .S(_2540_),
    .X(_2619_));
 sky130_fd_sc_hd__clkbuf_1 _5845_ (.A(_2619_),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _5846_ (.A(\cu.reg_file.reg_sp[13] ),
    .B(_2538_),
    .X(_2620_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(\cu.reg_file.reg_sp[13] ),
    .B(_2538_),
    .Y(_2621_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_2620_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__a21bo_1 _5849_ (.A1(_2613_),
    .A2(_2616_),
    .B1_N(_2614_),
    .X(_2623_));
 sky130_fd_sc_hd__xnor2_1 _5850_ (.A(_2622_),
    .B(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(_1208_),
    .A1(_2624_),
    .S(_2119_),
    .X(_2625_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(\cu.reg_file.reg_sp[13] ),
    .A1(_2625_),
    .S(_2540_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_1 _5853_ (.A(_2626_),
    .X(_0238_));
 sky130_fd_sc_hd__xnor2_1 _5854_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1286_),
    .Y(_2627_));
 sky130_fd_sc_hd__a21boi_2 _5855_ (.A1(_2620_),
    .A2(_2623_),
    .B1_N(_2621_),
    .Y(_2628_));
 sky130_fd_sc_hd__xnor2_1 _5856_ (.A(_2627_),
    .B(_2628_),
    .Y(_2629_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(_1626_),
    .A1(_2629_),
    .S(_2119_),
    .X(_2630_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(\cu.reg_file.reg_sp[14] ),
    .A1(_2630_),
    .S(_2540_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _5859_ (.A(_2631_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _5860_ (.A(\cu.reg_file.reg_sp[14] ),
    .B(_1286_),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(_1591_),
    .A1(_2632_),
    .S(_2628_),
    .X(_2633_));
 sky130_fd_sc_hd__xnor2_1 _5862_ (.A(\cu.reg_file.reg_sp[15] ),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(_1262_),
    .A1(_2634_),
    .S(_2119_),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(\cu.reg_file.reg_sp[15] ),
    .A1(_2635_),
    .S(_2540_),
    .X(_2636_));
 sky130_fd_sc_hd__clkbuf_1 _5865_ (.A(_2636_),
    .X(_0240_));
 sky130_fd_sc_hd__and3_2 _5866_ (.A(_1357_),
    .B(_1633_),
    .C(_2317_),
    .X(_2637_));
 sky130_fd_sc_hd__o21ai_4 _5867_ (.A1(_1671_),
    .A2(_2191_),
    .B1(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(_2141_),
    .A1(\ih.t.timer_max[8] ),
    .S(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _5869_ (.A(_2639_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(_2152_),
    .A1(\ih.t.timer_max[9] ),
    .S(_2638_),
    .X(_2640_));
 sky130_fd_sc_hd__clkbuf_1 _5871_ (.A(_2640_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(_2154_),
    .A1(\ih.t.timer_max[10] ),
    .S(_2638_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _5873_ (.A(_2641_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(_2156_),
    .A1(\ih.t.timer_max[11] ),
    .S(_2638_),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_1 _5875_ (.A(_2642_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(_2158_),
    .A1(\ih.t.timer_max[12] ),
    .S(_2638_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5877_ (.A(_2643_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_2160_),
    .A1(\ih.t.timer_max[13] ),
    .S(_2638_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_1 _5879_ (.A(_2644_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(_2162_),
    .A1(\ih.t.timer_max[14] ),
    .S(_2638_),
    .X(_2645_));
 sky130_fd_sc_hd__clkbuf_1 _5881_ (.A(_2645_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(_2164_),
    .A1(\ih.t.timer_max[15] ),
    .S(_2638_),
    .X(_2646_));
 sky130_fd_sc_hd__clkbuf_1 _5883_ (.A(_2646_),
    .X(_0248_));
 sky130_fd_sc_hd__o21ai_4 _5884_ (.A1(_1671_),
    .A2(_2177_),
    .B1(_2637_),
    .Y(_2647_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(_2025_),
    .A1(\ih.t.timer_max[0] ),
    .S(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _5886_ (.A(_2648_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5887_ (.A0(_1049_),
    .A1(\ih.t.timer_max[1] ),
    .S(_2647_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _5888_ (.A(_2649_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(_1071_),
    .A1(\ih.t.timer_max[2] ),
    .S(_2647_),
    .X(_2650_));
 sky130_fd_sc_hd__clkbuf_1 _5890_ (.A(_2650_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5891_ (.A0(_1186_),
    .A1(\ih.t.timer_max[3] ),
    .S(_2647_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _5892_ (.A(_2651_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5893_ (.A0(_1188_),
    .A1(\ih.t.timer_max[4] ),
    .S(_2647_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5894_ (.A(_2652_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5895_ (.A0(_1190_),
    .A1(\ih.t.timer_max[5] ),
    .S(_2647_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5896_ (.A(_2653_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(_1192_),
    .A1(\ih.t.timer_max[6] ),
    .S(_2647_),
    .X(_2654_));
 sky130_fd_sc_hd__clkbuf_1 _5898_ (.A(_2654_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5899_ (.A0(_1259_),
    .A1(\ih.t.timer_max[7] ),
    .S(_2647_),
    .X(_2655_));
 sky130_fd_sc_hd__clkbuf_1 _5900_ (.A(_2655_),
    .X(_0256_));
 sky130_fd_sc_hd__o21a_4 _5901_ (.A1(_1671_),
    .A2(_2202_),
    .B1(_2149_),
    .X(_2656_));
 sky130_fd_sc_hd__mux2_1 _5902_ (.A0(\ih.t.timer_max[16] ),
    .A1(_0617_),
    .S(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _5903_ (.A(_2657_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(\ih.t.timer_max[17] ),
    .A1(_1049_),
    .S(_2656_),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _5905_ (.A(_2658_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(\ih.t.timer_max[18] ),
    .A1(_1071_),
    .S(_2656_),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _5907_ (.A(_2659_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(\ih.t.timer_max[19] ),
    .A1(_1186_),
    .S(_2656_),
    .X(_2660_));
 sky130_fd_sc_hd__clkbuf_1 _5909_ (.A(_2660_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(\ih.t.timer_max[20] ),
    .A1(_1188_),
    .S(_2656_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _5911_ (.A(_2661_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(\ih.t.timer_max[21] ),
    .A1(_1190_),
    .S(_2656_),
    .X(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _5913_ (.A(_2662_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5914_ (.A0(\ih.t.timer_max[22] ),
    .A1(_1192_),
    .S(_2656_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_1 _5915_ (.A(_2663_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(\ih.t.timer_max[23] ),
    .A1(_1259_),
    .S(_2656_),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_1 _5917_ (.A(_2664_),
    .X(_0264_));
 sky130_fd_sc_hd__inv_2 _5918_ (.A(\cu.ir.idx[0] ),
    .Y(_2665_));
 sky130_fd_sc_hd__o21a_1 _5919_ (.A1(_2665_),
    .A2(_1646_),
    .B1(_1483_),
    .X(_2666_));
 sky130_fd_sc_hd__a21o_1 _5920_ (.A1(_2951_),
    .A2(_1481_),
    .B1(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__a22o_1 _5921_ (.A1(_1659_),
    .A2(_2666_),
    .B1(_2667_),
    .B2(net222),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_4 _5922_ (.A(_2665_),
    .B(\cu.ir.idx[1] ),
    .Y(_2668_));
 sky130_fd_sc_hd__a32o_1 _5923_ (.A1(_1483_),
    .A2(_1659_),
    .A3(_2668_),
    .B1(_2667_),
    .B2(net236),
    .X(_0266_));
 sky130_fd_sc_hd__o21ai_1 _5924_ (.A1(_1783_),
    .A2(_2534_),
    .B1(net202),
    .Y(_2669_));
 sky130_fd_sc_hd__o21ai_1 _5925_ (.A1(net203),
    .A2(_2669_),
    .B1(_1784_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_4 _5926_ (.A(\cu.ir.idx[0] ),
    .B(\cu.ir.idx[1] ),
    .Y(_2670_));
 sky130_fd_sc_hd__mux2_1 _5927_ (.A0(_2934_),
    .A1(_2347_),
    .S(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_1 _5928_ (.A(_2671_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5929_ (.A0(_2903_),
    .A1(_2368_),
    .S(_2670_),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_1 _5930_ (.A(_2672_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(_2902_),
    .A1(_2387_),
    .S(_2670_),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_1 _5932_ (.A(_2673_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5933_ (.A0(_2896_),
    .A1(_2406_),
    .S(_2670_),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _5934_ (.A(_2674_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(_0359_),
    .A1(_2425_),
    .S(_2670_),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_1 _5936_ (.A(_2675_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(_2922_),
    .A1(_2444_),
    .S(_2670_),
    .X(_2676_));
 sky130_fd_sc_hd__clkbuf_1 _5938_ (.A(_2676_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(_2878_),
    .A1(_2463_),
    .S(_2670_),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_1 _5940_ (.A(_2677_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(_2879_),
    .A1(_2482_),
    .S(_2670_),
    .X(_2678_));
 sky130_fd_sc_hd__clkbuf_1 _5942_ (.A(_2678_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(_0344_),
    .A1(_2347_),
    .S(_2668_),
    .X(_2679_));
 sky130_fd_sc_hd__clkbuf_1 _5944_ (.A(_2679_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(_0341_),
    .A1(_2368_),
    .S(_2668_),
    .X(_2680_));
 sky130_fd_sc_hd__clkbuf_1 _5946_ (.A(_2680_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5947_ (.A0(_0342_),
    .A1(_2387_),
    .S(_2668_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_1 _5948_ (.A(_2681_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5949_ (.A0(\cu.id.cb_opcode_y[0] ),
    .A1(_2406_),
    .S(_2668_),
    .X(_2682_));
 sky130_fd_sc_hd__clkbuf_1 _5950_ (.A(_2682_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5951_ (.A0(_0374_),
    .A1(_2425_),
    .S(_2668_),
    .X(_2683_));
 sky130_fd_sc_hd__clkbuf_1 _5952_ (.A(_2683_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5953_ (.A0(_0373_),
    .A1(_2444_),
    .S(_2668_),
    .X(_2684_));
 sky130_fd_sc_hd__clkbuf_1 _5954_ (.A(_2684_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5955_ (.A0(_0387_),
    .A1(_2463_),
    .S(_2668_),
    .X(_2685_));
 sky130_fd_sc_hd__clkbuf_1 _5956_ (.A(_2685_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5957_ (.A0(_1232_),
    .A1(_2482_),
    .S(_2668_),
    .X(_2686_));
 sky130_fd_sc_hd__clkbuf_1 _5958_ (.A(_2686_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _5959_ (.A(_2665_),
    .B(\cu.ir.idx[1] ),
    .X(_2687_));
 sky130_fd_sc_hd__buf_2 _5960_ (.A(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__mux2_1 _5961_ (.A0(\cu.id.imm_i[8] ),
    .A1(_2347_),
    .S(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__clkbuf_1 _5962_ (.A(_2689_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _5963_ (.A0(\cu.id.imm_i[9] ),
    .A1(_2368_),
    .S(_2688_),
    .X(_2690_));
 sky130_fd_sc_hd__clkbuf_1 _5964_ (.A(_2690_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _5965_ (.A0(\cu.id.imm_i[10] ),
    .A1(_2387_),
    .S(_2688_),
    .X(_2691_));
 sky130_fd_sc_hd__clkbuf_1 _5966_ (.A(_2691_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5967_ (.A0(\cu.id.imm_i[11] ),
    .A1(_2406_),
    .S(_2688_),
    .X(_2692_));
 sky130_fd_sc_hd__clkbuf_1 _5968_ (.A(_2692_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(\cu.id.imm_i[12] ),
    .A1(_2425_),
    .S(_2688_),
    .X(_2693_));
 sky130_fd_sc_hd__clkbuf_1 _5970_ (.A(_2693_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(\cu.id.imm_i[13] ),
    .A1(_2444_),
    .S(_2688_),
    .X(_2694_));
 sky130_fd_sc_hd__clkbuf_1 _5972_ (.A(_2694_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5973_ (.A0(\cu.id.imm_i[14] ),
    .A1(_2463_),
    .S(_2688_),
    .X(_2695_));
 sky130_fd_sc_hd__clkbuf_1 _5974_ (.A(_2695_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(\cu.id.imm_i[15] ),
    .A1(_2482_),
    .S(_2688_),
    .X(_2696_));
 sky130_fd_sc_hd__clkbuf_1 _5976_ (.A(_2696_),
    .X(_0291_));
 sky130_fd_sc_hd__dfrtp_4 _5977_ (.CLK(clknet_leaf_39_clk),
    .D(_0007_),
    .RESET_B(net151),
    .Q(\alu.Cin ));
 sky130_fd_sc_hd__dfrtp_1 _5978_ (.CLK(clknet_leaf_38_clk),
    .D(_0008_),
    .RESET_B(net151),
    .Q(\cu.alu_f[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5979_ (.CLK(clknet_leaf_38_clk),
    .D(_0009_),
    .RESET_B(net151),
    .Q(\cu.alu_f[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5980_ (.CLK(clknet_leaf_38_clk),
    .D(_0010_),
    .RESET_B(net152),
    .Q(\cu.alu_f[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5981_ (.CLK(clknet_leaf_38_clk),
    .D(_0011_),
    .RESET_B(net152),
    .Q(\cu.alu_f[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5982_ (.CLK(clknet_leaf_38_clk),
    .D(_0012_),
    .RESET_B(net152),
    .Q(\cu.alu_f[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5983_ (.CLK(clknet_leaf_38_clk),
    .D(_0013_),
    .RESET_B(net152),
    .Q(\cu.alu_f[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5984_ (.CLK(clknet_leaf_38_clk),
    .D(_0014_),
    .RESET_B(net152),
    .Q(\cu.alu_f[7] ));
 sky130_fd_sc_hd__dfrtp_2 _5985_ (.CLK(clknet_leaf_33_clk),
    .D(_0016_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[0] ));
 sky130_fd_sc_hd__dfrtp_4 _5986_ (.CLK(clknet_leaf_33_clk),
    .D(_0017_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5987_ (.CLK(clknet_leaf_33_clk),
    .D(_0018_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _5988_ (.CLK(clknet_leaf_34_clk),
    .D(_0019_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5989_ (.CLK(clknet_leaf_34_clk),
    .D(_0020_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _5990_ (.CLK(clknet_leaf_33_clk),
    .D(_0021_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _5991_ (.CLK(clknet_leaf_28_clk),
    .D(_0022_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _5992_ (.CLK(clknet_leaf_28_clk),
    .D(_0023_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _5993_ (.CLK(clknet_leaf_27_clk),
    .D(_0024_),
    .RESET_B(net184),
    .Q(\cu.pc.pc_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _5994_ (.CLK(clknet_leaf_27_clk),
    .D(_0025_),
    .RESET_B(net184),
    .Q(\cu.pc.pc_o[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5995_ (.CLK(clknet_leaf_29_clk),
    .D(_0026_),
    .RESET_B(net184),
    .Q(\cu.pc.pc_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _5996_ (.CLK(clknet_leaf_27_clk),
    .D(_0027_),
    .RESET_B(net184),
    .Q(\cu.pc.pc_o[11] ));
 sky130_fd_sc_hd__dfstp_2 _5997_ (.CLK(clknet_leaf_29_clk),
    .D(_0028_),
    .SET_B(net186),
    .Q(\cu.pc.pc_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _5998_ (.CLK(clknet_leaf_28_clk),
    .D(_0029_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _5999_ (.CLK(clknet_leaf_28_clk),
    .D(_0030_),
    .RESET_B(net186),
    .Q(\cu.pc.pc_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6000_ (.CLK(clknet_leaf_33_clk),
    .D(_0031_),
    .RESET_B(net160),
    .Q(\cu.pc.pc_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6001_ (.CLK(clknet_leaf_30_clk),
    .D(_0032_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_a[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6002_ (.CLK(clknet_leaf_3_clk),
    .D(_0033_),
    .RESET_B(net168),
    .Q(\cu.reg_file.reg_a[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6003_ (.CLK(clknet_leaf_30_clk),
    .D(_0034_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_a[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6004_ (.CLK(clknet_leaf_30_clk),
    .D(_0035_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_a[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6005_ (.CLK(clknet_leaf_32_clk),
    .D(_0036_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_a[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6006_ (.CLK(clknet_leaf_32_clk),
    .D(_0037_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_a[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6007_ (.CLK(clknet_leaf_30_clk),
    .D(_0038_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_a[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6008_ (.CLK(clknet_leaf_37_clk),
    .D(_0039_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_a[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6009_ (.CLK(clknet_leaf_30_clk),
    .D(_0040_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6010_ (.CLK(clknet_leaf_2_clk),
    .D(_0041_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_b[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6011_ (.CLK(clknet_leaf_29_clk),
    .D(_0042_),
    .RESET_B(net184),
    .Q(\cu.reg_file.reg_b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6012_ (.CLK(clknet_leaf_30_clk),
    .D(_0043_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_b[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6013_ (.CLK(clknet_leaf_29_clk),
    .D(_0044_),
    .RESET_B(net184),
    .Q(\cu.reg_file.reg_b[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6014_ (.CLK(clknet_leaf_29_clk),
    .D(_0045_),
    .RESET_B(net186),
    .Q(\cu.reg_file.reg_b[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6015_ (.CLK(clknet_leaf_29_clk),
    .D(_0046_),
    .RESET_B(net186),
    .Q(\cu.reg_file.reg_b[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6016_ (.CLK(clknet_leaf_29_clk),
    .D(_0047_),
    .RESET_B(net186),
    .Q(\cu.reg_file.reg_b[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6017_ (.CLK(clknet_leaf_16_clk),
    .D(_0048_),
    .RESET_B(net168),
    .Q(\cu.reg_file.reg_c[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6018_ (.CLK(clknet_leaf_2_clk),
    .D(_0049_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_c[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6019_ (.CLK(clknet_leaf_17_clk),
    .D(_0050_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_c[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6020_ (.CLK(clknet_leaf_17_clk),
    .D(_0051_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_c[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6021_ (.CLK(clknet_leaf_17_clk),
    .D(_0052_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_c[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6022_ (.CLK(clknet_leaf_31_clk),
    .D(_0053_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_c[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6023_ (.CLK(clknet_leaf_30_clk),
    .D(_0054_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_c[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6024_ (.CLK(clknet_leaf_16_clk),
    .D(_0055_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_c[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6025_ (.CLK(clknet_leaf_32_clk),
    .D(_0056_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_d[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6026_ (.CLK(clknet_leaf_3_clk),
    .D(_0057_),
    .RESET_B(net167),
    .Q(\cu.reg_file.reg_d[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6027_ (.CLK(clknet_leaf_30_clk),
    .D(_0058_),
    .RESET_B(net186),
    .Q(\cu.reg_file.reg_d[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6028_ (.CLK(clknet_leaf_30_clk),
    .D(_0059_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_d[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6029_ (.CLK(clknet_leaf_35_clk),
    .D(_0060_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_d[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6030_ (.CLK(clknet_leaf_35_clk),
    .D(_0061_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_d[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6031_ (.CLK(clknet_leaf_29_clk),
    .D(_0062_),
    .RESET_B(net186),
    .Q(\cu.reg_file.reg_d[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6032_ (.CLK(clknet_leaf_32_clk),
    .D(_0063_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_d[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6033_ (.CLK(clknet_leaf_2_clk),
    .D(_0064_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_e[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6034_ (.CLK(clknet_leaf_2_clk),
    .D(_0065_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_e[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6035_ (.CLK(clknet_leaf_3_clk),
    .D(_0066_),
    .RESET_B(net167),
    .Q(\cu.reg_file.reg_e[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6036_ (.CLK(clknet_leaf_3_clk),
    .D(_0067_),
    .RESET_B(net168),
    .Q(\cu.reg_file.reg_e[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6037_ (.CLK(clknet_leaf_3_clk),
    .D(_0068_),
    .RESET_B(net167),
    .Q(\cu.reg_file.reg_e[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6038_ (.CLK(clknet_leaf_3_clk),
    .D(_0069_),
    .RESET_B(net168),
    .Q(\cu.reg_file.reg_e[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6039_ (.CLK(clknet_leaf_17_clk),
    .D(_0070_),
    .RESET_B(net168),
    .Q(\cu.reg_file.reg_e[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6040_ (.CLK(clknet_leaf_17_clk),
    .D(_0071_),
    .RESET_B(net169),
    .Q(\cu.reg_file.reg_e[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6041_ (.CLK(clknet_leaf_35_clk),
    .D(_0072_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_h[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6042_ (.CLK(clknet_leaf_35_clk),
    .D(_0073_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_h[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6043_ (.CLK(clknet_leaf_35_clk),
    .D(_0074_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_h[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6044_ (.CLK(clknet_leaf_36_clk),
    .D(_0075_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_h[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6045_ (.CLK(clknet_leaf_34_clk),
    .D(_0076_),
    .RESET_B(net159),
    .Q(\cu.reg_file.reg_h[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6046_ (.CLK(clknet_leaf_36_clk),
    .D(_0077_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_h[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6047_ (.CLK(clknet_leaf_36_clk),
    .D(_0078_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_h[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6048_ (.CLK(clknet_leaf_36_clk),
    .D(_0079_),
    .RESET_B(net161),
    .Q(\cu.reg_file.reg_h[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6049_ (.CLK(clknet_leaf_16_clk),
    .D(_0080_),
    .RESET_B(net169),
    .Q(\cu.reg_file.reg_l[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6050_ (.CLK(clknet_leaf_3_clk),
    .D(_0081_),
    .RESET_B(net167),
    .Q(\cu.reg_file.reg_l[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6051_ (.CLK(clknet_leaf_17_clk),
    .D(_0082_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_l[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6052_ (.CLK(clknet_leaf_16_clk),
    .D(_0083_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_l[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6053_ (.CLK(clknet_leaf_17_clk),
    .D(_0084_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_l[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6054_ (.CLK(clknet_leaf_31_clk),
    .D(_0085_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_l[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6055_ (.CLK(clknet_leaf_30_clk),
    .D(_0086_),
    .RESET_B(net181),
    .Q(\cu.reg_file.reg_l[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6056_ (.CLK(clknet_leaf_16_clk),
    .D(_0087_),
    .RESET_B(net169),
    .Q(\cu.reg_file.reg_l[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6057_ (.CLK(clknet_leaf_20_clk),
    .D(_0088_),
    .RESET_B(net188),
    .Q(\mc.cl.next_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6058_ (.CLK(clknet_leaf_20_clk),
    .D(_0089_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6059_ (.CLK(clknet_leaf_20_clk),
    .D(_0090_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6060_ (.CLK(clknet_leaf_21_clk),
    .D(_0091_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6061_ (.CLK(clknet_leaf_20_clk),
    .D(_0092_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6062_ (.CLK(clknet_leaf_23_clk),
    .D(_0093_),
    .RESET_B(net190),
    .Q(\mc.cl.next_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6063_ (.CLK(clknet_leaf_20_clk),
    .D(_0094_),
    .RESET_B(net189),
    .Q(\mc.cl.next_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6064_ (.CLK(clknet_leaf_20_clk),
    .D(_0095_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6065_ (.CLK(clknet_leaf_24_clk),
    .D(\mc.cc.enable ),
    .RESET_B(net192),
    .Q(\mc.cc.enable_edge_detector.prev_data ));
 sky130_fd_sc_hd__dfrtp_2 _6066_ (.CLK(clknet_leaf_2_clk),
    .D(_0096_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_sp[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6067_ (.CLK(clknet_leaf_23_clk),
    .D(\mc.rw.next_state[0] ),
    .RESET_B(net188),
    .Q(\mc.rw.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6068_ (.CLK(clknet_leaf_23_clk),
    .D(\mc.rw.next_state[1] ),
    .RESET_B(net192),
    .Q(\mc.rw.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6069_ (.CLK(clknet_leaf_23_clk),
    .D(\mc.rw.next_state[2] ),
    .RESET_B(net188),
    .Q(\mc.rw.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6070_ (.CLK(clknet_leaf_24_clk),
    .D(\mc.rw.cmp_check ),
    .RESET_B(net192),
    .Q(\mc.cl.cmp_o ));
 sky130_fd_sc_hd__dfrtp_1 _6071_ (.CLK(clknet_leaf_15_clk),
    .D(_0097_),
    .RESET_B(net175),
    .Q(\ih.gpio_interrupt_mask[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6072_ (.CLK(clknet_leaf_8_clk),
    .D(_0098_),
    .RESET_B(net171),
    .Q(\ih.gpio_interrupt_mask[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6073_ (.CLK(clknet_leaf_7_clk),
    .D(_0099_),
    .RESET_B(net166),
    .Q(\ih.gpio_interrupt_mask[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6074_ (.CLK(clknet_leaf_7_clk),
    .D(_0100_),
    .RESET_B(net166),
    .Q(\ih.gpio_interrupt_mask[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6075_ (.CLK(clknet_leaf_7_clk),
    .D(_0101_),
    .RESET_B(net166),
    .Q(\ih.gpio_interrupt_mask[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6076_ (.CLK(clknet_leaf_11_clk),
    .D(_0102_),
    .RESET_B(net171),
    .Q(\ih.gpio_interrupt_mask[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6077_ (.CLK(clknet_leaf_11_clk),
    .D(_0103_),
    .RESET_B(net175),
    .Q(\ih.gpio_interrupt_mask[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6078_ (.CLK(clknet_leaf_11_clk),
    .D(_0104_),
    .RESET_B(net175),
    .Q(\ih.gpio_interrupt_mask[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6079_ (.CLK(clknet_leaf_15_clk),
    .D(_0105_),
    .RESET_B(net175),
    .Q(\ih.t.enable ));
 sky130_fd_sc_hd__dfrtp_2 _6080_ (.CLK(clknet_leaf_21_clk),
    .D(_0106_),
    .RESET_B(net189),
    .Q(\ih.t.timer_max[24] ));
 sky130_fd_sc_hd__dfrtp_4 _6081_ (.CLK(clknet_leaf_14_clk),
    .D(_0107_),
    .RESET_B(net189),
    .Q(\ih.t.timer_max[25] ));
 sky130_fd_sc_hd__dfrtp_2 _6082_ (.CLK(clknet_leaf_21_clk),
    .D(_0108_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[26] ));
 sky130_fd_sc_hd__dfrtp_2 _6083_ (.CLK(clknet_leaf_23_clk),
    .D(_0109_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[27] ));
 sky130_fd_sc_hd__dfrtp_4 _6084_ (.CLK(clknet_leaf_21_clk),
    .D(_0110_),
    .RESET_B(net189),
    .Q(\ih.t.timer_max[28] ));
 sky130_fd_sc_hd__dfrtp_2 _6085_ (.CLK(clknet_leaf_23_clk),
    .D(_0111_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[29] ));
 sky130_fd_sc_hd__dfrtp_2 _6086_ (.CLK(clknet_leaf_22_clk),
    .D(_0112_),
    .RESET_B(net193),
    .Q(\ih.t.timer_max[30] ));
 sky130_fd_sc_hd__dfrtp_4 _6087_ (.CLK(clknet_leaf_22_clk),
    .D(_0113_),
    .RESET_B(net193),
    .Q(\ih.t.timer_max[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6088_ (.CLK(clknet_leaf_15_clk),
    .D(_0114_),
    .RESET_B(net175),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _6089_ (.CLK(clknet_leaf_11_clk),
    .D(_0115_),
    .RESET_B(net171),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _6090_ (.CLK(clknet_leaf_8_clk),
    .D(_0116_),
    .RESET_B(net172),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_4 _6091_ (.CLK(clknet_leaf_29_clk),
    .D(_0117_),
    .RESET_B(net184),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_4 _6092_ (.CLK(clknet_leaf_24_clk),
    .D(_0118_),
    .RESET_B(net192),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_4 _6093_ (.CLK(clknet_leaf_7_clk),
    .D(_0119_),
    .RESET_B(net166),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_4 _6094_ (.CLK(clknet_leaf_27_clk),
    .D(_0120_),
    .RESET_B(net184),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_4 _6095_ (.CLK(clknet_leaf_27_clk),
    .D(_0121_),
    .RESET_B(net184),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_2 _6096_ (.CLK(clknet_leaf_20_clk),
    .D(_0122_),
    .RESET_B(net188),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _6097_ (.CLK(clknet_leaf_9_clk),
    .D(_0123_),
    .RESET_B(net172),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_4 _6098_ (.CLK(clknet_leaf_27_clk),
    .D(_0124_),
    .RESET_B(net184),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _6099_ (.CLK(clknet_leaf_6_clk),
    .D(_0125_),
    .RESET_B(net162),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_2 _6100_ (.CLK(clknet_leaf_6_clk),
    .D(_0126_),
    .RESET_B(net162),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_4 _6101_ (.CLK(clknet_leaf_26_clk),
    .D(_0127_),
    .RESET_B(net192),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_4 _6102_ (.CLK(clknet_leaf_5_clk),
    .D(_0128_),
    .RESET_B(net163),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_2 _6103_ (.CLK(clknet_leaf_5_clk),
    .D(_0129_),
    .RESET_B(net163),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_4 _6104_ (.CLK(clknet_leaf_39_clk),
    .D(_0130_),
    .RESET_B(net151),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_4 _6105_ (.CLK(clknet_leaf_26_clk),
    .D(_0131_),
    .RESET_B(net192),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_2 _6106_ (.CLK(clknet_leaf_8_clk),
    .D(_0132_),
    .RESET_B(net172),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_4 _6107_ (.CLK(clknet_leaf_36_clk),
    .D(_0133_),
    .RESET_B(net161),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_2 _6108_ (.CLK(clknet_leaf_6_clk),
    .D(_0134_),
    .RESET_B(net162),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_4 _6109_ (.CLK(clknet_leaf_5_clk),
    .D(_0135_),
    .RESET_B(net163),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_4 _6110_ (.CLK(clknet_leaf_27_clk),
    .D(_0136_),
    .RESET_B(net185),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_2 _6111_ (.CLK(clknet_leaf_26_clk),
    .D(_0137_),
    .RESET_B(net192),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _6112_ (.CLK(clknet_leaf_26_clk),
    .D(_0138_),
    .RESET_B(net192),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _6113_ (.CLK(clknet_leaf_26_clk),
    .D(_0139_),
    .RESET_B(net193),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _6114_ (.CLK(clknet_leaf_7_clk),
    .D(_0140_),
    .RESET_B(net165),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _6115_ (.CLK(clknet_leaf_27_clk),
    .D(_0141_),
    .RESET_B(net185),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _6116_ (.CLK(clknet_leaf_7_clk),
    .D(_0142_),
    .RESET_B(net165),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_2 _6117_ (.CLK(clknet_leaf_27_clk),
    .D(_0143_),
    .RESET_B(net185),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _6118_ (.CLK(clknet_leaf_26_clk),
    .D(_0144_),
    .RESET_B(net193),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _6119_ (.CLK(clknet_leaf_27_clk),
    .D(_0145_),
    .RESET_B(net185),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _6120_ (.CLK(clknet_leaf_19_clk),
    .D(_0146_),
    .RESET_B(net188),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _6121_ (.CLK(clknet_leaf_9_clk),
    .D(_0147_),
    .RESET_B(net172),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 _6122_ (.CLK(clknet_leaf_6_clk),
    .D(_0148_),
    .RESET_B(net165),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_2 _6123_ (.CLK(clknet_leaf_6_clk),
    .D(_0149_),
    .RESET_B(net165),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _6124_ (.CLK(clknet_leaf_7_clk),
    .D(_0150_),
    .RESET_B(net165),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 _6125_ (.CLK(clknet_leaf_19_clk),
    .D(_0151_),
    .RESET_B(net183),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _6126_ (.CLK(clknet_leaf_8_clk),
    .D(_0152_),
    .RESET_B(net172),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_2 _6127_ (.CLK(clknet_leaf_11_clk),
    .D(_0153_),
    .RESET_B(net171),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_2 _6128_ (.CLK(clknet_leaf_14_clk),
    .D(_0154_),
    .RESET_B(net175),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _6129_ (.CLK(clknet_leaf_8_clk),
    .D(_0155_),
    .RESET_B(net172),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _6130_ (.CLK(clknet_leaf_7_clk),
    .D(_0156_),
    .RESET_B(net165),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _6131_ (.CLK(clknet_leaf_6_clk),
    .D(_0157_),
    .RESET_B(net165),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _6132_ (.CLK(clknet_leaf_18_clk),
    .D(_0158_),
    .RESET_B(net182),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_2 _6133_ (.CLK(clknet_leaf_16_clk),
    .D(_0159_),
    .RESET_B(net182),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _6134_ (.CLK(clknet_leaf_16_clk),
    .D(_0160_),
    .RESET_B(net170),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_4 _6135_ (.CLK(clknet_leaf_14_clk),
    .D(_0161_),
    .RESET_B(net175),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _6136_ (.CLK(clknet_leaf_26_clk),
    .D(_0162_),
    .RESET_B(net193),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_2 _6137_ (.CLK(clknet_leaf_8_clk),
    .D(_0163_),
    .RESET_B(net172),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_2 _6138_ (.CLK(clknet_leaf_6_clk),
    .D(_0164_),
    .RESET_B(net162),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_2 _6139_ (.CLK(clknet_leaf_5_clk),
    .D(_0165_),
    .RESET_B(net163),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _6140_ (.CLK(clknet_leaf_5_clk),
    .D(_0166_),
    .RESET_B(net162),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_2 _6141_ (.CLK(clknet_leaf_6_clk),
    .D(_0167_),
    .RESET_B(net162),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_2 _6142_ (.CLK(clknet_leaf_27_clk),
    .D(_0168_),
    .RESET_B(net185),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_4 _6143_ (.CLK(clknet_leaf_16_clk),
    .D(_0169_),
    .RESET_B(net182),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_2 _6144_ (.CLK(clknet_leaf_14_clk),
    .D(_0170_),
    .RESET_B(net178),
    .Q(net132));
 sky130_fd_sc_hd__dfrtp_4 _6145_ (.CLK(clknet_leaf_8_clk),
    .D(_0171_),
    .RESET_B(net171),
    .Q(net133));
 sky130_fd_sc_hd__dfrtp_1 _6146_ (.CLK(clknet_leaf_8_clk),
    .D(_0172_),
    .RESET_B(net172),
    .Q(net134));
 sky130_fd_sc_hd__dfrtp_2 _6147_ (.CLK(clknet_leaf_5_clk),
    .D(_0173_),
    .RESET_B(net162),
    .Q(net135));
 sky130_fd_sc_hd__dfrtp_4 _6148_ (.CLK(clknet_leaf_6_clk),
    .D(_0174_),
    .RESET_B(net162),
    .Q(net136));
 sky130_fd_sc_hd__dfrtp_1 _6149_ (.CLK(clknet_leaf_6_clk),
    .D(_0175_),
    .RESET_B(net162),
    .Q(net137));
 sky130_fd_sc_hd__dfrtp_2 _6150_ (.CLK(clknet_leaf_7_clk),
    .D(_0176_),
    .RESET_B(net166),
    .Q(net138));
 sky130_fd_sc_hd__dfrtp_4 _6151_ (.CLK(clknet_leaf_16_clk),
    .D(_0177_),
    .RESET_B(net170),
    .Q(net139));
 sky130_fd_sc_hd__dfrtp_4 _6152_ (.CLK(clknet_leaf_16_clk),
    .D(_0178_),
    .RESET_B(net170),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_4 _6153_ (.CLK(clknet_leaf_7_clk),
    .D(_0179_),
    .RESET_B(net166),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_4 _6154_ (.CLK(clknet_leaf_8_clk),
    .D(_0180_),
    .RESET_B(net171),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_4 _6155_ (.CLK(clknet_leaf_7_clk),
    .D(_0181_),
    .RESET_B(net166),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_4 _6156_ (.CLK(clknet_leaf_11_clk),
    .D(_0182_),
    .RESET_B(net171),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_4 _6157_ (.CLK(clknet_leaf_11_clk),
    .D(_0183_),
    .RESET_B(net171),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_4 _6158_ (.CLK(clknet_leaf_8_clk),
    .D(_0184_),
    .RESET_B(net172),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_2 _6159_ (.CLK(clknet_leaf_7_clk),
    .D(_0185_),
    .RESET_B(net166),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _6160_ (.CLK(clknet_leaf_16_clk),
    .D(_0186_),
    .RESET_B(net170),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_4 _6161_ (.CLK(clknet_leaf_16_clk),
    .D(_0187_),
    .RESET_B(net170),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_4 _6162_ (.CLK(clknet_leaf_4_clk),
    .D(_0188_),
    .RESET_B(net167),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_4 _6163_ (.CLK(clknet_leaf_4_clk),
    .D(_0189_),
    .RESET_B(net167),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_4 _6164_ (.CLK(clknet_leaf_4_clk),
    .D(_0190_),
    .RESET_B(net167),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _6165_ (.CLK(clknet_leaf_6_clk),
    .D(_0191_),
    .RESET_B(net165),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_4 _6166_ (.CLK(clknet_leaf_6_clk),
    .D(_0192_),
    .RESET_B(net162),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_2 _6167_ (.CLK(clknet_leaf_6_clk),
    .D(_0193_),
    .RESET_B(net164),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_2 _6168_ (.CLK(clknet_leaf_40_clk),
    .D(_0194_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6169_ (.CLK(clknet_leaf_40_clk),
    .D(_0195_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6170_ (.CLK(clknet_leaf_40_clk),
    .D(_0196_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6171_ (.CLK(clknet_leaf_0_clk),
    .D(_0197_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_mem[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6172_ (.CLK(clknet_leaf_40_clk),
    .D(_0198_),
    .RESET_B(net156),
    .Q(\cu.reg_file.reg_mem[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6173_ (.CLK(clknet_leaf_0_clk),
    .D(_0199_),
    .RESET_B(net154),
    .Q(\cu.reg_file.reg_mem[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6174_ (.CLK(clknet_leaf_2_clk),
    .D(_0200_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_mem[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6175_ (.CLK(clknet_leaf_2_clk),
    .D(_0201_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_mem[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6176_ (.CLK(clknet_leaf_19_clk),
    .D(_0202_),
    .RESET_B(net183),
    .Q(\cu.reg_file.reg_mem[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6177_ (.CLK(clknet_leaf_18_clk),
    .D(_0203_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6178_ (.CLK(clknet_leaf_18_clk),
    .D(_0204_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6179_ (.CLK(clknet_leaf_18_clk),
    .D(_0205_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6180_ (.CLK(clknet_leaf_18_clk),
    .D(_0206_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6181_ (.CLK(clknet_leaf_18_clk),
    .D(_0207_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6182_ (.CLK(clknet_leaf_18_clk),
    .D(_0208_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6183_ (.CLK(clknet_leaf_18_clk),
    .D(_0209_),
    .RESET_B(net182),
    .Q(\cu.reg_file.reg_mem[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6184_ (.CLK(clknet_leaf_39_clk),
    .D(_0000_),
    .RESET_B(net151),
    .Q(\ih.interrupt_source[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6185_ (.CLK(clknet_leaf_4_clk),
    .D(_0210_),
    .RESET_B(net167),
    .Q(\ih.input_handler_enable ));
 sky130_fd_sc_hd__dfrtp_4 _6186_ (.CLK(clknet_leaf_23_clk),
    .D(_0211_),
    .RESET_B(net188),
    .Q(\mc.count ));
 sky130_fd_sc_hd__dfrtp_1 _6187_ (.CLK(clknet_leaf_39_clk),
    .D(net200),
    .RESET_B(net151),
    .Q(\ih.interrupt_source[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6188_ (.CLK(clknet_leaf_39_clk),
    .D(_0213_),
    .RESET_B(net151),
    .Q(\ih.interrupt_source[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6189_ (.CLK(clknet_leaf_19_clk),
    .D(_0214_),
    .RESET_B(net188),
    .Q(\mc.cl.next_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6190_ (.CLK(clknet_leaf_20_clk),
    .D(_0215_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6191_ (.CLK(clknet_leaf_20_clk),
    .D(_0216_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6192_ (.CLK(clknet_leaf_20_clk),
    .D(_0217_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6193_ (.CLK(clknet_leaf_20_clk),
    .D(_0218_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6194_ (.CLK(clknet_leaf_23_clk),
    .D(_0219_),
    .RESET_B(net188),
    .Q(\mc.cl.next_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6195_ (.CLK(clknet_leaf_14_clk),
    .D(_0220_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6196_ (.CLK(clknet_leaf_20_clk),
    .D(_0221_),
    .RESET_B(net187),
    .Q(\mc.cl.next_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6197_ (.CLK(clknet_leaf_24_clk),
    .D(net215),
    .RESET_B(net192),
    .Q(\mc.cc.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _6198_ (.CLK(clknet_leaf_24_clk),
    .D(_0223_),
    .SET_B(net193),
    .Q(\mc.cc.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6199_ (.CLK(clknet_leaf_24_clk),
    .D(net211),
    .RESET_B(net193),
    .Q(\mc.cc.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6200_ (.CLK(clknet_leaf_24_clk),
    .D(_0225_),
    .RESET_B(net193),
    .Q(\mc.cc.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6201_ (.CLK(clknet_leaf_39_clk),
    .D(net1),
    .RESET_B(net151),
    .Q(\ih.ip_ed.prev_data ));
 sky130_fd_sc_hd__dfrtp_1 _6202_ (.CLK(clknet_leaf_4_clk),
    .D(net2),
    .RESET_B(net167),
    .Q(\ih.ih.ih.prev_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6203_ (.CLK(clknet_leaf_5_clk),
    .D(net9),
    .RESET_B(net164),
    .Q(\ih.ih.ih.prev_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6204_ (.CLK(clknet_leaf_7_clk),
    .D(net10),
    .RESET_B(net165),
    .Q(\ih.ih.ih.prev_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6205_ (.CLK(clknet_leaf_7_clk),
    .D(net11),
    .RESET_B(net165),
    .Q(\ih.ih.ih.prev_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6206_ (.CLK(clknet_leaf_5_clk),
    .D(net12),
    .RESET_B(net163),
    .Q(\ih.ih.ih.prev_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6207_ (.CLK(clknet_leaf_5_clk),
    .D(net13),
    .RESET_B(net163),
    .Q(\ih.ih.ih.prev_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6208_ (.CLK(clknet_leaf_4_clk),
    .D(net14),
    .RESET_B(net163),
    .Q(\ih.ih.ih.prev_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6209_ (.CLK(clknet_leaf_4_clk),
    .D(net15),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6210_ (.CLK(clknet_leaf_4_clk),
    .D(net16),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6211_ (.CLK(clknet_leaf_5_clk),
    .D(net17),
    .RESET_B(net163),
    .Q(\ih.ih.ih.prev_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6212_ (.CLK(clknet_leaf_5_clk),
    .D(net3),
    .RESET_B(net163),
    .Q(\ih.ih.ih.prev_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6213_ (.CLK(clknet_leaf_6_clk),
    .D(net4),
    .RESET_B(net164),
    .Q(\ih.ih.ih.prev_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6214_ (.CLK(clknet_leaf_5_clk),
    .D(net5),
    .RESET_B(net164),
    .Q(\ih.ih.ih.prev_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6215_ (.CLK(clknet_leaf_5_clk),
    .D(net6),
    .RESET_B(net164),
    .Q(\ih.ih.ih.prev_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6216_ (.CLK(clknet_leaf_4_clk),
    .D(net7),
    .RESET_B(net164),
    .Q(\ih.ih.ih.prev_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6217_ (.CLK(clknet_leaf_4_clk),
    .D(net8),
    .RESET_B(net168),
    .Q(\ih.ih.ih.prev_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6218_ (.CLK(clknet_leaf_4_clk),
    .D(\ih.ih.int_f.data_in ),
    .RESET_B(net168),
    .Q(\ih.ih.int_f.prev_data ));
 sky130_fd_sc_hd__dfrtp_4 _6219_ (.CLK(clknet_leaf_9_clk),
    .D(\ih.t.next_count[0] ),
    .RESET_B(net173),
    .Q(\ih.t.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6220_ (.CLK(clknet_leaf_9_clk),
    .D(\ih.t.next_count[1] ),
    .RESET_B(net173),
    .Q(\ih.t.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6221_ (.CLK(clknet_leaf_9_clk),
    .D(\ih.t.next_count[2] ),
    .RESET_B(net173),
    .Q(\ih.t.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6222_ (.CLK(clknet_leaf_9_clk),
    .D(\ih.t.next_count[3] ),
    .RESET_B(net173),
    .Q(\ih.t.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6223_ (.CLK(clknet_leaf_9_clk),
    .D(\ih.t.next_count[4] ),
    .RESET_B(net173),
    .Q(\ih.t.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6224_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[5] ),
    .RESET_B(net173),
    .Q(\ih.t.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6225_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[6] ),
    .RESET_B(net173),
    .Q(\ih.t.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6226_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[7] ),
    .RESET_B(net173),
    .Q(\ih.t.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6227_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[8] ),
    .RESET_B(net173),
    .Q(\ih.t.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6228_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[9] ),
    .RESET_B(net173),
    .Q(\ih.t.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6229_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[10] ),
    .RESET_B(net174),
    .Q(\ih.t.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6230_ (.CLK(clknet_leaf_10_clk),
    .D(\ih.t.next_count[11] ),
    .RESET_B(net174),
    .Q(\ih.t.count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6231_ (.CLK(clknet_leaf_12_clk),
    .D(\ih.t.next_count[12] ),
    .RESET_B(net176),
    .Q(\ih.t.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6232_ (.CLK(clknet_leaf_12_clk),
    .D(\ih.t.next_count[13] ),
    .RESET_B(net176),
    .Q(\ih.t.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6233_ (.CLK(clknet_leaf_12_clk),
    .D(\ih.t.next_count[14] ),
    .RESET_B(net176),
    .Q(\ih.t.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6234_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[15] ),
    .RESET_B(net176),
    .Q(\ih.t.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6235_ (.CLK(clknet_leaf_12_clk),
    .D(\ih.t.next_count[16] ),
    .RESET_B(net176),
    .Q(\ih.t.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6236_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[17] ),
    .RESET_B(net176),
    .Q(\ih.t.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6237_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[18] ),
    .RESET_B(net177),
    .Q(\ih.t.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6238_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[19] ),
    .RESET_B(net177),
    .Q(\ih.t.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6239_ (.CLK(clknet_leaf_13_clk),
    .D(\ih.t.next_count[20] ),
    .RESET_B(net177),
    .Q(\ih.t.count[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6240_ (.CLK(clknet_leaf_21_clk),
    .D(\ih.t.next_count[21] ),
    .RESET_B(net189),
    .Q(\ih.t.count[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6241_ (.CLK(clknet_leaf_21_clk),
    .D(\ih.t.next_count[22] ),
    .RESET_B(net189),
    .Q(\ih.t.count[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6242_ (.CLK(clknet_leaf_21_clk),
    .D(\ih.t.next_count[23] ),
    .RESET_B(net189),
    .Q(\ih.t.count[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6243_ (.CLK(clknet_leaf_21_clk),
    .D(\ih.t.next_count[24] ),
    .RESET_B(net191),
    .Q(\ih.t.count[24] ));
 sky130_fd_sc_hd__dfrtp_2 _6244_ (.CLK(clknet_leaf_22_clk),
    .D(\ih.t.next_count[25] ),
    .RESET_B(net190),
    .Q(\ih.t.count[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6245_ (.CLK(clknet_leaf_22_clk),
    .D(\ih.t.next_count[26] ),
    .RESET_B(net190),
    .Q(\ih.t.count[26] ));
 sky130_fd_sc_hd__dfrtp_1 _6246_ (.CLK(clknet_leaf_22_clk),
    .D(\ih.t.next_count[27] ),
    .RESET_B(net191),
    .Q(\ih.t.count[27] ));
 sky130_fd_sc_hd__dfrtp_2 _6247_ (.CLK(clknet_leaf_22_clk),
    .D(\ih.t.next_count[28] ),
    .RESET_B(net191),
    .Q(\ih.t.count[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6248_ (.CLK(clknet_leaf_22_clk),
    .D(\ih.t.next_count[29] ),
    .RESET_B(net191),
    .Q(\ih.t.count[29] ));
 sky130_fd_sc_hd__dfrtp_1 _6249_ (.CLK(clknet_leaf_25_clk),
    .D(\ih.t.next_count[30] ),
    .RESET_B(net193),
    .Q(\ih.t.count[30] ));
 sky130_fd_sc_hd__dfrtp_1 _6250_ (.CLK(clknet_leaf_25_clk),
    .D(\ih.t.next_count[31] ),
    .RESET_B(net194),
    .Q(\ih.t.count[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6251_ (.CLK(clknet_leaf_39_clk),
    .D(_0015_),
    .RESET_B(net151),
    .Q(\cu.id.interrupt_requested ));
 sky130_fd_sc_hd__dfrtp_4 _6252_ (.CLK(clknet_leaf_2_clk),
    .D(_0226_),
    .RESET_B(net157),
    .Q(\cu.reg_file.reg_sp[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6253_ (.CLK(clknet_leaf_37_clk),
    .D(_0227_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_sp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6254_ (.CLK(clknet_leaf_3_clk),
    .D(_0228_),
    .RESET_B(net158),
    .Q(\cu.reg_file.reg_sp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6255_ (.CLK(clknet_leaf_3_clk),
    .D(_0229_),
    .RESET_B(net169),
    .Q(\cu.reg_file.reg_sp[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6256_ (.CLK(clknet_leaf_3_clk),
    .D(_0230_),
    .RESET_B(net169),
    .Q(\cu.reg_file.reg_sp[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6257_ (.CLK(clknet_leaf_17_clk),
    .D(_0231_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_sp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6258_ (.CLK(clknet_leaf_17_clk),
    .D(_0232_),
    .RESET_B(net180),
    .Q(\cu.reg_file.reg_sp[7] ));
 sky130_fd_sc_hd__dfstp_2 _6259_ (.CLK(clknet_leaf_37_clk),
    .D(_0233_),
    .SET_B(net158),
    .Q(\cu.reg_file.reg_sp[8] ));
 sky130_fd_sc_hd__dfstp_2 _6260_ (.CLK(clknet_leaf_37_clk),
    .D(_0234_),
    .SET_B(net158),
    .Q(\cu.reg_file.reg_sp[9] ));
 sky130_fd_sc_hd__dfstp_2 _6261_ (.CLK(clknet_leaf_34_clk),
    .D(_0235_),
    .SET_B(net159),
    .Q(\cu.reg_file.reg_sp[10] ));
 sky130_fd_sc_hd__dfstp_2 _6262_ (.CLK(clknet_leaf_34_clk),
    .D(_0236_),
    .SET_B(net159),
    .Q(\cu.reg_file.reg_sp[11] ));
 sky130_fd_sc_hd__dfstp_2 _6263_ (.CLK(clknet_leaf_34_clk),
    .D(_0237_),
    .SET_B(net159),
    .Q(\cu.reg_file.reg_sp[12] ));
 sky130_fd_sc_hd__dfstp_2 _6264_ (.CLK(clknet_leaf_34_clk),
    .D(_0238_),
    .SET_B(net159),
    .Q(\cu.reg_file.reg_sp[13] ));
 sky130_fd_sc_hd__dfstp_2 _6265_ (.CLK(clknet_leaf_35_clk),
    .D(_0239_),
    .SET_B(net160),
    .Q(\cu.reg_file.reg_sp[14] ));
 sky130_fd_sc_hd__dfstp_2 _6266_ (.CLK(clknet_leaf_35_clk),
    .D(_0240_),
    .SET_B(net160),
    .Q(\cu.reg_file.reg_sp[15] ));
 sky130_fd_sc_hd__dfstp_2 _6267_ (.CLK(clknet_leaf_21_clk),
    .D(_0241_),
    .SET_B(net189),
    .Q(\ih.t.timer_max[8] ));
 sky130_fd_sc_hd__dfstp_1 _6268_ (.CLK(clknet_leaf_14_clk),
    .D(_0242_),
    .SET_B(net189),
    .Q(\ih.t.timer_max[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6269_ (.CLK(clknet_leaf_21_clk),
    .D(_0243_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6270_ (.CLK(clknet_leaf_21_clk),
    .D(_0244_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[11] ));
 sky130_fd_sc_hd__dfrtp_2 _6271_ (.CLK(clknet_leaf_21_clk),
    .D(_0245_),
    .RESET_B(net191),
    .Q(\ih.t.timer_max[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6272_ (.CLK(clknet_leaf_22_clk),
    .D(_0246_),
    .RESET_B(net190),
    .Q(\ih.t.timer_max[13] ));
 sky130_fd_sc_hd__dfstp_2 _6273_ (.CLK(clknet_leaf_23_clk),
    .D(_0247_),
    .SET_B(net190),
    .Q(\ih.t.timer_max[14] ));
 sky130_fd_sc_hd__dfstp_2 _6274_ (.CLK(clknet_leaf_24_clk),
    .D(_0248_),
    .SET_B(net192),
    .Q(\ih.t.timer_max[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6275_ (.CLK(clknet_leaf_8_clk),
    .D(_0249_),
    .RESET_B(net171),
    .Q(\ih.t.timer_max[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6276_ (.CLK(clknet_leaf_11_clk),
    .D(_0250_),
    .RESET_B(net174),
    .Q(\ih.t.timer_max[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6277_ (.CLK(clknet_leaf_11_clk),
    .D(_0251_),
    .RESET_B(net171),
    .Q(\ih.t.timer_max[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6278_ (.CLK(clknet_leaf_11_clk),
    .D(_0252_),
    .RESET_B(net174),
    .Q(\ih.t.timer_max[3] ));
 sky130_fd_sc_hd__dfstp_1 _6279_ (.CLK(clknet_leaf_12_clk),
    .D(_0253_),
    .SET_B(net176),
    .Q(\ih.t.timer_max[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6280_ (.CLK(clknet_leaf_11_clk),
    .D(_0254_),
    .RESET_B(net174),
    .Q(\ih.t.timer_max[5] ));
 sky130_fd_sc_hd__dfstp_1 _6281_ (.CLK(clknet_leaf_11_clk),
    .D(_0255_),
    .SET_B(net175),
    .Q(\ih.t.timer_max[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6282_ (.CLK(clknet_leaf_11_clk),
    .D(_0256_),
    .RESET_B(net179),
    .Q(\ih.t.timer_max[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6283_ (.CLK(clknet_leaf_11_clk),
    .D(_0257_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[16] ));
 sky130_fd_sc_hd__dfrtp_2 _6284_ (.CLK(clknet_leaf_11_clk),
    .D(_0258_),
    .RESET_B(net176),
    .Q(\ih.t.timer_max[17] ));
 sky130_fd_sc_hd__dfrtp_2 _6285_ (.CLK(clknet_leaf_11_clk),
    .D(_0259_),
    .RESET_B(net175),
    .Q(\ih.t.timer_max[18] ));
 sky130_fd_sc_hd__dfrtp_2 _6286_ (.CLK(clknet_leaf_12_clk),
    .D(_0260_),
    .RESET_B(net176),
    .Q(\ih.t.timer_max[19] ));
 sky130_fd_sc_hd__dfrtp_2 _6287_ (.CLK(clknet_leaf_12_clk),
    .D(_0261_),
    .RESET_B(net176),
    .Q(\ih.t.timer_max[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6288_ (.CLK(clknet_leaf_13_clk),
    .D(_0262_),
    .RESET_B(net177),
    .Q(\ih.t.timer_max[21] ));
 sky130_fd_sc_hd__dfrtp_4 _6289_ (.CLK(clknet_leaf_14_clk),
    .D(_0263_),
    .RESET_B(net177),
    .Q(\ih.t.timer_max[22] ));
 sky130_fd_sc_hd__dfrtp_2 _6290_ (.CLK(clknet_leaf_14_clk),
    .D(_0264_),
    .RESET_B(net178),
    .Q(\ih.t.timer_max[23] ));
 sky130_fd_sc_hd__dfrtp_2 _6291_ (.CLK(clknet_leaf_0_clk),
    .D(_0265_),
    .RESET_B(net154),
    .Q(\cu.ir.idx[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6292_ (.CLK(clknet_leaf_1_clk),
    .D(_0266_),
    .RESET_B(net154),
    .Q(\cu.ir.idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6293_ (.CLK(clknet_leaf_39_clk),
    .D(_0267_),
    .RESET_B(net151),
    .Q(\cu.id.can_be_interrupted ));
 sky130_fd_sc_hd__dfrtp_4 _6294_ (.CLK(clknet_leaf_40_clk),
    .D(_0268_),
    .RESET_B(net156),
    .Q(\cu.id.opcode[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6295_ (.CLK(clknet_leaf_40_clk),
    .D(_0269_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6296_ (.CLK(clknet_leaf_40_clk),
    .D(_0270_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6297_ (.CLK(clknet_leaf_40_clk),
    .D(_0271_),
    .RESET_B(net156),
    .Q(\cu.id.alu_opcode[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6298_ (.CLK(clknet_leaf_40_clk),
    .D(_0272_),
    .RESET_B(net156),
    .Q(\cu.id.alu_opcode[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6299_ (.CLK(clknet_leaf_40_clk),
    .D(_0273_),
    .RESET_B(net156),
    .Q(\cu.id.alu_opcode[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6300_ (.CLK(clknet_leaf_40_clk),
    .D(_0274_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6301_ (.CLK(clknet_leaf_40_clk),
    .D(_0275_),
    .RESET_B(net153),
    .Q(\cu.id.opcode[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6302_ (.CLK(clknet_leaf_0_clk),
    .D(_0276_),
    .RESET_B(net155),
    .Q(\cu.id.cb_opcode_z[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6303_ (.CLK(clknet_leaf_0_clk),
    .D(_0277_),
    .RESET_B(net155),
    .Q(\cu.id.cb_opcode_z[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6304_ (.CLK(clknet_leaf_0_clk),
    .D(_0278_),
    .RESET_B(net155),
    .Q(\cu.id.cb_opcode_z[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6305_ (.CLK(clknet_leaf_0_clk),
    .D(_0279_),
    .RESET_B(net155),
    .Q(\cu.id.cb_opcode_y[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6306_ (.CLK(clknet_leaf_1_clk),
    .D(_0280_),
    .RESET_B(net155),
    .Q(\cu.id.cb_opcode_y[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6307_ (.CLK(clknet_leaf_2_clk),
    .D(_0281_),
    .RESET_B(net157),
    .Q(\cu.id.cb_opcode_y[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6308_ (.CLK(clknet_leaf_2_clk),
    .D(_0282_),
    .RESET_B(net157),
    .Q(\cu.id.cb_opcode_x[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6309_ (.CLK(clknet_leaf_3_clk),
    .D(_0283_),
    .RESET_B(net167),
    .Q(\cu.id.cb_opcode_x[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6310_ (.CLK(clknet_leaf_0_clk),
    .D(_0284_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6311_ (.CLK(clknet_leaf_0_clk),
    .D(_0285_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6312_ (.CLK(clknet_leaf_0_clk),
    .D(_0286_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6313_ (.CLK(clknet_leaf_0_clk),
    .D(_0287_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6314_ (.CLK(clknet_leaf_0_clk),
    .D(_0288_),
    .RESET_B(net155),
    .Q(\cu.id.imm_i[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6315_ (.CLK(clknet_leaf_0_clk),
    .D(_0289_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6316_ (.CLK(clknet_leaf_0_clk),
    .D(_0290_),
    .RESET_B(net154),
    .Q(\cu.id.imm_i[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6317_ (.CLK(clknet_leaf_0_clk),
    .D(_0291_),
    .RESET_B(net155),
    .Q(\cu.id.imm_i[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6318_ (.CLK(clknet_leaf_1_clk),
    .D(_0004_),
    .RESET_B(net155),
    .Q(\cu.id.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6319_ (.CLK(clknet_leaf_1_clk),
    .D(_0005_),
    .RESET_B(net155),
    .Q(\cu.id.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6320_ (.CLK(clknet_leaf_5_clk),
    .D(_0006_),
    .RESET_B(net163),
    .Q(\cu.id.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6321_ (.CLK(clknet_leaf_39_clk),
    .D(_0001_),
    .RESET_B(net153),
    .Q(\cu.id.is_halted ));
 sky130_fd_sc_hd__dfrtp_4 _6322_ (.CLK(clknet_leaf_39_clk),
    .D(_0003_),
    .RESET_B(net153),
    .Q(\cu.id.starting_int_service ));
 sky130_fd_sc_hd__dfrtp_1 _6323_ (.CLK(clknet_leaf_39_clk),
    .D(_0002_),
    .RESET_B(net153),
    .Q(\cu.id.is_interrupted ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net197),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net197),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(net197),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net197),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net196),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net196),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net170),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net196),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net179),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net179),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(net179),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net178),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 fanout179 (.A(net196),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net183),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 fanout183 (.A(net195),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(net195),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net195),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net195),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net194),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net194),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net194),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net26),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 hold1 (.A(\cu.id.is_halted ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\cu.alu_f[3] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\cu.alu_f[4] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\cu.alu_f[5] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\mc.cc.count[3] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0224_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\ih.t.count[16] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\ih.t.count[10] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\mc.cc.count[0] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0222_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ih.t.count[22] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\ih.ip_ed.prev_data ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\ih.t.count[25] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ih.t.count[13] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\ih.t.count[28] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\ih.t.count[4] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\ih.t.count[19] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\cu.ir.idx[0] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\ih.t.count[7] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\ih.t.count[9] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\ih.ih.ih.prev_data[11] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_2717_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0212_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\mc.cc.count[1] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\ih.t.count[18] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\ih.t.count[24] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ih.t.count[27] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\ih.t.count[21] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\ih.t.count[15] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\ih.input_handler_enable ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ih.t.count[8] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\ih.t.count[6] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\cu.ir.idx[1] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\cu.id.interrupt_requested ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\cu.id.can_be_interrupted ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\cu.id.is_interrupted ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ih.interrupt_source[1] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\ih.interrupt_source[2] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\ih.t.count[30] ),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(interrupt_gpio_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(keypad_input[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(keypad_input[3]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(keypad_input[4]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(keypad_input[5]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(keypad_input[6]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(keypad_input[7]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(keypad_input[8]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(keypad_input[9]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(memory_data_in[0]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(memory_data_in[1]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(keypad_input[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(memory_data_in[2]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(memory_data_in[3]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(memory_data_in[4]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(memory_data_in[5]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(memory_data_in[6]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(memory_data_in[7]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(nrst),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(programmable_gpio_in[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(programmable_gpio_in[1]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(programmable_gpio_in[2]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(keypad_input[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(programmable_gpio_in[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(programmable_gpio_in[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(programmable_gpio_in[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(programmable_gpio_in[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(programmable_gpio_in[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input4 (.A(keypad_input[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(keypad_input[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(keypad_input[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(keypad_input[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(keypad_input[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(keypad_input[1]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap141 (.A(_2321_),
    .X(net141));
 sky130_fd_sc_hd__buf_2 max_cap142 (.A(_0510_),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap145 (.A(net239),
    .X(net145));
 sky130_fd_sc_hd__buf_1 max_cap146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 max_cap147 (.A(net240),
    .X(net147));
 sky130_fd_sc_hd__buf_1 max_cap149 (.A(_1654_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 max_cap150 (.A(_2898_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(ss3[0]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(ss3[1]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(ss3[2]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(ss3[3]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(ss3[4]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(ss3[5]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(ss3[6]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(ss3[7]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(ss4[0]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(ss4[1]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(ss4[2]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(ss4[3]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(ss4[4]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(ss4[5]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(ss4[6]));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(ss4[7]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(ss5[0]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(ss5[1]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(ss5[2]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(ss5[3]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(ss5[4]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(ss5[5]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(ss5[6]));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net123),
    .X(ss5[7]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(ss6[0]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(ss6[1]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(ss6[2]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(ss6[3]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(ss6[4]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(ss6[5]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(ss6[6]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(ss6[7]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(ss7[0]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(ss7[1]));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net134),
    .X(ss7[2]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(ss7[3]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(ss7[4]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(ss7[5]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(ss7[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(ss7[7]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(memory_address_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(memory_address_out[10]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(memory_address_out[11]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(memory_address_out[12]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(memory_address_out[13]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(memory_address_out[14]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(memory_address_out[15]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(memory_address_out[1]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(memory_address_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(memory_address_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .X(memory_address_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(memory_address_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(memory_address_out[6]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(memory_address_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(memory_address_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(memory_address_out[9]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(memory_data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(memory_data_out[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(memory_data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(memory_data_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(memory_data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(memory_data_out[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(memory_data_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(memory_data_out[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(memory_wr));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(programmable_gpio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(programmable_gpio_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(programmable_gpio_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(programmable_gpio_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(programmable_gpio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(programmable_gpio_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(programmable_gpio_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(programmable_gpio_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(programmable_gpio_wr[0]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(programmable_gpio_wr[1]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(programmable_gpio_wr[2]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(programmable_gpio_wr[3]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(programmable_gpio_wr[4]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(programmable_gpio_wr[5]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(programmable_gpio_wr[6]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(programmable_gpio_wr[7]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(ss0[0]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(ss0[1]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(ss0[2]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(ss0[3]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(ss0[4]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(ss0[5]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(ss0[6]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(ss0[7]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(ss1[0]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(ss1[1]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(ss1[2]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(ss1[3]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(ss1[4]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(ss1[5]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(ss1[6]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(ss1[7]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(ss2[0]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(ss2[1]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(ss2[2]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(ss2[3]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(ss2[4]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(ss2[5]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(ss2[6]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(ss2[7]));
 sky130_fd_sc_hd__buf_1 wire1 (.A(_0985_),
    .X(net237));
 sky130_fd_sc_hd__buf_4 wire140 (.A(_1811_),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire144 (.A(_1279_),
    .X(net144));
 sky130_fd_sc_hd__buf_1 wire148 (.A(net241),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 wire3 (.A(_0482_),
    .X(net239));
 sky130_fd_sc_hd__buf_1 wire4 (.A(_0333_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 wire5 (.A(_0448_),
    .X(net241));
endmodule

