magic
tech sky130A
magscale 1 2
timestamp 1694454425
<< viali >>
rect 1409 45441 1443 45475
rect 6561 45441 6595 45475
rect 14933 45441 14967 45475
rect 23949 45441 23983 45475
rect 32505 45441 32539 45475
rect 41521 45441 41555 45475
rect 1593 45237 1627 45271
rect 6745 45237 6779 45271
rect 15117 45237 15151 45271
rect 24133 45237 24167 45271
rect 32321 45237 32355 45271
rect 41337 45237 41371 45271
rect 5917 44965 5951 44999
rect 18705 44965 18739 44999
rect 31953 44965 31987 44999
rect 36829 44965 36863 44999
rect 5641 44897 5675 44931
rect 11989 44897 12023 44931
rect 16405 44897 16439 44931
rect 18429 44897 18463 44931
rect 18889 44897 18923 44931
rect 10241 44829 10275 44863
rect 12633 44829 12667 44863
rect 13645 44829 13679 44863
rect 15853 44829 15887 44863
rect 16129 44829 16163 44863
rect 19533 44829 19567 44863
rect 10517 44761 10551 44795
rect 14473 44761 14507 44795
rect 31585 44761 31619 44795
rect 36461 44761 36495 44795
rect 6101 44693 6135 44727
rect 12081 44693 12115 44727
rect 13461 44693 13495 44727
rect 14381 44693 14415 44727
rect 16037 44693 16071 44727
rect 17877 44693 17911 44727
rect 19717 44693 19751 44727
rect 32045 44693 32079 44727
rect 36921 44693 36955 44727
rect 10793 44489 10827 44523
rect 11897 44489 11931 44523
rect 16681 44489 16715 44523
rect 8585 44421 8619 44455
rect 13369 44421 13403 44455
rect 18981 44421 19015 44455
rect 20177 44421 20211 44455
rect 6377 44353 6411 44387
rect 8309 44353 8343 44387
rect 10977 44353 11011 44387
rect 17049 44353 17083 44387
rect 18797 44353 18831 44387
rect 19073 44353 19107 44387
rect 19349 44353 19383 44387
rect 31861 44353 31895 44387
rect 36461 44353 36495 44387
rect 11989 44285 12023 44319
rect 12081 44285 12115 44319
rect 12909 44285 12943 44319
rect 13093 44285 13127 44319
rect 14841 44285 14875 44319
rect 15485 44285 15519 44319
rect 17141 44285 17175 44319
rect 17325 44285 17359 44319
rect 19901 44285 19935 44319
rect 11529 44217 11563 44251
rect 12357 44217 12391 44251
rect 6561 44149 6595 44183
rect 8217 44149 8251 44183
rect 8861 44149 8895 44183
rect 14933 44149 14967 44183
rect 18613 44149 18647 44183
rect 19533 44149 19567 44183
rect 21649 44149 21683 44183
rect 31677 44149 31711 44183
rect 36277 44149 36311 44183
rect 12357 43945 12391 43979
rect 14105 43945 14139 43979
rect 17785 43945 17819 43979
rect 15025 43877 15059 43911
rect 6745 43809 6779 43843
rect 14749 43809 14783 43843
rect 15301 43809 15335 43843
rect 17049 43809 17083 43843
rect 17141 43809 17175 43843
rect 18981 43809 19015 43843
rect 21097 43809 21131 43843
rect 25421 43809 25455 43843
rect 31585 43809 31619 43843
rect 36369 43809 36403 43843
rect 10609 43741 10643 43775
rect 13185 43741 13219 43775
rect 13921 43741 13955 43775
rect 14473 43741 14507 43775
rect 14933 43741 14967 43775
rect 18153 43741 18187 43775
rect 19257 43741 19291 43775
rect 21649 43741 21683 43775
rect 31309 43741 31343 43775
rect 36093 43741 36127 43775
rect 7021 43673 7055 43707
rect 10885 43673 10919 43707
rect 15577 43673 15611 43707
rect 19533 43673 19567 43707
rect 43453 43673 43487 43707
rect 44281 43673 44315 43707
rect 8493 43605 8527 43639
rect 12541 43605 12575 43639
rect 13277 43605 13311 43639
rect 14565 43605 14599 43639
rect 18337 43605 18371 43639
rect 18429 43605 18463 43639
rect 21005 43605 21039 43639
rect 26065 43605 26099 43639
rect 33057 43605 33091 43639
rect 37841 43605 37875 43639
rect 11529 43401 11563 43435
rect 14473 43401 14507 43435
rect 15761 43401 15795 43435
rect 17877 43401 17911 43435
rect 19901 43401 19935 43435
rect 20361 43401 20395 43435
rect 10977 43333 11011 43367
rect 13001 43333 13035 43367
rect 29193 43333 29227 43367
rect 10885 43265 10919 43299
rect 11161 43265 11195 43299
rect 12449 43265 12483 43299
rect 17693 43265 17727 43299
rect 17969 43265 18003 43299
rect 21005 43265 21039 43299
rect 28917 43265 28951 43299
rect 33425 43265 33459 43299
rect 11345 43197 11379 43231
rect 12081 43197 12115 43231
rect 12725 43197 12759 43231
rect 15577 43197 15611 43231
rect 16405 43197 16439 43231
rect 17325 43197 17359 43231
rect 18153 43197 18187 43231
rect 18429 43197 18463 43231
rect 20453 43197 20487 43231
rect 20545 43197 20579 43231
rect 24041 43197 24075 43231
rect 36185 43197 36219 43231
rect 38945 43197 38979 43231
rect 39221 43197 39255 43231
rect 17509 43129 17543 43163
rect 19993 43129 20027 43163
rect 24317 43129 24351 43163
rect 12541 43061 12575 43095
rect 15025 43061 15059 43095
rect 16773 43061 16807 43095
rect 20913 43061 20947 43095
rect 24501 43061 24535 43095
rect 30665 43061 30699 43095
rect 34069 43061 34103 43095
rect 35541 43061 35575 43095
rect 40693 43061 40727 43095
rect 12817 42857 12851 42891
rect 13461 42857 13495 42891
rect 16681 42857 16715 42891
rect 39037 42857 39071 42891
rect 6653 42721 6687 42755
rect 12357 42721 12391 42755
rect 12909 42721 12943 42755
rect 18613 42721 18647 42755
rect 19257 42721 19291 42755
rect 38853 42721 38887 42755
rect 40509 42721 40543 42755
rect 5825 42653 5859 42687
rect 9597 42653 9631 42687
rect 9873 42653 9907 42687
rect 10977 42653 11011 42687
rect 11713 42653 11747 42687
rect 12449 42653 12483 42687
rect 12633 42653 12667 42687
rect 13093 42653 13127 42687
rect 13645 42653 13679 42687
rect 13829 42653 13863 42687
rect 13921 42653 13955 42687
rect 14933 42653 14967 42687
rect 21649 42653 21683 42687
rect 24961 42653 24995 42687
rect 34713 42653 34747 42687
rect 38761 42653 38795 42687
rect 39865 42653 39899 42687
rect 40785 42653 40819 42687
rect 13277 42585 13311 42619
rect 15209 42585 15243 42619
rect 18337 42585 18371 42619
rect 21005 42585 21039 42619
rect 34989 42585 35023 42619
rect 8953 42517 8987 42551
rect 9689 42517 9723 42551
rect 10333 42517 10367 42551
rect 16865 42517 16899 42551
rect 21097 42517 21131 42551
rect 25145 42517 25179 42551
rect 36461 42517 36495 42551
rect 40601 42517 40635 42551
rect 10701 42313 10735 42347
rect 14841 42313 14875 42347
rect 15577 42313 15611 42347
rect 16037 42313 16071 42347
rect 17877 42313 17911 42347
rect 27169 42313 27203 42347
rect 38853 42313 38887 42347
rect 42257 42313 42291 42347
rect 9229 42245 9263 42279
rect 15301 42245 15335 42279
rect 25329 42245 25363 42279
rect 33701 42245 33735 42279
rect 35081 42245 35115 42279
rect 36705 42245 36739 42279
rect 36921 42245 36955 42279
rect 40141 42245 40175 42279
rect 42717 42245 42751 42279
rect 7113 42177 7147 42211
rect 8953 42177 8987 42211
rect 11897 42177 11931 42211
rect 12357 42177 12391 42211
rect 14933 42177 14967 42211
rect 15026 42177 15060 42211
rect 15209 42177 15243 42211
rect 15439 42177 15473 42211
rect 15669 42177 15703 42211
rect 15853 42177 15887 42211
rect 18337 42177 18371 42211
rect 18485 42177 18519 42211
rect 18613 42177 18647 42211
rect 18705 42177 18739 42211
rect 18802 42177 18836 42211
rect 19073 42177 19107 42211
rect 21833 42177 21867 42211
rect 26985 42177 27019 42211
rect 27353 42177 27387 42211
rect 33977 42177 34011 42211
rect 34621 42177 34655 42211
rect 35265 42177 35299 42211
rect 38853 42177 38887 42211
rect 39037 42177 39071 42211
rect 42073 42177 42107 42211
rect 7389 42109 7423 42143
rect 8861 42109 8895 42143
rect 11989 42109 12023 42143
rect 12173 42109 12207 42143
rect 12909 42109 12943 42143
rect 13093 42109 13127 42143
rect 13369 42109 13403 42143
rect 17325 42109 17359 42143
rect 19349 42109 19383 42143
rect 21465 42109 21499 42143
rect 22109 42109 22143 42143
rect 25053 42109 25087 42143
rect 34713 42109 34747 42143
rect 34989 42109 35023 42143
rect 35817 42109 35851 42143
rect 39865 42109 39899 42143
rect 42441 42109 42475 42143
rect 27537 42041 27571 42075
rect 11529 41973 11563 42007
rect 18981 41973 19015 42007
rect 20821 41973 20855 42007
rect 20913 41973 20947 42007
rect 23581 41973 23615 42007
rect 26801 41973 26835 42007
rect 32229 41973 32263 42007
rect 36461 41973 36495 42007
rect 36553 41973 36587 42007
rect 36737 41973 36771 42007
rect 41613 41973 41647 42007
rect 44189 41973 44223 42007
rect 7757 41769 7791 41803
rect 10149 41769 10183 41803
rect 11989 41769 12023 41803
rect 14105 41769 14139 41803
rect 17325 41769 17359 41803
rect 17969 41769 18003 41803
rect 19901 41769 19935 41803
rect 21465 41769 21499 41803
rect 31309 41769 31343 41803
rect 35173 41769 35207 41803
rect 36737 41769 36771 41803
rect 39313 41769 39347 41803
rect 41797 41769 41831 41803
rect 42073 41769 42107 41803
rect 42257 41769 42291 41803
rect 13645 41701 13679 41735
rect 8677 41633 8711 41667
rect 9597 41633 9631 41667
rect 10241 41633 10275 41667
rect 14657 41633 14691 41667
rect 19257 41633 19291 41667
rect 24961 41633 24995 41667
rect 40693 41633 40727 41667
rect 41153 41633 41187 41667
rect 42533 41633 42567 41667
rect 42809 41633 42843 41667
rect 7941 41565 7975 41599
rect 8401 41565 8435 41599
rect 12265 41565 12299 41599
rect 13001 41565 13035 41599
rect 13094 41565 13128 41599
rect 13466 41565 13500 41599
rect 16681 41565 16715 41599
rect 16774 41565 16808 41599
rect 17049 41565 17083 41599
rect 17146 41565 17180 41599
rect 17601 41565 17635 41599
rect 17785 41565 17819 41599
rect 20821 41565 20855 41599
rect 20914 41565 20948 41599
rect 21286 41565 21320 41599
rect 32689 41565 32723 41599
rect 33057 41565 33091 41599
rect 34483 41565 34517 41599
rect 35357 41565 35391 41599
rect 36093 41565 36127 41599
rect 36185 41565 36219 41599
rect 36369 41565 36403 41599
rect 38209 41565 38243 41599
rect 40233 41565 40267 41599
rect 40877 41565 40911 41599
rect 40969 41565 41003 41599
rect 41061 41565 41095 41599
rect 10517 41497 10551 41531
rect 12909 41497 12943 41531
rect 13277 41497 13311 41531
rect 13369 41497 13403 41531
rect 16957 41497 16991 41531
rect 21097 41497 21131 41531
rect 21189 41497 21223 41531
rect 24409 41497 24443 41531
rect 32597 41497 32631 41531
rect 39497 41497 39531 41531
rect 40325 41497 40359 41531
rect 40417 41497 40451 41531
rect 40601 41497 40635 41531
rect 41429 41497 41463 41531
rect 41613 41497 41647 41531
rect 41889 41497 41923 41531
rect 8033 41429 8067 41463
rect 8493 41429 8527 41463
rect 9689 41429 9723 41463
rect 9781 41429 9815 41463
rect 35449 41429 35483 41463
rect 36277 41429 36311 41463
rect 39129 41429 39163 41463
rect 39297 41429 39331 41463
rect 40049 41429 40083 41463
rect 42089 41429 42123 41463
rect 44281 41429 44315 41463
rect 10977 41225 11011 41259
rect 11897 41225 11931 41259
rect 33977 41225 34011 41259
rect 34805 41225 34839 41259
rect 39037 41225 39071 41259
rect 39129 41225 39163 41259
rect 40509 41225 40543 41259
rect 42073 41225 42107 41259
rect 13369 41157 13403 41191
rect 13737 41157 13771 41191
rect 15669 41157 15703 41191
rect 16681 41157 16715 41191
rect 21925 41157 21959 41191
rect 22385 41157 22419 41191
rect 35081 41157 35115 41191
rect 35633 41157 35667 41191
rect 39497 41157 39531 41191
rect 44065 41157 44099 41191
rect 44281 41157 44315 41191
rect 9137 41089 9171 41123
rect 11161 41089 11195 41123
rect 16313 41089 16347 41123
rect 17325 41089 17359 41123
rect 18153 41089 18187 41123
rect 18337 41089 18371 41123
rect 19349 41089 19383 41123
rect 19533 41089 19567 41123
rect 19625 41089 19659 41123
rect 21833 41089 21867 41123
rect 22109 41089 22143 41123
rect 22293 41089 22327 41123
rect 23305 41089 23339 41123
rect 34069 41089 34103 41123
rect 37289 41089 37323 41123
rect 39313 41089 39347 41123
rect 40049 41089 40083 41123
rect 41981 41089 42015 41123
rect 42165 41089 42199 41123
rect 42625 41089 42659 41123
rect 43085 41089 43119 41123
rect 13645 41021 13679 41055
rect 14289 41021 14323 41055
rect 15485 41021 15519 41055
rect 15577 41021 15611 41055
rect 17969 41021 18003 41055
rect 20453 41021 20487 41055
rect 22937 41021 22971 41055
rect 35357 41021 35391 41055
rect 37105 41021 37139 41055
rect 37565 41021 37599 41055
rect 42809 41021 42843 41055
rect 43821 41021 43855 41055
rect 16037 40953 16071 40987
rect 40417 40953 40451 40987
rect 10425 40885 10459 40919
rect 16129 40885 16163 40919
rect 19165 40885 19199 40919
rect 19901 40885 19935 40919
rect 23949 40885 23983 40919
rect 42441 40885 42475 40919
rect 42809 40885 42843 40919
rect 43177 40885 43211 40919
rect 43913 40885 43947 40919
rect 44097 40885 44131 40919
rect 12909 40681 12943 40715
rect 17049 40681 17083 40715
rect 18245 40681 18279 40715
rect 20624 40681 20658 40715
rect 22201 40681 22235 40715
rect 35265 40681 35299 40715
rect 36737 40681 36771 40715
rect 38025 40681 38059 40715
rect 40601 40681 40635 40715
rect 43361 40681 43395 40715
rect 35817 40613 35851 40647
rect 42993 40613 43027 40647
rect 10885 40545 10919 40579
rect 11713 40545 11747 40579
rect 13001 40545 13035 40579
rect 15577 40545 15611 40579
rect 19809 40545 19843 40579
rect 20361 40545 20395 40579
rect 23673 40545 23707 40579
rect 23949 40545 23983 40579
rect 35725 40545 35759 40579
rect 40141 40545 40175 40579
rect 8217 40477 8251 40511
rect 9137 40477 9171 40511
rect 12265 40477 12299 40511
rect 12413 40477 12447 40511
rect 12771 40477 12805 40511
rect 13553 40477 13587 40511
rect 15301 40477 15335 40511
rect 17693 40477 17727 40511
rect 18061 40477 18095 40511
rect 18797 40477 18831 40511
rect 24409 40477 24443 40511
rect 34713 40477 34747 40511
rect 34897 40477 34931 40511
rect 34989 40477 35023 40511
rect 35081 40477 35115 40511
rect 35541 40477 35575 40511
rect 36369 40477 36403 40511
rect 36737 40477 36771 40511
rect 36829 40477 36863 40511
rect 38209 40477 38243 40511
rect 40233 40477 40267 40511
rect 40601 40477 40635 40511
rect 42717 40477 42751 40511
rect 42993 40477 43027 40511
rect 43177 40477 43211 40511
rect 43361 40477 43395 40511
rect 43453 40477 43487 40511
rect 44005 40477 44039 40511
rect 9413 40409 9447 40443
rect 12541 40409 12575 40443
rect 12633 40409 12667 40443
rect 17141 40409 17175 40443
rect 35265 40409 35299 40443
rect 36553 40409 36587 40443
rect 42809 40409 42843 40443
rect 8769 40341 8803 40375
rect 11161 40341 11195 40375
rect 17877 40341 17911 40375
rect 19257 40341 19291 40375
rect 22109 40341 22143 40375
rect 25053 40341 25087 40375
rect 34805 40341 34839 40375
rect 35357 40341 35391 40375
rect 37013 40341 37047 40375
rect 40785 40341 40819 40375
rect 8585 40137 8619 40171
rect 9045 40137 9079 40171
rect 10241 40137 10275 40171
rect 11345 40137 11379 40171
rect 21097 40137 21131 40171
rect 21833 40137 21867 40171
rect 22293 40137 22327 40171
rect 24133 40137 24167 40171
rect 36001 40137 36035 40171
rect 13921 40069 13955 40103
rect 16129 40069 16163 40103
rect 16957 40069 16991 40103
rect 18797 40069 18831 40103
rect 23765 40069 23799 40103
rect 23857 40069 23891 40103
rect 9689 40001 9723 40035
rect 9781 40001 9815 40035
rect 9965 40001 9999 40035
rect 10977 40001 11011 40035
rect 11161 40001 11195 40035
rect 18521 40001 18555 40035
rect 21281 40001 21315 40035
rect 22201 40001 22235 40035
rect 23489 40001 23523 40035
rect 23609 40001 23643 40035
rect 23954 40001 23988 40035
rect 25881 40001 25915 40035
rect 27169 40001 27203 40035
rect 40601 40001 40635 40035
rect 41245 40001 41279 40035
rect 41429 40001 41463 40035
rect 43361 40001 43395 40035
rect 43453 40001 43487 40035
rect 43637 40001 43671 40035
rect 6837 39933 6871 39967
rect 7113 39933 7147 39967
rect 9137 39933 9171 39967
rect 9321 39933 9355 39967
rect 10149 39933 10183 39967
rect 10793 39933 10827 39967
rect 12541 39933 12575 39967
rect 12817 39933 12851 39967
rect 16221 39933 16255 39967
rect 16313 39933 16347 39967
rect 16681 39933 16715 39967
rect 20269 39933 20303 39967
rect 22477 39933 22511 39967
rect 24593 39933 24627 39967
rect 32413 39933 32447 39967
rect 34253 39933 34287 39967
rect 34529 39933 34563 39967
rect 38485 39933 38519 39967
rect 38761 39933 38795 39967
rect 40233 39933 40267 39967
rect 42717 39933 42751 39967
rect 18429 39865 18463 39899
rect 8677 39797 8711 39831
rect 11989 39797 12023 39831
rect 13369 39797 13403 39831
rect 15209 39797 15243 39831
rect 15761 39797 15795 39831
rect 25237 39797 25271 39831
rect 25329 39797 25363 39831
rect 26985 39797 27019 39831
rect 33057 39797 33091 39831
rect 41153 39797 41187 39831
rect 41245 39797 41279 39831
rect 43637 39797 43671 39831
rect 7389 39593 7423 39627
rect 13277 39593 13311 39627
rect 17049 39593 17083 39627
rect 26157 39593 26191 39627
rect 35081 39593 35115 39627
rect 39405 39593 39439 39627
rect 40049 39593 40083 39627
rect 40233 39593 40267 39627
rect 42441 39593 42475 39627
rect 16037 39525 16071 39559
rect 17509 39525 17543 39559
rect 9597 39457 9631 39491
rect 11529 39457 11563 39491
rect 11805 39457 11839 39491
rect 16405 39457 16439 39491
rect 17141 39457 17175 39491
rect 18245 39457 18279 39491
rect 19257 39457 19291 39491
rect 24409 39457 24443 39491
rect 26433 39457 26467 39491
rect 26709 39457 26743 39491
rect 28181 39457 28215 39491
rect 31769 39457 31803 39491
rect 32045 39457 32079 39491
rect 32137 39457 32171 39491
rect 32413 39457 32447 39491
rect 40601 39457 40635 39491
rect 44189 39457 44223 39491
rect 7573 39389 7607 39423
rect 13737 39389 13771 39423
rect 14289 39389 14323 39423
rect 17325 39389 17359 39423
rect 18889 39389 18923 39423
rect 22293 39389 22327 39423
rect 22569 39389 22603 39423
rect 29009 39389 29043 39423
rect 35081 39389 35115 39423
rect 35265 39389 35299 39423
rect 38025 39389 38059 39423
rect 38209 39389 38243 39423
rect 39221 39389 39255 39423
rect 39405 39389 39439 39423
rect 40509 39389 40543 39423
rect 40693 39389 40727 39423
rect 42165 39389 42199 39423
rect 42349 39389 42383 39423
rect 9873 39321 9907 39355
rect 14565 39321 14599 39355
rect 16681 39321 16715 39355
rect 17601 39321 17635 39355
rect 19533 39321 19567 39355
rect 24685 39321 24719 39355
rect 28825 39321 28859 39355
rect 40417 39321 40451 39355
rect 42257 39321 42291 39355
rect 43913 39321 43947 39355
rect 11345 39253 11379 39287
rect 13921 39253 13955 39287
rect 16589 39253 16623 39287
rect 19073 39253 19107 39287
rect 21005 39253 21039 39287
rect 22109 39253 22143 39287
rect 22477 39253 22511 39287
rect 28641 39253 28675 39287
rect 30297 39253 30331 39287
rect 33885 39253 33919 39287
rect 38117 39253 38151 39287
rect 40212 39253 40246 39287
rect 7665 39049 7699 39083
rect 9597 39049 9631 39083
rect 10057 39049 10091 39083
rect 10517 39049 10551 39083
rect 10977 39049 11011 39083
rect 12081 39049 12115 39083
rect 12817 39049 12851 39083
rect 15485 39049 15519 39083
rect 19533 39049 19567 39083
rect 19993 39049 20027 39083
rect 24409 39049 24443 39083
rect 32137 39049 32171 39083
rect 44005 39049 44039 39083
rect 12449 38981 12483 39015
rect 18153 38981 18187 39015
rect 24133 38981 24167 39015
rect 26709 38981 26743 39015
rect 32643 38981 32677 39015
rect 33149 38981 33183 39015
rect 33254 38981 33288 39015
rect 36737 38981 36771 39015
rect 42533 38981 42567 39015
rect 7297 38913 7331 38947
rect 8033 38913 8067 38947
rect 8493 38913 8527 38947
rect 9321 38913 9355 38947
rect 10241 38913 10275 38947
rect 10885 38913 10919 38947
rect 12260 38913 12294 38947
rect 12357 38913 12391 38947
rect 12632 38913 12666 38947
rect 12725 38913 12759 38947
rect 14565 38913 14599 38947
rect 15761 38913 15795 38947
rect 17969 38913 18003 38947
rect 19901 38913 19935 38947
rect 20453 38913 20487 38947
rect 23765 38913 23799 38947
rect 23913 38913 23947 38947
rect 24041 38913 24075 38947
rect 24230 38913 24264 38947
rect 24501 38913 24535 38947
rect 26341 38913 26375 38947
rect 27353 38913 27387 38947
rect 27997 38913 28031 38947
rect 32321 38913 32355 38947
rect 32413 38913 32447 38947
rect 32505 38913 32539 38947
rect 33057 38913 33091 38947
rect 33359 38913 33393 38947
rect 34253 38913 34287 38947
rect 40325 38913 40359 38947
rect 40601 38913 40635 38947
rect 40785 38913 40819 38947
rect 8125 38845 8159 38879
rect 8309 38845 8343 38879
rect 9045 38845 9079 38879
rect 11161 38845 11195 38879
rect 14289 38845 14323 38879
rect 14657 38845 14691 38879
rect 15209 38845 15243 38879
rect 17785 38845 17819 38879
rect 20177 38845 20211 38879
rect 22017 38845 22051 38879
rect 23029 38845 23063 38879
rect 23581 38845 23615 38879
rect 24777 38845 24811 38879
rect 27445 38845 27479 38879
rect 27629 38845 27663 38879
rect 28273 38845 28307 38879
rect 29745 38845 29779 38879
rect 30389 38845 30423 38879
rect 32781 38845 32815 38879
rect 33517 38845 33551 38879
rect 33701 38845 33735 38879
rect 36553 38845 36587 38879
rect 38761 38845 38795 38879
rect 39037 38845 39071 38879
rect 40141 38845 40175 38879
rect 29837 38777 29871 38811
rect 32873 38777 32907 38811
rect 37013 38777 37047 38811
rect 40601 38777 40635 38811
rect 7113 38709 7147 38743
rect 20545 38709 20579 38743
rect 22661 38709 22695 38743
rect 26249 38709 26283 38743
rect 26985 38709 27019 38743
rect 35909 38709 35943 38743
rect 37289 38709 37323 38743
rect 40509 38709 40543 38743
rect 13645 38505 13679 38539
rect 23581 38505 23615 38539
rect 28365 38505 28399 38539
rect 32689 38505 32723 38539
rect 33241 38505 33275 38539
rect 33701 38505 33735 38539
rect 41613 38505 41647 38539
rect 9321 38437 9355 38471
rect 6469 38369 6503 38403
rect 8217 38369 8251 38403
rect 8953 38369 8987 38403
rect 9413 38369 9447 38403
rect 10517 38369 10551 38403
rect 15485 38369 15519 38403
rect 16497 38369 16531 38403
rect 18245 38369 18279 38403
rect 19993 38369 20027 38403
rect 21833 38369 21867 38403
rect 22109 38369 22143 38403
rect 25421 38369 25455 38403
rect 29009 38369 29043 38403
rect 29653 38369 29687 38403
rect 31401 38369 31435 38403
rect 32045 38369 32079 38403
rect 38025 38369 38059 38403
rect 42717 38369 42751 38403
rect 43453 38369 43487 38403
rect 9137 38301 9171 38335
rect 9597 38301 9631 38335
rect 9873 38301 9907 38335
rect 11437 38301 11471 38335
rect 13001 38301 13035 38335
rect 13149 38301 13183 38335
rect 13277 38301 13311 38335
rect 13369 38301 13403 38335
rect 13507 38301 13541 38335
rect 18889 38301 18923 38335
rect 28549 38301 28583 38335
rect 29101 38301 29135 38335
rect 29285 38301 29319 38335
rect 32873 38301 32907 38335
rect 33149 38301 33183 38335
rect 33241 38301 33275 38335
rect 33333 38301 33367 38335
rect 33609 38301 33643 38335
rect 33793 38301 33827 38335
rect 34989 38301 35023 38335
rect 37749 38301 37783 38335
rect 37933 38301 37967 38335
rect 39865 38301 39899 38335
rect 42625 38301 42659 38335
rect 43269 38301 43303 38335
rect 6745 38233 6779 38267
rect 9781 38233 9815 38267
rect 10885 38233 10919 38267
rect 17969 38233 18003 38267
rect 20269 38233 20303 38267
rect 27169 38233 27203 38267
rect 28641 38233 28675 38267
rect 28733 38233 28767 38267
rect 28871 38233 28905 38267
rect 29929 38233 29963 38267
rect 33517 38233 33551 38267
rect 35265 38233 35299 38267
rect 37841 38233 37875 38267
rect 40141 38233 40175 38267
rect 43085 38233 43119 38267
rect 9965 38165 9999 38199
rect 14841 38165 14875 38199
rect 18337 38165 18371 38199
rect 21741 38165 21775 38199
rect 29193 38165 29227 38199
rect 31493 38165 31527 38199
rect 33057 38165 33091 38199
rect 36737 38165 36771 38199
rect 38669 38165 38703 38199
rect 42993 38165 43027 38199
rect 11161 37961 11195 37995
rect 18521 37961 18555 37995
rect 21189 37961 21223 37995
rect 21833 37961 21867 37995
rect 22201 37961 22235 37995
rect 25237 37961 25271 37995
rect 30573 37961 30607 37995
rect 33149 37961 33183 37995
rect 35633 37961 35667 37995
rect 38025 37961 38059 37995
rect 38853 37961 38887 37995
rect 40233 37961 40267 37995
rect 42625 37961 42659 37995
rect 9689 37893 9723 37927
rect 22293 37893 22327 37927
rect 29161 37893 29195 37927
rect 29377 37893 29411 37927
rect 31059 37893 31093 37927
rect 36061 37893 36095 37927
rect 36277 37893 36311 37927
rect 38269 37893 38303 37927
rect 38485 37893 38519 37927
rect 6561 37825 6595 37859
rect 9413 37825 9447 37859
rect 13185 37825 13219 37859
rect 13369 37825 13403 37859
rect 13461 37825 13495 37859
rect 17049 37825 17083 37859
rect 17197 37825 17231 37859
rect 17325 37825 17359 37859
rect 17417 37825 17451 37859
rect 17553 37825 17587 37859
rect 20361 37825 20395 37859
rect 21373 37825 21407 37859
rect 24777 37825 24811 37859
rect 25329 37825 25363 37859
rect 27169 37825 27203 37859
rect 27261 37825 27295 37859
rect 27353 37825 27387 37859
rect 27471 37825 27505 37859
rect 28641 37825 28675 37859
rect 28825 37825 28859 37859
rect 28917 37825 28951 37859
rect 30757 37825 30791 37859
rect 30849 37825 30883 37859
rect 30941 37825 30975 37859
rect 31217 37825 31251 37859
rect 33333 37825 33367 37859
rect 33517 37825 33551 37859
rect 34989 37825 35023 37859
rect 35541 37825 35575 37859
rect 35817 37825 35851 37859
rect 36369 37825 36403 37859
rect 37013 37825 37047 37859
rect 37473 37825 37507 37859
rect 37841 37825 37875 37859
rect 38577 37825 38611 37859
rect 40233 37825 40267 37859
rect 43545 37825 43579 37859
rect 6837 37757 6871 37791
rect 8309 37757 8343 37791
rect 8953 37757 8987 37791
rect 14289 37757 14323 37791
rect 14565 37757 14599 37791
rect 17877 37757 17911 37791
rect 20085 37757 20119 37791
rect 20453 37757 20487 37791
rect 21005 37757 21039 37791
rect 22385 37757 22419 37791
rect 27629 37757 27663 37791
rect 27721 37757 27755 37791
rect 28273 37757 28307 37791
rect 35081 37757 35115 37791
rect 35357 37757 35391 37791
rect 37381 37757 37415 37791
rect 38853 37757 38887 37791
rect 39957 37757 39991 37791
rect 40141 37757 40175 37791
rect 43177 37757 43211 37791
rect 17693 37689 17727 37723
rect 24593 37689 24627 37723
rect 28457 37689 28491 37723
rect 8401 37621 8435 37655
rect 13001 37621 13035 37655
rect 16037 37621 16071 37655
rect 18613 37621 18647 37655
rect 26985 37621 27019 37655
rect 29009 37621 29043 37655
rect 29193 37621 29227 37655
rect 35817 37621 35851 37655
rect 35909 37621 35943 37655
rect 36093 37621 36127 37655
rect 37841 37621 37875 37655
rect 38117 37621 38151 37655
rect 38301 37621 38335 37655
rect 38669 37621 38703 37655
rect 44189 37621 44223 37655
rect 7113 37417 7147 37451
rect 16681 37417 16715 37451
rect 20729 37417 20763 37451
rect 25237 37417 25271 37451
rect 27813 37417 27847 37451
rect 36829 37417 36863 37451
rect 40509 37417 40543 37451
rect 42257 37417 42291 37451
rect 41061 37349 41095 37383
rect 8217 37281 8251 37315
rect 8953 37281 8987 37315
rect 11161 37281 11195 37315
rect 11345 37281 11379 37315
rect 12633 37281 12667 37315
rect 14657 37281 14691 37315
rect 16037 37281 16071 37315
rect 16313 37281 16347 37315
rect 26065 37281 26099 37315
rect 26341 37281 26375 37315
rect 35081 37281 35115 37315
rect 37841 37281 37875 37315
rect 44005 37281 44039 37315
rect 1409 37213 1443 37247
rect 7297 37213 7331 37247
rect 8033 37213 8067 37247
rect 9137 37213 9171 37247
rect 13277 37213 13311 37247
rect 13921 37213 13955 37247
rect 16497 37213 16531 37247
rect 17049 37213 17083 37247
rect 19257 37213 19291 37247
rect 22477 37213 22511 37247
rect 23857 37213 23891 37247
rect 24409 37213 24443 37247
rect 25513 37213 25547 37247
rect 25697 37213 25731 37247
rect 25881 37213 25915 37247
rect 33241 37213 33275 37247
rect 38025 37213 38059 37247
rect 38209 37213 38243 37247
rect 40141 37213 40175 37247
rect 40509 37213 40543 37247
rect 40785 37213 40819 37247
rect 40969 37213 41003 37247
rect 44281 37213 44315 37247
rect 9321 37145 9355 37179
rect 14841 37145 14875 37179
rect 15485 37145 15519 37179
rect 17325 37145 17359 37179
rect 23121 37145 23155 37179
rect 25789 37145 25823 37179
rect 33425 37145 33459 37179
rect 35357 37145 35391 37179
rect 41337 37145 41371 37179
rect 42073 37145 42107 37179
rect 42289 37145 42323 37179
rect 1593 37077 1627 37111
rect 7665 37077 7699 37111
rect 8125 37077 8159 37111
rect 10701 37077 10735 37111
rect 11069 37077 11103 37111
rect 13185 37077 13219 37111
rect 14749 37077 14783 37111
rect 15209 37077 15243 37111
rect 18797 37077 18831 37111
rect 23213 37077 23247 37111
rect 25053 37077 25087 37111
rect 33057 37077 33091 37111
rect 41245 37077 41279 37111
rect 41429 37077 41463 37111
rect 41613 37077 41647 37111
rect 42441 37077 42475 37111
rect 42533 37077 42567 37111
rect 12265 36873 12299 36907
rect 15301 36873 15335 36907
rect 17325 36873 17359 36907
rect 19441 36873 19475 36907
rect 23857 36873 23891 36907
rect 28365 36873 28399 36907
rect 32229 36873 32263 36907
rect 33057 36873 33091 36907
rect 33885 36873 33919 36907
rect 34069 36873 34103 36907
rect 35909 36873 35943 36907
rect 41889 36873 41923 36907
rect 13737 36805 13771 36839
rect 16037 36805 16071 36839
rect 19165 36805 19199 36839
rect 22661 36805 22695 36839
rect 25329 36805 25363 36839
rect 33701 36805 33735 36839
rect 35633 36805 35667 36839
rect 38117 36805 38151 36839
rect 40693 36805 40727 36839
rect 4353 36737 4387 36771
rect 6929 36737 6963 36771
rect 14013 36737 14047 36771
rect 15485 36737 15519 36771
rect 16405 36737 16439 36771
rect 16773 36737 16807 36771
rect 16865 36737 16899 36771
rect 17049 36737 17083 36771
rect 18705 36737 18739 36771
rect 18797 36737 18831 36771
rect 18945 36737 18979 36771
rect 19073 36737 19107 36771
rect 19262 36737 19296 36771
rect 19901 36737 19935 36771
rect 20453 36737 20487 36771
rect 21373 36737 21407 36771
rect 22569 36737 22603 36771
rect 25605 36737 25639 36771
rect 25973 36737 26007 36771
rect 27169 36737 27203 36771
rect 27905 36737 27939 36771
rect 28181 36737 28215 36771
rect 28457 36737 28491 36771
rect 30297 36737 30331 36771
rect 32413 36737 32447 36771
rect 32873 36737 32907 36771
rect 32965 36737 32999 36771
rect 33333 36737 33367 36771
rect 33517 36737 33551 36771
rect 33793 36737 33827 36771
rect 33977 36737 34011 36771
rect 34069 36737 34103 36771
rect 34253 36737 34287 36771
rect 35909 36737 35943 36771
rect 37749 36737 37783 36771
rect 37933 36737 37967 36771
rect 38025 36737 38059 36771
rect 38209 36737 38243 36771
rect 38577 36737 38611 36771
rect 41613 36737 41647 36771
rect 42073 36737 42107 36771
rect 42257 36737 42291 36771
rect 42441 36737 42475 36771
rect 1777 36669 1811 36703
rect 4629 36669 4663 36703
rect 6101 36669 6135 36703
rect 8677 36669 8711 36703
rect 9597 36669 9631 36703
rect 9873 36669 9907 36703
rect 17233 36669 17267 36703
rect 17877 36669 17911 36703
rect 19625 36669 19659 36703
rect 19809 36669 19843 36703
rect 21005 36669 21039 36703
rect 22753 36669 22787 36703
rect 23673 36669 23707 36703
rect 27813 36669 27847 36703
rect 28089 36669 28123 36703
rect 32505 36669 32539 36703
rect 32597 36669 32631 36703
rect 32689 36669 32723 36703
rect 33241 36669 33275 36703
rect 39129 36669 39163 36703
rect 42717 36669 42751 36703
rect 2145 36601 2179 36635
rect 18061 36601 18095 36635
rect 20269 36601 20303 36635
rect 26249 36601 26283 36635
rect 33149 36601 33183 36635
rect 35817 36601 35851 36635
rect 40417 36601 40451 36635
rect 41797 36601 41831 36635
rect 2237 36533 2271 36567
rect 11345 36533 11379 36567
rect 21189 36533 21223 36567
rect 22201 36533 22235 36567
rect 23121 36533 23155 36567
rect 26985 36533 27019 36567
rect 27537 36533 27571 36567
rect 27721 36533 27755 36567
rect 30113 36533 30147 36567
rect 37749 36533 37783 36567
rect 44189 36533 44223 36567
rect 5917 36329 5951 36363
rect 20747 36329 20781 36363
rect 21741 36329 21775 36363
rect 23581 36329 23615 36363
rect 24409 36329 24443 36363
rect 27997 36329 28031 36363
rect 32413 36329 32447 36363
rect 33241 36329 33275 36363
rect 33885 36329 33919 36363
rect 38853 36329 38887 36363
rect 42441 36329 42475 36363
rect 43085 36329 43119 36363
rect 8677 36261 8711 36295
rect 10333 36261 10367 36295
rect 16681 36261 16715 36295
rect 21649 36261 21683 36295
rect 25329 36261 25363 36295
rect 31769 36261 31803 36295
rect 33793 36261 33827 36295
rect 3801 36193 3835 36227
rect 6929 36193 6963 36227
rect 11805 36193 11839 36227
rect 14933 36193 14967 36227
rect 17417 36193 17451 36227
rect 21005 36193 21039 36227
rect 23213 36193 23247 36227
rect 23489 36193 23523 36227
rect 26249 36193 26283 36227
rect 26525 36193 26559 36227
rect 31401 36193 31435 36227
rect 32505 36193 32539 36227
rect 37381 36193 37415 36227
rect 40141 36193 40175 36227
rect 42625 36193 42659 36227
rect 6101 36125 6135 36159
rect 10517 36125 10551 36159
rect 14657 36125 14691 36159
rect 21465 36125 21499 36159
rect 23765 36125 23799 36159
rect 23949 36125 23983 36159
rect 24041 36125 24075 36159
rect 24588 36125 24622 36159
rect 24960 36125 24994 36159
rect 25053 36125 25087 36159
rect 25605 36125 25639 36159
rect 28273 36125 28307 36159
rect 28549 36125 28583 36159
rect 29837 36125 29871 36159
rect 29929 36125 29963 36159
rect 30297 36125 30331 36159
rect 30389 36125 30423 36159
rect 30941 36125 30975 36159
rect 31493 36125 31527 36159
rect 31953 36125 31987 36159
rect 32229 36125 32263 36159
rect 32597 36125 32631 36159
rect 33149 36125 33183 36159
rect 33333 36125 33367 36159
rect 33425 36125 33459 36159
rect 34253 36125 34287 36159
rect 37105 36125 37139 36159
rect 39865 36125 39899 36159
rect 39957 36125 39991 36159
rect 42717 36125 42751 36159
rect 42809 36125 42843 36159
rect 42993 36125 43027 36159
rect 43177 36125 43211 36159
rect 4077 36057 4111 36091
rect 7205 36057 7239 36091
rect 12081 36057 12115 36091
rect 15209 36057 15243 36091
rect 24685 36057 24719 36091
rect 24777 36057 24811 36091
rect 30021 36057 30055 36091
rect 30139 36057 30173 36091
rect 32321 36057 32355 36091
rect 33609 36057 33643 36091
rect 34069 36057 34103 36091
rect 5549 35989 5583 36023
rect 13553 35989 13587 36023
rect 14105 35989 14139 36023
rect 16773 35989 16807 36023
rect 19257 35989 19291 36023
rect 28089 35989 28123 36023
rect 28457 35989 28491 36023
rect 29653 35989 29687 36023
rect 31125 35989 31159 36023
rect 32137 35989 32171 36023
rect 32781 35989 32815 36023
rect 39865 35989 39899 36023
rect 2881 35785 2915 35819
rect 5825 35785 5859 35819
rect 7481 35785 7515 35819
rect 12541 35785 12575 35819
rect 13461 35785 13495 35819
rect 14841 35785 14875 35819
rect 15393 35785 15427 35819
rect 17325 35785 17359 35819
rect 25513 35785 25547 35819
rect 27169 35785 27203 35819
rect 27337 35785 27371 35819
rect 30389 35785 30423 35819
rect 30665 35785 30699 35819
rect 31401 35785 31435 35819
rect 5457 35717 5491 35751
rect 5657 35717 5691 35751
rect 13553 35717 13587 35751
rect 15485 35717 15519 35751
rect 26341 35717 26375 35751
rect 27537 35717 27571 35751
rect 28917 35717 28951 35751
rect 30941 35717 30975 35751
rect 32597 35717 32631 35751
rect 33241 35717 33275 35751
rect 39681 35717 39715 35751
rect 2697 35649 2731 35683
rect 7665 35649 7699 35683
rect 12081 35649 12115 35683
rect 12725 35649 12759 35683
rect 14657 35649 14691 35683
rect 17141 35649 17175 35683
rect 20453 35649 20487 35683
rect 23581 35649 23615 35683
rect 27813 35649 27847 35683
rect 27997 35649 28031 35683
rect 28457 35649 28491 35683
rect 30665 35649 30699 35683
rect 30757 35649 30791 35683
rect 31309 35649 31343 35683
rect 31493 35649 31527 35683
rect 31585 35649 31619 35683
rect 31769 35649 31803 35683
rect 32137 35649 32171 35683
rect 32302 35649 32336 35683
rect 32689 35649 32723 35683
rect 33425 35649 33459 35683
rect 33517 35649 33551 35683
rect 13737 35581 13771 35615
rect 15577 35581 15611 35615
rect 18613 35581 18647 35615
rect 23305 35581 23339 35615
rect 26065 35581 26099 35615
rect 27905 35581 27939 35615
rect 28089 35581 28123 35615
rect 28365 35581 28399 35615
rect 28641 35581 28675 35615
rect 36093 35581 36127 35615
rect 36369 35581 36403 35615
rect 39405 35581 39439 35615
rect 41153 35581 41187 35615
rect 41797 35581 41831 35615
rect 13093 35513 13127 35547
rect 15025 35513 15059 35547
rect 21833 35513 21867 35547
rect 32505 35513 32539 35547
rect 5641 35445 5675 35479
rect 12173 35445 12207 35479
rect 19165 35445 19199 35479
rect 20361 35445 20395 35479
rect 26617 35445 26651 35479
rect 27353 35445 27387 35479
rect 27629 35445 27663 35479
rect 31953 35445 31987 35479
rect 32413 35445 32447 35479
rect 34621 35445 34655 35479
rect 41245 35445 41279 35479
rect 7665 35241 7699 35275
rect 7849 35241 7883 35275
rect 8125 35241 8159 35275
rect 16957 35241 16991 35275
rect 18797 35241 18831 35275
rect 26065 35241 26099 35275
rect 39681 35241 39715 35275
rect 40049 35241 40083 35275
rect 41153 35241 41187 35275
rect 7481 35173 7515 35207
rect 11437 35173 11471 35207
rect 39865 35173 39899 35207
rect 40417 35173 40451 35207
rect 5733 35105 5767 35139
rect 17049 35105 17083 35139
rect 19257 35105 19291 35139
rect 26433 35105 26467 35139
rect 34989 35105 35023 35139
rect 35909 35105 35943 35139
rect 38761 35105 38795 35139
rect 39221 35105 39255 35139
rect 40969 35105 41003 35139
rect 42717 35105 42751 35139
rect 5253 35037 5287 35071
rect 5365 35037 5399 35071
rect 5457 35037 5491 35071
rect 5641 35037 5675 35071
rect 8493 35037 8527 35071
rect 8585 35037 8619 35071
rect 8769 35037 8803 35071
rect 8953 35037 8987 35071
rect 9137 35037 9171 35071
rect 9229 35037 9263 35071
rect 9321 35037 9355 35071
rect 9689 35037 9723 35071
rect 14565 35037 14599 35071
rect 16313 35037 16347 35071
rect 16589 35037 16623 35071
rect 16773 35037 16807 35071
rect 18889 35037 18923 35071
rect 22569 35037 22603 35071
rect 23489 35037 23523 35071
rect 25053 35037 25087 35071
rect 26249 35037 26283 35071
rect 31769 35037 31803 35071
rect 31953 35037 31987 35071
rect 39129 35037 39163 35071
rect 39405 35037 39439 35071
rect 39684 35037 39718 35071
rect 40877 35037 40911 35071
rect 43361 35037 43395 35071
rect 43545 35037 43579 35071
rect 4997 34969 5031 35003
rect 6009 34969 6043 35003
rect 8033 34969 8067 35003
rect 8309 34969 8343 35003
rect 9597 34969 9631 35003
rect 9965 34969 9999 35003
rect 17325 34969 17359 35003
rect 19533 34969 19567 35003
rect 23213 34969 23247 35003
rect 31861 34969 31895 35003
rect 36185 34969 36219 35003
rect 40233 34969 40267 35003
rect 40417 34969 40451 35003
rect 7833 34901 7867 34935
rect 8769 34901 8803 34935
rect 14473 34901 14507 34935
rect 15761 34901 15795 34935
rect 19073 34901 19107 34935
rect 21005 34901 21039 34935
rect 22845 34901 22879 34935
rect 24501 34901 24535 34935
rect 35633 34901 35667 34935
rect 37657 34901 37691 34935
rect 39497 34901 39531 34935
rect 40033 34901 40067 34935
rect 43269 34901 43303 34935
rect 43453 34901 43487 34935
rect 5641 34697 5675 34731
rect 6469 34697 6503 34731
rect 6745 34697 6779 34731
rect 8309 34697 8343 34731
rect 16221 34697 16255 34731
rect 17601 34697 17635 34731
rect 18889 34697 18923 34731
rect 19349 34697 19383 34731
rect 25973 34697 26007 34731
rect 35633 34697 35667 34731
rect 38025 34697 38059 34731
rect 40233 34697 40267 34731
rect 42257 34697 42291 34731
rect 42533 34697 42567 34731
rect 5825 34629 5859 34663
rect 17509 34629 17543 34663
rect 18705 34629 18739 34663
rect 23949 34629 23983 34663
rect 24501 34629 24535 34663
rect 27445 34629 27479 34663
rect 27813 34629 27847 34663
rect 35265 34629 35299 34663
rect 35357 34629 35391 34663
rect 36461 34629 36495 34663
rect 36661 34629 36695 34663
rect 41889 34629 41923 34663
rect 44005 34629 44039 34663
rect 42119 34595 42153 34629
rect 6009 34561 6043 34595
rect 6377 34561 6411 34595
rect 6561 34561 6595 34595
rect 6653 34561 6687 34595
rect 6837 34561 6871 34595
rect 7113 34561 7147 34595
rect 7205 34561 7239 34595
rect 8125 34561 8159 34595
rect 8309 34561 8343 34595
rect 8401 34561 8435 34595
rect 8585 34561 8619 34595
rect 8953 34561 8987 34595
rect 9045 34561 9079 34595
rect 11529 34561 11563 34595
rect 12449 34561 12483 34595
rect 12541 34561 12575 34595
rect 12725 34561 12759 34595
rect 13001 34561 13035 34595
rect 13185 34561 13219 34595
rect 14473 34561 14507 34595
rect 17233 34561 17267 34595
rect 17325 34561 17359 34595
rect 18521 34561 18555 34595
rect 18797 34561 18831 34595
rect 19257 34561 19291 34595
rect 23765 34561 23799 34595
rect 24041 34561 24075 34595
rect 27261 34561 27295 34595
rect 27537 34561 27571 34595
rect 27905 34561 27939 34595
rect 28181 34561 28215 34595
rect 28733 34561 28767 34595
rect 30757 34561 30791 34595
rect 30941 34561 30975 34595
rect 35081 34561 35115 34595
rect 35449 34561 35483 34595
rect 37473 34561 37507 34595
rect 37933 34561 37967 34595
rect 38393 34561 38427 34595
rect 40785 34561 40819 34595
rect 44281 34561 44315 34595
rect 8677 34493 8711 34527
rect 12909 34493 12943 34527
rect 14749 34493 14783 34527
rect 18245 34493 18279 34527
rect 18337 34493 18371 34527
rect 19441 34493 19475 34527
rect 22845 34493 22879 34527
rect 24225 34493 24259 34527
rect 30849 34493 30883 34527
rect 8585 34425 8619 34459
rect 8861 34425 8895 34459
rect 8769 34357 8803 34391
rect 9308 34357 9342 34391
rect 10793 34357 10827 34391
rect 11621 34357 11655 34391
rect 13001 34357 13035 34391
rect 23489 34357 23523 34391
rect 23581 34357 23615 34391
rect 27261 34357 27295 34391
rect 36645 34357 36679 34391
rect 36829 34357 36863 34391
rect 37657 34357 37691 34391
rect 39681 34357 39715 34391
rect 42073 34357 42107 34391
rect 6193 34153 6227 34187
rect 9229 34153 9263 34187
rect 12357 34153 12391 34187
rect 14289 34153 14323 34187
rect 14749 34153 14783 34187
rect 15945 34153 15979 34187
rect 17785 34153 17819 34187
rect 25053 34153 25087 34187
rect 28457 34153 28491 34187
rect 30389 34153 30423 34187
rect 31125 34153 31159 34187
rect 32873 34153 32907 34187
rect 34069 34153 34103 34187
rect 35173 34153 35207 34187
rect 39589 34153 39623 34187
rect 42993 34153 43027 34187
rect 13277 34085 13311 34119
rect 13369 34085 13403 34119
rect 13645 34085 13679 34119
rect 25145 34085 25179 34119
rect 10609 34017 10643 34051
rect 22569 34017 22603 34051
rect 22661 34017 22695 34051
rect 23949 34017 23983 34051
rect 25697 34017 25731 34051
rect 26985 34017 27019 34051
rect 33609 34017 33643 34051
rect 34161 34017 34195 34051
rect 34805 34017 34839 34051
rect 37473 34017 37507 34051
rect 37841 34017 37875 34051
rect 40969 34017 41003 34051
rect 41429 34017 41463 34051
rect 41889 34017 41923 34051
rect 5733 33949 5767 33983
rect 6101 33949 6135 33983
rect 6285 33949 6319 33983
rect 8953 33949 8987 33983
rect 9229 33949 9263 33983
rect 11437 33949 11471 33983
rect 11529 33949 11563 33983
rect 11621 33949 11655 33983
rect 11713 33949 11747 33983
rect 12081 33949 12115 33983
rect 12541 33949 12575 33983
rect 12633 33949 12667 33983
rect 13185 33949 13219 33983
rect 13461 33949 13495 33983
rect 13737 33949 13771 33983
rect 13921 33949 13955 33983
rect 14105 33949 14139 33983
rect 14289 33949 14323 33983
rect 14933 33949 14967 33983
rect 17417 33949 17451 33983
rect 20269 33949 20303 33983
rect 20453 33949 20487 33983
rect 24409 33949 24443 33983
rect 24557 33949 24591 33983
rect 24874 33949 24908 33983
rect 26709 33949 26743 33983
rect 30205 33949 30239 33983
rect 31033 33949 31067 33983
rect 31217 33949 31251 33983
rect 31401 33949 31435 33983
rect 32321 33949 32355 33983
rect 32505 33949 32539 33983
rect 32597 33949 32631 33983
rect 33701 33949 33735 33983
rect 34069 33949 34103 33983
rect 34897 33949 34931 33983
rect 40325 33949 40359 33983
rect 40509 33949 40543 33983
rect 40785 33949 40819 33983
rect 41521 33949 41555 33983
rect 42073 33949 42107 33983
rect 42717 33949 42751 33983
rect 42993 33949 43027 33983
rect 44281 33949 44315 33983
rect 11897 33881 11931 33915
rect 11989 33881 12023 33915
rect 12909 33881 12943 33915
rect 13001 33881 13035 33915
rect 17877 33881 17911 33915
rect 24685 33881 24719 33915
rect 24777 33881 24811 33915
rect 30021 33881 30055 33915
rect 30849 33881 30883 33915
rect 32781 33881 32815 33915
rect 38117 33881 38151 33915
rect 42625 33881 42659 33915
rect 42809 33881 42843 33915
rect 5641 33813 5675 33847
rect 9045 33813 9079 33847
rect 9965 33813 9999 33847
rect 12265 33813 12299 33847
rect 13829 33813 13863 33847
rect 20361 33813 20395 33847
rect 22753 33813 22787 33847
rect 23121 33813 23155 33847
rect 23397 33813 23431 33847
rect 30573 33813 30607 33847
rect 32045 33813 32079 33847
rect 32137 33813 32171 33847
rect 33333 33813 33367 33847
rect 34437 33813 34471 33847
rect 36921 33813 36955 33847
rect 40417 33813 40451 33847
rect 40601 33813 40635 33847
rect 44097 33813 44131 33847
rect 6377 33609 6411 33643
rect 12173 33609 12207 33643
rect 14841 33609 14875 33643
rect 15209 33609 15243 33643
rect 20269 33609 20303 33643
rect 22017 33609 22051 33643
rect 28733 33609 28767 33643
rect 31033 33609 31067 33643
rect 32305 33609 32339 33643
rect 33977 33609 34011 33643
rect 37289 33609 37323 33643
rect 41061 33609 41095 33643
rect 42441 33609 42475 33643
rect 14749 33541 14783 33575
rect 23489 33541 23523 33575
rect 26065 33541 26099 33575
rect 27261 33541 27295 33575
rect 31769 33541 31803 33575
rect 32505 33541 32539 33575
rect 33149 33541 33183 33575
rect 33609 33541 33643 33575
rect 36369 33541 36403 33575
rect 36461 33541 36495 33575
rect 43913 33541 43947 33575
rect 6009 33473 6043 33507
rect 6193 33473 6227 33507
rect 6561 33473 6595 33507
rect 9321 33473 9355 33507
rect 11805 33473 11839 33507
rect 11897 33473 11931 33507
rect 11989 33473 12023 33507
rect 12081 33473 12115 33507
rect 12357 33473 12391 33507
rect 12449 33473 12483 33507
rect 12725 33473 12759 33507
rect 16037 33473 16071 33507
rect 17049 33473 17083 33507
rect 17509 33473 17543 33507
rect 18429 33473 18463 33507
rect 18889 33473 18923 33507
rect 19257 33473 19291 33507
rect 19349 33473 19383 33507
rect 19717 33473 19751 33507
rect 20266 33473 20300 33507
rect 21097 33473 21131 33507
rect 21465 33473 21499 33507
rect 24041 33473 24075 33507
rect 26709 33473 26743 33507
rect 31401 33473 31435 33507
rect 32597 33473 32631 33507
rect 32781 33473 32815 33507
rect 33057 33473 33091 33507
rect 33241 33473 33275 33507
rect 33333 33473 33367 33507
rect 33426 33473 33460 33507
rect 33701 33473 33735 33507
rect 33798 33473 33832 33507
rect 34253 33473 34287 33507
rect 34529 33473 34563 33507
rect 34713 33473 34747 33507
rect 35173 33473 35207 33507
rect 36185 33473 36219 33507
rect 36553 33473 36587 33507
rect 3893 33405 3927 33439
rect 4169 33405 4203 33439
rect 5641 33405 5675 33439
rect 6745 33405 6779 33439
rect 12541 33405 12575 33439
rect 15301 33405 15335 33439
rect 15485 33405 15519 33439
rect 17141 33405 17175 33439
rect 17233 33405 17267 33439
rect 18061 33405 18095 33439
rect 18521 33405 18555 33439
rect 20729 33405 20763 33439
rect 21005 33405 21039 33439
rect 21373 33405 21407 33439
rect 23765 33405 23799 33439
rect 26341 33405 26375 33439
rect 26985 33405 27019 33439
rect 29285 33405 29319 33439
rect 29561 33405 29595 33439
rect 31309 33405 31343 33439
rect 31677 33405 31711 33439
rect 32689 33405 32723 33439
rect 35081 33405 35115 33439
rect 35541 33405 35575 33439
rect 38761 33405 38795 33439
rect 39037 33405 39071 33439
rect 39313 33405 39347 33439
rect 39589 33405 39623 33439
rect 44189 33405 44223 33439
rect 12357 33337 12391 33371
rect 13461 33337 13495 33371
rect 16681 33337 16715 33371
rect 20085 33337 20119 33371
rect 20821 33337 20855 33371
rect 24593 33337 24627 33371
rect 31125 33337 31159 33371
rect 32137 33337 32171 33371
rect 34069 33337 34103 33371
rect 36737 33337 36771 33371
rect 5825 33269 5859 33303
rect 9413 33269 9447 33303
rect 12541 33269 12575 33303
rect 12909 33269 12943 33303
rect 15853 33269 15887 33303
rect 18613 33269 18647 33303
rect 18797 33269 18831 33303
rect 19717 33269 19751 33303
rect 20637 33269 20671 33303
rect 23857 33269 23891 33303
rect 26525 33269 26559 33303
rect 32321 33269 32355 33303
rect 4629 33065 4663 33099
rect 5457 33065 5491 33099
rect 8677 33065 8711 33099
rect 13461 33065 13495 33099
rect 14105 33065 14139 33099
rect 17417 33065 17451 33099
rect 17969 33065 18003 33099
rect 19441 33065 19475 33099
rect 19901 33065 19935 33099
rect 21833 33065 21867 33099
rect 26525 33065 26559 33099
rect 28641 33065 28675 33099
rect 34897 33065 34931 33099
rect 35173 33065 35207 33099
rect 37933 33065 37967 33099
rect 40141 33065 40175 33099
rect 13829 32997 13863 33031
rect 21281 32997 21315 33031
rect 25053 32997 25087 33031
rect 34345 32997 34379 33031
rect 40233 32997 40267 33031
rect 43729 32997 43763 33031
rect 6929 32929 6963 32963
rect 13277 32929 13311 32963
rect 14657 32929 14691 32963
rect 15669 32929 15703 32963
rect 17601 32929 17635 32963
rect 19717 32929 19751 32963
rect 23305 32929 23339 32963
rect 25881 32929 25915 32963
rect 26893 32929 26927 32963
rect 34805 32929 34839 32963
rect 34989 32929 35023 32963
rect 43361 32929 43395 32963
rect 4813 32861 4847 32895
rect 13185 32861 13219 32895
rect 13461 32861 13495 32895
rect 13921 32861 13955 32895
rect 14289 32861 14323 32895
rect 14381 32861 14415 32895
rect 17785 32861 17819 32895
rect 19993 32861 20027 32895
rect 20269 32861 20303 32895
rect 20545 32861 20579 32895
rect 20729 32861 20763 32895
rect 21005 32861 21039 32895
rect 21281 32861 21315 32895
rect 23581 32861 23615 32895
rect 24409 32861 24443 32895
rect 24557 32861 24591 32895
rect 24777 32861 24811 32895
rect 24874 32861 24908 32895
rect 25789 32861 25823 32895
rect 26617 32861 26651 32895
rect 27169 32861 27203 32895
rect 31125 32861 31159 32895
rect 31401 32861 31435 32895
rect 31585 32861 31619 32895
rect 33701 32861 33735 32895
rect 33885 32861 33919 32895
rect 34161 32861 34195 32895
rect 34713 32861 34747 32895
rect 35081 32861 35115 32895
rect 35265 32861 35299 32895
rect 37657 32861 37691 32895
rect 40325 32861 40359 32895
rect 5441 32793 5475 32827
rect 5641 32793 5675 32827
rect 7205 32793 7239 32827
rect 14749 32793 14783 32827
rect 15945 32793 15979 32827
rect 20361 32793 20395 32827
rect 24685 32793 24719 32827
rect 31309 32793 31343 32827
rect 40049 32793 40083 32827
rect 5273 32725 5307 32759
rect 13645 32725 13679 32759
rect 20545 32725 20579 32759
rect 21097 32725 21131 32759
rect 25145 32725 25179 32759
rect 30941 32725 30975 32759
rect 31401 32725 31435 32759
rect 43821 32725 43855 32759
rect 7849 32521 7883 32555
rect 8401 32521 8435 32555
rect 16497 32521 16531 32555
rect 27905 32521 27939 32555
rect 34069 32521 34103 32555
rect 35633 32521 35667 32555
rect 7113 32453 7147 32487
rect 16957 32453 16991 32487
rect 34529 32453 34563 32487
rect 35449 32453 35483 32487
rect 6193 32385 6227 32419
rect 6837 32385 6871 32419
rect 8033 32385 8067 32419
rect 8309 32385 8343 32419
rect 8493 32385 8527 32419
rect 10609 32385 10643 32419
rect 16313 32385 16347 32419
rect 19441 32385 19475 32419
rect 22293 32385 22327 32419
rect 24869 32385 24903 32419
rect 27997 32385 28031 32419
rect 30941 32385 30975 32419
rect 31125 32385 31159 32419
rect 34161 32385 34195 32419
rect 34437 32385 34471 32419
rect 34621 32385 34655 32419
rect 34805 32385 34839 32419
rect 35265 32385 35299 32419
rect 42073 32385 42107 32419
rect 43545 32385 43579 32419
rect 7297 32317 7331 32351
rect 10517 32317 10551 32351
rect 16681 32317 16715 32351
rect 18429 32317 18463 32351
rect 19073 32317 19107 32351
rect 19257 32317 19291 32351
rect 19625 32317 19659 32351
rect 25145 32317 25179 32351
rect 26617 32317 26651 32351
rect 6653 32249 6687 32283
rect 34989 32249 35023 32283
rect 6009 32181 6043 32215
rect 10977 32181 11011 32215
rect 18521 32181 18555 32215
rect 22201 32181 22235 32215
rect 31033 32181 31067 32215
rect 42257 32181 42291 32215
rect 43361 32181 43395 32215
rect 7205 31977 7239 32011
rect 7849 31977 7883 32011
rect 8125 31977 8159 32011
rect 11069 31977 11103 32011
rect 16773 31977 16807 32011
rect 19993 31977 20027 32011
rect 21281 31977 21315 32011
rect 25329 31977 25363 32011
rect 31585 31977 31619 32011
rect 34069 31977 34103 32011
rect 37013 31977 37047 32011
rect 37362 31977 37396 32011
rect 39865 31977 39899 32011
rect 41613 31977 41647 32011
rect 8033 31909 8067 31943
rect 12265 31909 12299 31943
rect 19625 31909 19659 31943
rect 20177 31909 20211 31943
rect 31033 31909 31067 31943
rect 41061 31909 41095 31943
rect 5457 31841 5491 31875
rect 5733 31841 5767 31875
rect 9321 31841 9355 31875
rect 17325 31841 17359 31875
rect 30205 31841 30239 31875
rect 30297 31841 30331 31875
rect 31953 31841 31987 31875
rect 37105 31841 37139 31875
rect 40509 31841 40543 31875
rect 42533 31841 42567 31875
rect 42809 31841 42843 31875
rect 44281 31841 44315 31875
rect 8953 31773 8987 31807
rect 9137 31773 9171 31807
rect 11253 31773 11287 31807
rect 11621 31773 11655 31807
rect 11714 31773 11748 31807
rect 11897 31773 11931 31807
rect 12127 31773 12161 31807
rect 15020 31773 15054 31807
rect 15117 31773 15151 31807
rect 15392 31773 15426 31807
rect 15485 31773 15519 31807
rect 17233 31773 17267 31807
rect 20913 31773 20947 31807
rect 21097 31773 21131 31807
rect 24685 31773 24719 31807
rect 24833 31773 24867 31807
rect 25053 31773 25087 31807
rect 25150 31773 25184 31807
rect 29746 31783 29780 31817
rect 29837 31773 29871 31807
rect 29929 31773 29963 31807
rect 30067 31773 30101 31807
rect 30849 31773 30883 31807
rect 31217 31773 31251 31807
rect 31493 31773 31527 31807
rect 31585 31773 31619 31807
rect 31861 31773 31895 31807
rect 32137 31773 32171 31807
rect 32229 31773 32263 31807
rect 36461 31773 36495 31807
rect 36645 31773 36679 31807
rect 36737 31773 36771 31807
rect 36853 31773 36887 31807
rect 40785 31773 40819 31807
rect 40877 31773 40911 31807
rect 41153 31773 41187 31807
rect 42165 31773 42199 31807
rect 7665 31705 7699 31739
rect 7865 31705 7899 31739
rect 8309 31705 8343 31739
rect 8493 31705 8527 31739
rect 9597 31705 9631 31739
rect 11989 31705 12023 31739
rect 15209 31705 15243 31739
rect 17141 31705 17175 31739
rect 20637 31705 20671 31739
rect 20821 31705 20855 31739
rect 24961 31705 24995 31739
rect 31401 31705 31435 31739
rect 31677 31705 31711 31739
rect 31953 31705 31987 31739
rect 34253 31705 34287 31739
rect 34437 31705 34471 31739
rect 9045 31637 9079 31671
rect 11345 31637 11379 31671
rect 14841 31637 14875 31671
rect 19993 31637 20027 31671
rect 20269 31637 20303 31671
rect 20453 31637 20487 31671
rect 20545 31637 20579 31671
rect 29561 31637 29595 31671
rect 38853 31637 38887 31671
rect 40601 31637 40635 31671
rect 6193 31433 6227 31467
rect 8493 31433 8527 31467
rect 9413 31433 9447 31467
rect 11989 31433 12023 31467
rect 35265 31433 35299 31467
rect 42073 31433 42107 31467
rect 42441 31433 42475 31467
rect 42901 31433 42935 31467
rect 5825 31365 5859 31399
rect 6041 31365 6075 31399
rect 8125 31365 8159 31399
rect 14565 31365 14599 31399
rect 14657 31365 14691 31399
rect 16313 31365 16347 31399
rect 20085 31365 20119 31399
rect 20821 31365 20855 31399
rect 25329 31365 25363 31399
rect 26341 31365 26375 31399
rect 26433 31365 26467 31399
rect 33793 31365 33827 31399
rect 38761 31365 38795 31399
rect 8309 31297 8343 31331
rect 8493 31297 8527 31331
rect 8769 31297 8803 31331
rect 8953 31297 8987 31331
rect 9045 31297 9079 31331
rect 9137 31297 9171 31331
rect 11897 31297 11931 31331
rect 13645 31297 13679 31331
rect 13921 31297 13955 31331
rect 14013 31297 14047 31331
rect 14197 31297 14231 31331
rect 14427 31297 14461 31331
rect 14840 31297 14874 31331
rect 14933 31297 14967 31331
rect 15209 31297 15243 31331
rect 15301 31297 15335 31331
rect 15761 31297 15795 31331
rect 16129 31297 16163 31331
rect 16405 31297 16439 31331
rect 18889 31297 18923 31331
rect 19073 31297 19107 31331
rect 19809 31297 19843 31331
rect 21097 31297 21131 31331
rect 21373 31297 21407 31331
rect 26244 31297 26278 31331
rect 26616 31297 26650 31331
rect 26709 31297 26743 31331
rect 28273 31297 28307 31331
rect 30389 31297 30423 31331
rect 30481 31297 30515 31331
rect 30665 31297 30699 31331
rect 30849 31297 30883 31331
rect 32965 31297 32999 31331
rect 33130 31297 33164 31331
rect 33241 31297 33275 31331
rect 33425 31307 33459 31341
rect 38485 31297 38519 31331
rect 40325 31297 40359 31331
rect 42809 31297 42843 31331
rect 13737 31229 13771 31263
rect 15577 31229 15611 31263
rect 15669 31229 15703 31263
rect 15945 31229 15979 31263
rect 16037 31229 16071 31263
rect 19717 31229 19751 31263
rect 20177 31229 20211 31263
rect 21557 31229 21591 31263
rect 22569 31229 22603 31263
rect 22845 31229 22879 31263
rect 25881 31229 25915 31263
rect 27537 31229 27571 31263
rect 28181 31229 28215 31263
rect 28549 31229 28583 31263
rect 30021 31229 30055 31263
rect 40601 31229 40635 31263
rect 43085 31229 43119 31263
rect 18981 31161 19015 31195
rect 21649 31161 21683 31195
rect 30573 31161 30607 31195
rect 33333 31161 33367 31195
rect 40233 31161 40267 31195
rect 6009 31093 6043 31127
rect 6837 31093 6871 31127
rect 13829 31093 13863 31127
rect 14289 31093 14323 31127
rect 15025 31093 15059 31127
rect 15945 31093 15979 31127
rect 19533 31093 19567 31127
rect 24317 31093 24351 31127
rect 26065 31093 26099 31127
rect 30205 31093 30239 31127
rect 32781 31093 32815 31127
rect 7481 30889 7515 30923
rect 8033 30889 8067 30923
rect 12817 30889 12851 30923
rect 14270 30889 14304 30923
rect 14381 30889 14415 30923
rect 14565 30889 14599 30923
rect 19533 30889 19567 30923
rect 20177 30889 20211 30923
rect 20453 30889 20487 30923
rect 20913 30889 20947 30923
rect 21373 30889 21407 30923
rect 22569 30889 22603 30923
rect 25697 30889 25731 30923
rect 34345 30889 34379 30923
rect 37289 30889 37323 30923
rect 38117 30889 38151 30923
rect 38945 30889 38979 30923
rect 40601 30889 40635 30923
rect 41797 30889 41831 30923
rect 7021 30821 7055 30855
rect 20085 30821 20119 30855
rect 22661 30821 22695 30855
rect 23489 30821 23523 30855
rect 29285 30821 29319 30855
rect 3801 30753 3835 30787
rect 4077 30753 4111 30787
rect 6009 30753 6043 30787
rect 6653 30753 6687 30787
rect 10425 30753 10459 30787
rect 10885 30753 10919 30787
rect 13737 30753 13771 30787
rect 14473 30753 14507 30787
rect 15393 30753 15427 30787
rect 18705 30753 18739 30787
rect 23305 30753 23339 30787
rect 24133 30753 24167 30787
rect 27169 30753 27203 30787
rect 27445 30753 27479 30787
rect 27537 30753 27571 30787
rect 33057 30753 33091 30787
rect 33701 30753 33735 30787
rect 33977 30753 34011 30787
rect 34805 30753 34839 30787
rect 41153 30753 41187 30787
rect 42349 30753 42383 30787
rect 44097 30753 44131 30787
rect 5917 30685 5951 30719
rect 6101 30685 6135 30719
rect 6837 30685 6871 30719
rect 7573 30685 7607 30719
rect 8033 30685 8067 30719
rect 8217 30685 8251 30719
rect 10517 30685 10551 30719
rect 11621 30685 11655 30719
rect 11714 30685 11748 30719
rect 11989 30685 12023 30719
rect 12086 30685 12120 30719
rect 12541 30685 12575 30719
rect 12633 30685 12667 30719
rect 13068 30685 13102 30719
rect 13185 30685 13219 30719
rect 13405 30685 13439 30719
rect 13553 30685 13587 30719
rect 13653 30679 13687 30713
rect 14933 30685 14967 30719
rect 15117 30685 15151 30719
rect 15209 30685 15243 30719
rect 15485 30685 15519 30719
rect 18337 30685 18371 30719
rect 18521 30685 18555 30719
rect 18797 30685 18831 30719
rect 18981 30685 19015 30719
rect 19717 30685 19751 30719
rect 19901 30685 19935 30719
rect 20361 30685 20395 30719
rect 20545 30685 20579 30719
rect 20821 30685 20855 30719
rect 21097 30685 21131 30719
rect 21189 30685 21223 30719
rect 21465 30685 21499 30719
rect 21925 30685 21959 30719
rect 22017 30685 22051 30719
rect 22109 30685 22143 30719
rect 22385 30685 22419 30719
rect 23857 30685 23891 30719
rect 24961 30685 24995 30719
rect 30205 30685 30239 30719
rect 30389 30685 30423 30719
rect 31309 30685 31343 30719
rect 34069 30685 34103 30719
rect 34897 30685 34931 30719
rect 35541 30685 35575 30719
rect 37933 30685 37967 30719
rect 38209 30685 38243 30719
rect 38301 30685 38335 30719
rect 38669 30685 38703 30719
rect 39129 30685 39163 30719
rect 39497 30685 39531 30719
rect 40417 30685 40451 30719
rect 41521 30685 41555 30719
rect 41613 30685 41647 30719
rect 41889 30685 41923 30719
rect 42073 30685 42107 30719
rect 5825 30617 5859 30651
rect 7113 30617 7147 30651
rect 7297 30617 7331 30651
rect 7757 30617 7791 30651
rect 11897 30617 11931 30651
rect 12817 30617 12851 30651
rect 13277 30617 13311 30651
rect 14105 30617 14139 30651
rect 19441 30617 19475 30651
rect 23029 30617 23063 30651
rect 24409 30617 24443 30651
rect 27813 30617 27847 30651
rect 31585 30617 31619 30651
rect 35817 30617 35851 30651
rect 38485 30617 38519 30651
rect 38577 30617 38611 30651
rect 39221 30617 39255 30651
rect 39313 30617 39347 30651
rect 7941 30549 7975 30583
rect 12265 30549 12299 30583
rect 12357 30549 12391 30583
rect 12909 30549 12943 30583
rect 22293 30549 22327 30583
rect 23121 30549 23155 30583
rect 23949 30549 23983 30583
rect 31217 30549 31251 30583
rect 33149 30549 33183 30583
rect 35265 30549 35299 30583
rect 38853 30549 38887 30583
rect 39865 30549 39899 30583
rect 41337 30549 41371 30583
rect 5641 30345 5675 30379
rect 6101 30345 6135 30379
rect 7389 30345 7423 30379
rect 9505 30345 9539 30379
rect 11989 30345 12023 30379
rect 20545 30345 20579 30379
rect 23949 30345 23983 30379
rect 27629 30345 27663 30379
rect 33326 30345 33360 30379
rect 34713 30345 34747 30379
rect 35633 30345 35667 30379
rect 38301 30345 38335 30379
rect 43085 30345 43119 30379
rect 5733 30277 5767 30311
rect 12449 30277 12483 30311
rect 13921 30277 13955 30311
rect 15209 30277 15243 30311
rect 20269 30277 20303 30311
rect 27261 30277 27295 30311
rect 27353 30277 27387 30311
rect 29469 30277 29503 30311
rect 32229 30277 32263 30311
rect 32505 30277 32539 30311
rect 33425 30277 33459 30311
rect 33885 30277 33919 30311
rect 39037 30277 39071 30311
rect 5963 30243 5997 30277
rect 5365 30209 5399 30243
rect 7481 30209 7515 30243
rect 10793 30209 10827 30243
rect 11897 30209 11931 30243
rect 12541 30209 12575 30243
rect 12817 30209 12851 30243
rect 12909 30209 12943 30243
rect 13645 30209 13679 30243
rect 15117 30209 15151 30243
rect 18521 30209 18555 30243
rect 18705 30209 18739 30243
rect 18973 30209 19007 30243
rect 19165 30209 19199 30243
rect 19349 30209 19383 30243
rect 19625 30209 19659 30243
rect 19901 30209 19935 30243
rect 20386 30209 20420 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 26985 30209 27019 30243
rect 27133 30209 27167 30243
rect 27450 30209 27484 30243
rect 29285 30209 29319 30243
rect 29561 30209 29595 30243
rect 29653 30209 29687 30243
rect 30021 30209 30055 30243
rect 32413 30209 32447 30243
rect 32597 30209 32631 30243
rect 32735 30209 32769 30243
rect 32873 30209 32907 30243
rect 33149 30209 33183 30243
rect 33241 30209 33275 30243
rect 33701 30209 33735 30243
rect 34069 30209 34103 30243
rect 34253 30209 34287 30243
rect 34437 30209 34471 30243
rect 35081 30209 35115 30243
rect 35265 30209 35299 30243
rect 35357 30209 35391 30243
rect 35449 30209 35483 30243
rect 36277 30209 36311 30243
rect 36461 30209 36495 30243
rect 37841 30209 37875 30243
rect 38117 30209 38151 30243
rect 38761 30209 38795 30243
rect 41889 30209 41923 30243
rect 5641 30141 5675 30175
rect 7757 30141 7791 30175
rect 8033 30141 8067 30175
rect 13185 30141 13219 30175
rect 13277 30141 13311 30175
rect 13553 30141 13587 30175
rect 14013 30141 14047 30175
rect 16681 30141 16715 30175
rect 16957 30141 16991 30175
rect 19441 30141 19475 30175
rect 19533 30141 19567 30175
rect 20177 30141 20211 30175
rect 20821 30141 20855 30175
rect 21005 30141 21039 30175
rect 22201 30141 22235 30175
rect 22477 30141 22511 30175
rect 24133 30141 24167 30175
rect 24409 30141 24443 30175
rect 25881 30141 25915 30175
rect 29101 30141 29135 30175
rect 29837 30141 29871 30175
rect 33609 30141 33643 30175
rect 34345 30141 34379 30175
rect 34713 30141 34747 30175
rect 35725 30141 35759 30175
rect 36737 30141 36771 30175
rect 37933 30141 37967 30175
rect 41153 30141 41187 30175
rect 42533 30141 42567 30175
rect 12633 30073 12667 30107
rect 19073 30073 19107 30107
rect 19809 30073 19843 30107
rect 37013 30073 37047 30107
rect 40509 30073 40543 30107
rect 5457 30005 5491 30039
rect 5917 30005 5951 30039
rect 10701 30005 10735 30039
rect 13369 30005 13403 30039
rect 18429 30005 18463 30039
rect 18613 30005 18647 30039
rect 20637 30005 20671 30039
rect 34529 30005 34563 30039
rect 36829 30005 36863 30039
rect 38117 30005 38151 30039
rect 40601 30005 40635 30039
rect 41337 30005 41371 30039
rect 5733 29801 5767 29835
rect 8217 29801 8251 29835
rect 12633 29801 12667 29835
rect 24225 29801 24259 29835
rect 27261 29801 27295 29835
rect 27629 29801 27663 29835
rect 33885 29801 33919 29835
rect 35541 29801 35575 29835
rect 38945 29801 38979 29835
rect 42625 29801 42659 29835
rect 11345 29733 11379 29767
rect 12173 29733 12207 29767
rect 39037 29733 39071 29767
rect 3801 29665 3835 29699
rect 8953 29665 8987 29699
rect 12725 29665 12759 29699
rect 15761 29665 15795 29699
rect 17785 29665 17819 29699
rect 24961 29665 24995 29699
rect 41153 29665 41187 29699
rect 43177 29665 43211 29699
rect 43269 29665 43303 29699
rect 5917 29597 5951 29631
rect 6101 29597 6135 29631
rect 7573 29597 7607 29631
rect 7757 29597 7791 29631
rect 7849 29597 7883 29631
rect 7941 29597 7975 29631
rect 11437 29597 11471 29631
rect 11529 29597 11563 29631
rect 11622 29597 11656 29631
rect 11805 29597 11839 29631
rect 11897 29597 11931 29631
rect 11994 29597 12028 29631
rect 12633 29597 12667 29631
rect 12909 29597 12943 29631
rect 17969 29597 18003 29631
rect 24041 29597 24075 29631
rect 24777 29597 24811 29631
rect 27261 29597 27295 29631
rect 27445 29597 27479 29631
rect 33977 29597 34011 29631
rect 34161 29597 34195 29631
rect 35265 29597 35299 29631
rect 38393 29597 38427 29631
rect 38761 29597 38795 29631
rect 39681 29597 39715 29631
rect 39865 29597 39899 29631
rect 40877 29597 40911 29631
rect 4077 29529 4111 29563
rect 6377 29529 6411 29563
rect 6561 29529 6595 29563
rect 16037 29529 16071 29563
rect 33517 29529 33551 29563
rect 33701 29529 33735 29563
rect 38577 29529 38611 29563
rect 38669 29529 38703 29563
rect 5549 29461 5583 29495
rect 6193 29461 6227 29495
rect 9597 29461 9631 29495
rect 13093 29461 13127 29495
rect 17509 29461 17543 29495
rect 17877 29461 17911 29495
rect 18337 29461 18371 29495
rect 24409 29461 24443 29495
rect 24869 29461 24903 29495
rect 34161 29461 34195 29495
rect 40509 29461 40543 29495
rect 42717 29461 42751 29495
rect 43085 29461 43119 29495
rect 4169 29257 4203 29291
rect 5349 29257 5383 29291
rect 5733 29257 5767 29291
rect 9229 29257 9263 29291
rect 11069 29257 11103 29291
rect 16681 29257 16715 29291
rect 17969 29257 18003 29291
rect 18061 29257 18095 29291
rect 20361 29257 20395 29291
rect 21005 29257 21039 29291
rect 27537 29257 27571 29291
rect 32137 29257 32171 29291
rect 33609 29257 33643 29291
rect 37473 29257 37507 29291
rect 5549 29189 5583 29223
rect 9597 29189 9631 29223
rect 20085 29189 20119 29223
rect 20269 29189 20303 29223
rect 20637 29189 20671 29223
rect 21189 29189 21223 29223
rect 21373 29189 21407 29223
rect 23029 29189 23063 29223
rect 34897 29189 34931 29223
rect 40417 29189 40451 29223
rect 42901 29189 42935 29223
rect 4353 29121 4387 29155
rect 5825 29121 5859 29155
rect 9045 29121 9079 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17141 29121 17175 29155
rect 17417 29121 17451 29155
rect 18245 29121 18279 29155
rect 19901 29121 19935 29155
rect 20545 29121 20579 29155
rect 20775 29121 20809 29155
rect 20913 29121 20947 29155
rect 27169 29121 27203 29155
rect 27905 29121 27939 29155
rect 30297 29121 30331 29155
rect 30481 29121 30515 29155
rect 30665 29121 30699 29155
rect 31309 29121 31343 29155
rect 31493 29121 31527 29155
rect 33425 29121 33459 29155
rect 33609 29121 33643 29155
rect 37657 29121 37691 29155
rect 37933 29121 37967 29155
rect 38669 29121 38703 29155
rect 42073 29121 42107 29155
rect 9321 29053 9355 29087
rect 27261 29053 27295 29087
rect 27629 29053 27663 29087
rect 32781 29053 32815 29087
rect 36553 29053 36587 29087
rect 37841 29053 37875 29087
rect 40693 29053 40727 29087
rect 43453 29053 43487 29087
rect 5181 28985 5215 29019
rect 28089 28985 28123 29019
rect 31401 28985 31435 29019
rect 34621 28985 34655 29019
rect 38025 28985 38059 29019
rect 5365 28917 5399 28951
rect 24501 28917 24535 28951
rect 27721 28917 27755 28951
rect 36001 28917 36035 28951
rect 37933 28917 37967 28951
rect 38945 28917 38979 28951
rect 42257 28917 42291 28951
rect 7113 28713 7147 28747
rect 8401 28713 8435 28747
rect 9137 28713 9171 28747
rect 9321 28713 9355 28747
rect 11529 28713 11563 28747
rect 14749 28713 14783 28747
rect 20085 28713 20119 28747
rect 20821 28713 20855 28747
rect 29101 28713 29135 28747
rect 33977 28713 34011 28747
rect 37381 28713 37415 28747
rect 42165 28713 42199 28747
rect 6929 28645 6963 28679
rect 8585 28645 8619 28679
rect 13553 28645 13587 28679
rect 27997 28645 28031 28679
rect 32137 28645 32171 28679
rect 11253 28577 11287 28611
rect 14473 28577 14507 28611
rect 22753 28577 22787 28611
rect 27537 28577 27571 28611
rect 27813 28577 27847 28611
rect 31217 28577 31251 28611
rect 31677 28577 31711 28611
rect 32965 28577 32999 28611
rect 35909 28577 35943 28611
rect 40417 28577 40451 28611
rect 44281 28577 44315 28611
rect 6653 28509 6687 28543
rect 6837 28509 6871 28543
rect 7389 28509 7423 28543
rect 8309 28509 8343 28543
rect 8585 28509 8619 28543
rect 8769 28509 8803 28543
rect 9413 28509 9447 28543
rect 9597 28509 9631 28543
rect 11161 28509 11195 28543
rect 11989 28509 12023 28543
rect 12817 28509 12851 28543
rect 13185 28509 13219 28543
rect 13369 28509 13403 28543
rect 14381 28509 14415 28543
rect 16405 28509 16439 28543
rect 18521 28509 18555 28543
rect 19809 28509 19843 28543
rect 20367 28509 20401 28543
rect 20545 28509 20579 28543
rect 20913 28509 20947 28543
rect 23029 28509 23063 28543
rect 23949 28509 23983 28543
rect 24225 28509 24259 28543
rect 27445 28509 27479 28543
rect 27905 28509 27939 28543
rect 28089 28509 28123 28543
rect 29009 28509 29043 28543
rect 29929 28509 29963 28543
rect 30113 28509 30147 28543
rect 30389 28509 30423 28543
rect 30481 28509 30515 28543
rect 31033 28509 31067 28543
rect 31585 28509 31619 28543
rect 31861 28509 31895 28543
rect 32045 28509 32079 28543
rect 32229 28509 32263 28543
rect 32321 28509 32355 28543
rect 33057 28509 33091 28543
rect 34069 28509 34103 28543
rect 35633 28509 35667 28543
rect 38485 28509 38519 28543
rect 39681 28509 39715 28543
rect 42257 28509 42291 28543
rect 7297 28441 7331 28475
rect 8979 28441 9013 28475
rect 9169 28441 9203 28475
rect 9505 28441 9539 28475
rect 20085 28441 20119 28475
rect 20453 28441 20487 28475
rect 24133 28441 24167 28475
rect 30021 28441 30055 28475
rect 30251 28441 30285 28475
rect 32505 28441 32539 28475
rect 40693 28441 40727 28475
rect 42533 28441 42567 28475
rect 6469 28373 6503 28407
rect 7097 28373 7131 28407
rect 7573 28373 7607 28407
rect 12081 28373 12115 28407
rect 12265 28373 12299 28407
rect 16957 28373 16991 28407
rect 17969 28373 18003 28407
rect 19901 28373 19935 28407
rect 22201 28373 22235 28407
rect 22569 28373 22603 28407
rect 22661 28373 22695 28407
rect 23673 28373 23707 28407
rect 23765 28373 23799 28407
rect 29745 28373 29779 28407
rect 32689 28373 32723 28407
rect 37841 28373 37875 28407
rect 39037 28373 39071 28407
rect 5917 28169 5951 28203
rect 8585 28169 8619 28203
rect 8753 28169 8787 28203
rect 9597 28169 9631 28203
rect 11529 28169 11563 28203
rect 11897 28169 11931 28203
rect 12449 28169 12483 28203
rect 13921 28169 13955 28203
rect 15761 28169 15795 28203
rect 17509 28169 17543 28203
rect 18153 28169 18187 28203
rect 19901 28169 19935 28203
rect 21557 28169 21591 28203
rect 21833 28169 21867 28203
rect 26433 28169 26467 28203
rect 30481 28169 30515 28203
rect 30941 28169 30975 28203
rect 31769 28169 31803 28203
rect 32229 28169 32263 28203
rect 35725 28169 35759 28203
rect 41153 28169 41187 28203
rect 7849 28101 7883 28135
rect 8953 28101 8987 28135
rect 9413 28101 9447 28135
rect 11989 28101 12023 28135
rect 12817 28101 12851 28135
rect 14289 28101 14323 28135
rect 23305 28101 23339 28135
rect 28917 28101 28951 28135
rect 30665 28101 30699 28135
rect 30830 28101 30864 28135
rect 40601 28101 40635 28135
rect 5365 28033 5399 28067
rect 5549 28033 5583 28067
rect 5641 28033 5675 28067
rect 5837 28033 5871 28067
rect 6101 28033 6135 28067
rect 6193 28033 6227 28067
rect 6377 28033 6411 28067
rect 7021 28033 7055 28067
rect 7297 28033 7331 28067
rect 7389 28033 7423 28067
rect 8309 28033 8343 28067
rect 9229 28033 9263 28067
rect 9505 28033 9539 28067
rect 9597 28033 9631 28067
rect 9689 28033 9723 28067
rect 9873 28033 9907 28067
rect 11345 28033 11379 28067
rect 12628 28033 12662 28067
rect 12725 28033 12759 28067
rect 13000 28033 13034 28067
rect 13093 28033 13127 28067
rect 13737 28033 13771 28067
rect 16405 28033 16439 28067
rect 16773 28033 16807 28067
rect 16865 28033 16899 28067
rect 17325 28033 17359 28067
rect 17601 28033 17635 28067
rect 18061 28033 18095 28067
rect 18521 28033 18555 28067
rect 19901 28033 19935 28067
rect 20269 28033 20303 28067
rect 20637 28033 20671 28067
rect 21649 28033 21683 28067
rect 24409 28033 24443 28067
rect 27353 28033 27387 28067
rect 28089 28033 28123 28067
rect 30941 28033 30975 28067
rect 31125 28033 31159 28067
rect 31401 28033 31435 28067
rect 31769 28033 31803 28067
rect 31953 28033 31987 28067
rect 32137 28033 32171 28067
rect 32321 28033 32355 28067
rect 33333 28033 33367 28067
rect 35541 28033 35575 28067
rect 35909 28033 35943 28067
rect 36001 28033 36035 28067
rect 36093 28033 36127 28067
rect 36277 28033 36311 28067
rect 42533 28033 42567 28067
rect 5917 27965 5951 27999
rect 7113 27965 7147 27999
rect 12173 27965 12207 27999
rect 14013 27965 14047 27999
rect 18337 27965 18371 27999
rect 19165 27965 19199 27999
rect 19993 27965 20027 27999
rect 23581 27965 23615 27999
rect 24685 27965 24719 27999
rect 24961 27965 24995 27999
rect 28365 27965 28399 27999
rect 28641 27965 28675 27999
rect 30389 27965 30423 27999
rect 31677 27965 31711 27999
rect 33609 27965 33643 27999
rect 35081 27965 35115 27999
rect 36921 27965 36955 27999
rect 37289 27965 37323 27999
rect 37565 27965 37599 27999
rect 39037 27965 39071 27999
rect 40877 27965 40911 27999
rect 41705 27965 41739 27999
rect 5825 27897 5859 27931
rect 17049 27897 17083 27931
rect 31585 27897 31619 27931
rect 35357 27897 35391 27931
rect 5365 27829 5399 27863
rect 7205 27829 7239 27863
rect 7757 27829 7791 27863
rect 8493 27829 8527 27863
rect 8769 27829 8803 27863
rect 9045 27829 9079 27863
rect 11161 27829 11195 27863
rect 15853 27829 15887 27863
rect 17141 27829 17175 27863
rect 17693 27829 17727 27863
rect 20177 27829 20211 27863
rect 20545 27829 20579 27863
rect 24593 27829 24627 27863
rect 27905 27829 27939 27863
rect 31493 27829 31527 27863
rect 36369 27829 36403 27863
rect 39129 27829 39163 27863
rect 44005 27829 44039 27863
rect 4984 27625 5018 27659
rect 6910 27625 6944 27659
rect 8401 27625 8435 27659
rect 10964 27625 10998 27659
rect 12449 27625 12483 27659
rect 12909 27625 12943 27659
rect 16773 27625 16807 27659
rect 19533 27625 19567 27659
rect 19717 27625 19751 27659
rect 19901 27625 19935 27659
rect 20269 27625 20303 27659
rect 23397 27625 23431 27659
rect 24225 27625 24259 27659
rect 25310 27625 25344 27659
rect 33333 27625 33367 27659
rect 14473 27557 14507 27591
rect 15945 27557 15979 27591
rect 18889 27557 18923 27591
rect 39313 27557 39347 27591
rect 40969 27557 41003 27591
rect 43177 27557 43211 27591
rect 4721 27489 4755 27523
rect 13553 27489 13587 27523
rect 15117 27489 15151 27523
rect 23581 27489 23615 27523
rect 25053 27489 25087 27523
rect 26801 27489 26835 27523
rect 34069 27489 34103 27523
rect 41429 27489 41463 27523
rect 42625 27489 42659 27523
rect 42717 27489 42751 27523
rect 1409 27421 1443 27455
rect 6653 27421 6687 27455
rect 10701 27421 10735 27455
rect 13093 27421 13127 27455
rect 13185 27421 13219 27455
rect 13461 27421 13495 27455
rect 14841 27421 14875 27455
rect 16221 27421 16255 27455
rect 16405 27421 16439 27455
rect 16589 27421 16623 27455
rect 16865 27421 16899 27455
rect 17141 27421 17175 27455
rect 19257 27421 19291 27455
rect 19809 27421 19843 27455
rect 21649 27421 21683 27455
rect 23857 27421 23891 27455
rect 24409 27421 24443 27455
rect 28365 27421 28399 27455
rect 30665 27421 30699 27455
rect 32781 27421 32815 27455
rect 33149 27421 33183 27455
rect 34897 27421 34931 27455
rect 36921 27421 36955 27455
rect 38761 27421 38795 27455
rect 39129 27421 39163 27455
rect 40509 27421 40543 27455
rect 41153 27421 41187 27455
rect 41245 27421 41279 27455
rect 41521 27421 41555 27455
rect 43821 27421 43855 27455
rect 44189 27421 44223 27455
rect 17417 27353 17451 27387
rect 21925 27353 21959 27387
rect 32965 27353 32999 27387
rect 33057 27353 33091 27387
rect 33425 27353 33459 27387
rect 35173 27353 35207 27387
rect 38945 27353 38979 27387
rect 39037 27353 39071 27387
rect 1593 27285 1627 27319
rect 6469 27285 6503 27319
rect 14933 27285 14967 27319
rect 17049 27285 17083 27319
rect 23765 27285 23799 27319
rect 24593 27285 24627 27319
rect 28917 27285 28951 27319
rect 31953 27285 31987 27319
rect 36645 27285 36679 27319
rect 38209 27285 38243 27319
rect 39865 27285 39899 27319
rect 42809 27285 42843 27319
rect 43269 27285 43303 27319
rect 44005 27285 44039 27319
rect 10333 27081 10367 27115
rect 18429 27081 18463 27115
rect 22017 27081 22051 27115
rect 24777 27081 24811 27115
rect 31861 27081 31895 27115
rect 32321 27081 32355 27115
rect 35633 27081 35667 27115
rect 37933 27081 37967 27115
rect 8861 27013 8895 27047
rect 16957 27013 16991 27047
rect 28457 27013 28491 27047
rect 28825 27013 28859 27047
rect 29331 27013 29365 27047
rect 31677 27013 31711 27047
rect 38209 27013 38243 27047
rect 38301 27013 38335 27047
rect 16497 26945 16531 26979
rect 20453 26945 20487 26979
rect 22201 26945 22235 26979
rect 24409 26945 24443 26979
rect 29009 26945 29043 26979
rect 29101 26945 29135 26979
rect 29193 26945 29227 26979
rect 29469 26945 29503 26979
rect 29561 26945 29595 26979
rect 29745 26945 29779 26979
rect 31493 26945 31527 26979
rect 32137 26945 32171 26979
rect 32321 26945 32355 26979
rect 34345 26945 34379 26979
rect 34529 26945 34563 26979
rect 34621 26945 34655 26979
rect 34713 26945 34747 26979
rect 36645 26945 36679 26979
rect 36737 26945 36771 26979
rect 37013 26945 37047 26979
rect 37289 26945 37323 26979
rect 37473 26945 37507 26979
rect 37565 26945 37599 26979
rect 37841 26945 37875 26979
rect 38117 26945 38151 26979
rect 38485 26945 38519 26979
rect 40877 26945 40911 26979
rect 41153 26945 41187 26979
rect 41245 26945 41279 26979
rect 44281 26945 44315 26979
rect 8585 26877 8619 26911
rect 16221 26877 16255 26911
rect 16681 26877 16715 26911
rect 20177 26877 20211 26911
rect 20361 26877 20395 26911
rect 24133 26877 24167 26911
rect 24317 26877 24351 26911
rect 26985 26877 27019 26911
rect 28733 26877 28767 26911
rect 29653 26877 29687 26911
rect 34989 26877 35023 26911
rect 40693 26877 40727 26911
rect 40969 26877 41003 26911
rect 41429 26877 41463 26911
rect 41521 26877 41555 26911
rect 42533 26877 42567 26911
rect 44005 26877 44039 26911
rect 34897 26809 34931 26843
rect 20821 26741 20855 26775
rect 36461 26741 36495 26775
rect 36921 26741 36955 26775
rect 37749 26741 37783 26775
rect 40141 26741 40175 26775
rect 42165 26741 42199 26775
rect 9689 26537 9723 26571
rect 19441 26537 19475 26571
rect 30113 26537 30147 26571
rect 37933 26537 37967 26571
rect 41968 26537 42002 26571
rect 43453 26537 43487 26571
rect 4997 26469 5031 26503
rect 12357 26469 12391 26503
rect 21281 26469 21315 26503
rect 29837 26469 29871 26503
rect 30757 26469 30791 26503
rect 35449 26469 35483 26503
rect 4905 26401 4939 26435
rect 12817 26401 12851 26435
rect 13001 26401 13035 26435
rect 14749 26401 14783 26435
rect 15853 26401 15887 26435
rect 20913 26401 20947 26435
rect 21189 26401 21223 26435
rect 23489 26401 23523 26435
rect 30481 26401 30515 26435
rect 33885 26401 33919 26435
rect 36737 26401 36771 26435
rect 40141 26401 40175 26435
rect 41705 26401 41739 26435
rect 5365 26333 5399 26367
rect 9045 26333 9079 26367
rect 9229 26333 9263 26367
rect 11161 26333 11195 26367
rect 12265 26333 12299 26367
rect 13829 26333 13863 26367
rect 14473 26333 14507 26367
rect 15209 26333 15243 26367
rect 17969 26333 18003 26367
rect 21465 26333 21499 26367
rect 28273 26333 28307 26367
rect 28365 26333 28399 26367
rect 28825 26333 28859 26367
rect 29101 26333 29135 26367
rect 29285 26333 29319 26367
rect 29653 26333 29687 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 30389 26333 30423 26367
rect 31493 26333 31527 26367
rect 33977 26333 34011 26367
rect 34253 26333 34287 26367
rect 34345 26333 34379 26367
rect 35265 26333 35299 26367
rect 36001 26333 36035 26367
rect 37105 26333 37139 26367
rect 38485 26333 38519 26367
rect 39865 26333 39899 26367
rect 9137 26265 9171 26299
rect 12725 26265 12759 26299
rect 13185 26265 13219 26299
rect 16221 26265 16255 26299
rect 23673 26265 23707 26299
rect 28181 26265 28215 26299
rect 28917 26265 28951 26299
rect 33609 26265 33643 26299
rect 34161 26265 34195 26299
rect 37749 26265 37783 26299
rect 12081 26197 12115 26231
rect 14105 26197 14139 26231
rect 14565 26197 14599 26231
rect 23581 26197 23615 26231
rect 24041 26197 24075 26231
rect 28457 26197 28491 26231
rect 32045 26197 32079 26231
rect 32137 26197 32171 26231
rect 34529 26197 34563 26231
rect 34713 26197 34747 26231
rect 36185 26197 36219 26231
rect 41613 26197 41647 26231
rect 10073 25993 10107 26027
rect 10241 25993 10275 26027
rect 13369 25993 13403 26027
rect 15853 25993 15887 26027
rect 22385 25993 22419 26027
rect 22661 25993 22695 26027
rect 28733 25993 28767 26027
rect 29377 25993 29411 26027
rect 30113 25993 30147 26027
rect 32689 25993 32723 26027
rect 35265 25993 35299 26027
rect 37105 25993 37139 26027
rect 42717 25993 42751 26027
rect 43177 25993 43211 26027
rect 9873 25925 9907 25959
rect 11897 25925 11931 25959
rect 25421 25925 25455 25959
rect 28549 25925 28583 25959
rect 28917 25925 28951 25959
rect 29285 25925 29319 25959
rect 29561 25925 29595 25959
rect 32413 25925 32447 25959
rect 32873 25925 32907 25959
rect 33793 25925 33827 25959
rect 35633 25925 35667 25959
rect 6561 25857 6595 25891
rect 9045 25857 9079 25891
rect 9781 25857 9815 25891
rect 10517 25857 10551 25891
rect 10701 25857 10735 25891
rect 10977 25857 11011 25891
rect 13553 25857 13587 25891
rect 13737 25857 13771 25891
rect 17509 25857 17543 25891
rect 22201 25857 22235 25891
rect 22477 25857 22511 25891
rect 23397 25857 23431 25891
rect 26157 25857 26191 25891
rect 28365 25857 28399 25891
rect 28641 25857 28675 25891
rect 28825 25857 28859 25891
rect 29101 25857 29135 25891
rect 29745 25857 29779 25891
rect 29837 25857 29871 25891
rect 32137 25857 32171 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 32781 25857 32815 25891
rect 35357 25857 35391 25891
rect 37841 25857 37875 25891
rect 41705 25857 41739 25891
rect 42809 25857 42843 25891
rect 43269 25857 43303 25891
rect 7205 25789 7239 25823
rect 7573 25789 7607 25823
rect 11621 25789 11655 25823
rect 14105 25789 14139 25823
rect 14381 25789 14415 25823
rect 17325 25789 17359 25823
rect 19349 25789 19383 25823
rect 19625 25789 19659 25823
rect 23213 25789 23247 25823
rect 23673 25789 23707 25823
rect 25881 25789 25915 25823
rect 28181 25789 28215 25823
rect 30113 25789 30147 25823
rect 33517 25789 33551 25823
rect 38117 25789 38151 25823
rect 38393 25789 38427 25823
rect 39865 25789 39899 25823
rect 39957 25789 39991 25823
rect 42625 25789 42659 25823
rect 10333 25721 10367 25755
rect 6377 25653 6411 25687
rect 9137 25653 9171 25687
rect 10057 25653 10091 25687
rect 10793 25653 10827 25687
rect 13921 25653 13955 25687
rect 21097 25653 21131 25687
rect 22017 25653 22051 25687
rect 25973 25653 26007 25687
rect 26341 25653 26375 25687
rect 29929 25653 29963 25687
rect 37289 25653 37323 25687
rect 40601 25653 40635 25687
rect 41153 25653 41187 25687
rect 43453 25653 43487 25687
rect 7941 25449 7975 25483
rect 10713 25449 10747 25483
rect 14289 25449 14323 25483
rect 18889 25449 18923 25483
rect 19993 25449 20027 25483
rect 23489 25449 23523 25483
rect 23581 25449 23615 25483
rect 26065 25449 26099 25483
rect 26709 25449 26743 25483
rect 28641 25449 28675 25483
rect 29193 25449 29227 25483
rect 29653 25449 29687 25483
rect 36632 25449 36666 25483
rect 38485 25449 38519 25483
rect 39405 25449 39439 25483
rect 40509 25449 40543 25483
rect 40969 25449 41003 25483
rect 40325 25381 40359 25415
rect 5825 25313 5859 25347
rect 6101 25313 6135 25347
rect 10977 25313 11011 25347
rect 11069 25313 11103 25347
rect 12817 25313 12851 25347
rect 17785 25313 17819 25347
rect 20729 25313 20763 25347
rect 21281 25313 21315 25347
rect 21741 25313 21775 25347
rect 22017 25313 22051 25347
rect 25697 25313 25731 25347
rect 26525 25313 26559 25347
rect 27169 25313 27203 25347
rect 27445 25313 27479 25347
rect 36369 25313 36403 25347
rect 39129 25313 39163 25347
rect 39865 25313 39899 25347
rect 43913 25313 43947 25347
rect 44189 25313 44223 25347
rect 7849 25245 7883 25279
rect 8033 25245 8067 25279
rect 14105 25245 14139 25279
rect 18613 25245 18647 25279
rect 18797 25245 18831 25279
rect 19257 25245 19291 25279
rect 20177 25245 20211 25279
rect 20361 25245 20395 25279
rect 20453 25245 20487 25279
rect 23765 25245 23799 25279
rect 24961 25245 24995 25279
rect 25789 25245 25823 25279
rect 26433 25245 26467 25279
rect 27077 25245 27111 25279
rect 28549 25245 28583 25279
rect 28733 25245 28767 25279
rect 28825 25245 28859 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 31769 25245 31803 25279
rect 32505 25245 32539 25279
rect 39589 25245 39623 25279
rect 40049 25245 40083 25279
rect 40141 25245 40175 25279
rect 40417 25245 40451 25279
rect 40693 25245 40727 25279
rect 40785 25245 40819 25279
rect 41061 25245 41095 25279
rect 8953 25177 8987 25211
rect 11345 25177 11379 25211
rect 17509 25177 17543 25211
rect 18061 25177 18095 25211
rect 29009 25177 29043 25211
rect 31677 25177 31711 25211
rect 7573 25109 7607 25143
rect 17141 25109 17175 25143
rect 17601 25109 17635 25143
rect 19441 25109 19475 25143
rect 24409 25109 24443 25143
rect 31953 25109 31987 25143
rect 38117 25109 38151 25143
rect 42441 25109 42475 25143
rect 11897 24905 11931 24939
rect 15577 24905 15611 24939
rect 16129 24905 16163 24939
rect 18429 24905 18463 24939
rect 25697 24905 25731 24939
rect 27721 24905 27755 24939
rect 32137 24905 32171 24939
rect 39405 24837 39439 24871
rect 10701 24769 10735 24803
rect 11989 24769 12023 24803
rect 13829 24769 13863 24803
rect 16681 24769 16715 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 22201 24769 22235 24803
rect 22477 24769 22511 24803
rect 25881 24769 25915 24803
rect 26157 24769 26191 24803
rect 26985 24769 27019 24803
rect 27261 24769 27295 24803
rect 27629 24769 27663 24803
rect 27813 24769 27847 24803
rect 31401 24769 31435 24803
rect 31585 24769 31619 24803
rect 31677 24769 31711 24803
rect 31769 24769 31803 24803
rect 33885 24769 33919 24803
rect 36185 24769 36219 24803
rect 36737 24769 36771 24803
rect 39497 24769 39531 24803
rect 44281 24769 44315 24803
rect 12173 24701 12207 24735
rect 14105 24701 14139 24735
rect 16221 24701 16255 24735
rect 16405 24701 16439 24735
rect 16957 24701 16991 24735
rect 22753 24701 22787 24735
rect 27169 24701 27203 24735
rect 33609 24701 33643 24735
rect 36645 24701 36679 24735
rect 39589 24701 39623 24735
rect 10885 24633 10919 24667
rect 11529 24633 11563 24667
rect 22385 24633 22419 24667
rect 25973 24633 26007 24667
rect 26065 24633 26099 24667
rect 27445 24633 27479 24667
rect 31953 24633 31987 24667
rect 36553 24633 36587 24667
rect 44097 24633 44131 24667
rect 15761 24565 15795 24599
rect 24225 24565 24259 24599
rect 27077 24565 27111 24599
rect 36921 24565 36955 24599
rect 39037 24565 39071 24599
rect 13369 24361 13403 24395
rect 14473 24361 14507 24395
rect 16865 24361 16899 24395
rect 22109 24361 22143 24395
rect 31125 24361 31159 24395
rect 42901 24361 42935 24395
rect 14197 24293 14231 24327
rect 19073 24293 19107 24327
rect 29561 24293 29595 24327
rect 11621 24225 11655 24259
rect 17325 24225 17359 24259
rect 19809 24225 19843 24259
rect 20637 24225 20671 24259
rect 22661 24225 22695 24259
rect 30205 24225 30239 24259
rect 30757 24225 30791 24259
rect 32781 24225 32815 24259
rect 34529 24225 34563 24259
rect 35265 24225 35299 24259
rect 40509 24225 40543 24259
rect 43085 24225 43119 24259
rect 14289 24157 14323 24191
rect 14657 24157 14691 24191
rect 14841 24157 14875 24191
rect 16681 24157 16715 24191
rect 21005 24157 21039 24191
rect 22477 24157 22511 24191
rect 24961 24157 24995 24191
rect 29561 24157 29595 24191
rect 29837 24157 29871 24191
rect 30113 24157 30147 24191
rect 30297 24157 30331 24191
rect 30389 24157 30423 24191
rect 30849 24157 30883 24191
rect 36921 24157 36955 24191
rect 37565 24157 37599 24191
rect 38853 24157 38887 24191
rect 40233 24157 40267 24191
rect 42809 24157 42843 24191
rect 11897 24089 11931 24123
rect 17601 24089 17635 24123
rect 19625 24089 19659 24123
rect 20085 24089 20119 24123
rect 33057 24089 33091 24123
rect 40785 24089 40819 24123
rect 15025 24021 15059 24055
rect 19257 24021 19291 24055
rect 19717 24021 19751 24055
rect 20821 24021 20855 24055
rect 22569 24021 22603 24055
rect 24409 24021 24443 24055
rect 29745 24021 29779 24055
rect 30481 24021 30515 24055
rect 34713 24021 34747 24055
rect 37105 24021 37139 24055
rect 37381 24021 37415 24055
rect 39037 24021 39071 24055
rect 40417 24021 40451 24055
rect 42257 24021 42291 24055
rect 43085 24021 43119 24055
rect 12081 23817 12115 23851
rect 12357 23817 12391 23851
rect 12725 23817 12759 23851
rect 15301 23817 15335 23851
rect 18153 23817 18187 23851
rect 25145 23817 25179 23851
rect 31401 23817 31435 23851
rect 33701 23817 33735 23851
rect 34437 23817 34471 23851
rect 40969 23817 41003 23851
rect 41429 23817 41463 23851
rect 20177 23749 20211 23783
rect 29745 23749 29779 23783
rect 34805 23749 34839 23783
rect 36829 23749 36863 23783
rect 39037 23749 39071 23783
rect 39405 23749 39439 23783
rect 41337 23749 41371 23783
rect 12265 23681 12299 23715
rect 15945 23681 15979 23715
rect 18337 23681 18371 23715
rect 26433 23681 26467 23715
rect 29561 23681 29595 23715
rect 30113 23681 30147 23715
rect 30481 23681 30515 23715
rect 30665 23681 30699 23715
rect 31033 23681 31067 23715
rect 31401 23681 31435 23715
rect 31585 23681 31619 23715
rect 33885 23681 33919 23715
rect 33977 23681 34011 23715
rect 34069 23681 34103 23715
rect 34187 23681 34221 23715
rect 34345 23681 34379 23715
rect 34621 23681 34655 23715
rect 34897 23681 34931 23715
rect 35081 23681 35115 23715
rect 42809 23681 42843 23715
rect 43269 23681 43303 23715
rect 43453 23681 43487 23715
rect 43545 23681 43579 23715
rect 12817 23613 12851 23647
rect 13001 23613 13035 23647
rect 13553 23613 13587 23647
rect 13829 23613 13863 23647
rect 19901 23613 19935 23647
rect 23213 23613 23247 23647
rect 37105 23613 37139 23647
rect 39129 23613 39163 23647
rect 41521 23613 41555 23647
rect 42901 23613 42935 23647
rect 43085 23613 43119 23647
rect 43361 23613 43395 23647
rect 34989 23545 35023 23579
rect 37749 23545 37783 23579
rect 15393 23477 15427 23511
rect 21649 23477 21683 23511
rect 22661 23477 22695 23511
rect 35357 23477 35391 23511
rect 40877 23477 40911 23511
rect 42441 23477 42475 23511
rect 14105 23273 14139 23307
rect 15577 23273 15611 23307
rect 21189 23273 21223 23307
rect 24225 23273 24259 23307
rect 29193 23273 29227 23307
rect 32229 23273 32263 23307
rect 33241 23273 33275 23307
rect 33425 23273 33459 23307
rect 14565 23205 14599 23239
rect 33793 23205 33827 23239
rect 11621 23137 11655 23171
rect 15025 23137 15059 23171
rect 15117 23137 15151 23171
rect 21005 23137 21039 23171
rect 21741 23137 21775 23171
rect 26617 23137 26651 23171
rect 27813 23137 27847 23171
rect 37013 23137 37047 23171
rect 37289 23137 37323 23171
rect 43177 23137 43211 23171
rect 10517 23069 10551 23103
rect 10793 23069 10827 23103
rect 11345 23069 11379 23103
rect 14289 23069 14323 23103
rect 14933 23069 14967 23103
rect 15485 23069 15519 23103
rect 17049 23069 17083 23103
rect 18153 23069 18187 23103
rect 19257 23069 19291 23103
rect 21557 23069 21591 23103
rect 22477 23069 22511 23103
rect 25605 23069 25639 23103
rect 25789 23069 25823 23103
rect 26801 23069 26835 23103
rect 28089 23069 28123 23103
rect 28825 23069 28859 23103
rect 29561 23069 29595 23103
rect 31953 23069 31987 23103
rect 32137 23069 32171 23103
rect 32321 23069 32355 23103
rect 33517 23069 33551 23103
rect 33609 23069 33643 23103
rect 33885 23069 33919 23103
rect 34069 23069 34103 23103
rect 35725 23069 35759 23103
rect 43085 23069 43119 23103
rect 18061 23001 18095 23035
rect 19533 23001 19567 23035
rect 22753 23001 22787 23035
rect 24501 23001 24535 23035
rect 28733 23001 28767 23035
rect 29009 23001 29043 23035
rect 29837 23001 29871 23035
rect 33057 23001 33091 23035
rect 33793 23001 33827 23035
rect 10333 22933 10367 22967
rect 10609 22933 10643 22967
rect 10977 22933 11011 22967
rect 11437 22933 11471 22967
rect 17325 22933 17359 22967
rect 21649 22933 21683 22967
rect 24593 22933 24627 22967
rect 26893 22933 26927 22967
rect 31309 22933 31343 22967
rect 31401 22933 31435 22967
rect 33257 22933 33291 22967
rect 34253 22933 34287 22967
rect 35173 22933 35207 22967
rect 38761 22933 38795 22967
rect 42717 22933 42751 22967
rect 11529 22729 11563 22763
rect 16497 22729 16531 22763
rect 19165 22729 19199 22763
rect 23029 22729 23063 22763
rect 23673 22729 23707 22763
rect 24685 22729 24719 22763
rect 25789 22729 25823 22763
rect 28181 22729 28215 22763
rect 29377 22729 29411 22763
rect 32597 22729 32631 22763
rect 32965 22729 32999 22763
rect 35357 22729 35391 22763
rect 37565 22729 37599 22763
rect 37933 22729 37967 22763
rect 9781 22661 9815 22695
rect 13369 22661 13403 22695
rect 16957 22661 16991 22695
rect 30113 22661 30147 22695
rect 32873 22661 32907 22695
rect 38025 22661 38059 22695
rect 40049 22661 40083 22695
rect 43361 22661 43395 22695
rect 11897 22593 11931 22627
rect 13277 22593 13311 22627
rect 16313 22593 16347 22627
rect 19809 22593 19843 22627
rect 22017 22593 22051 22627
rect 23213 22593 23247 22627
rect 24869 22593 24903 22627
rect 25421 22593 25455 22627
rect 26065 22593 26099 22627
rect 26341 22593 26375 22627
rect 28089 22591 28123 22625
rect 29561 22593 29595 22627
rect 29653 22593 29687 22627
rect 29745 22593 29779 22627
rect 29863 22593 29897 22627
rect 30021 22593 30055 22627
rect 30297 22593 30331 22627
rect 30481 22593 30515 22627
rect 30573 22593 30607 22627
rect 30665 22593 30699 22627
rect 30757 22593 30791 22627
rect 32137 22593 32171 22627
rect 32229 22593 32263 22627
rect 32413 22593 32447 22627
rect 32689 22593 32723 22627
rect 32965 22593 32999 22627
rect 33701 22593 33735 22627
rect 33885 22593 33919 22627
rect 34161 22593 34195 22627
rect 35081 22593 35115 22627
rect 37105 22593 37139 22627
rect 39589 22593 39623 22627
rect 40325 22593 40359 22627
rect 43085 22593 43119 22627
rect 9505 22525 9539 22559
rect 11253 22525 11287 22559
rect 11989 22525 12023 22559
rect 12173 22525 12207 22559
rect 13553 22525 13587 22559
rect 16681 22525 16715 22559
rect 18981 22525 19015 22559
rect 19073 22525 19107 22559
rect 23765 22525 23799 22559
rect 23949 22525 23983 22559
rect 25145 22525 25179 22559
rect 25513 22525 25547 22559
rect 25881 22525 25915 22559
rect 34989 22525 35023 22559
rect 36829 22525 36863 22559
rect 38117 22525 38151 22559
rect 39681 22525 39715 22559
rect 40049 22525 40083 22559
rect 43177 22525 43211 22559
rect 23305 22457 23339 22491
rect 26157 22457 26191 22491
rect 26249 22457 26283 22491
rect 39957 22457 39991 22491
rect 12909 22389 12943 22423
rect 18429 22389 18463 22423
rect 19533 22389 19567 22423
rect 19625 22389 19659 22423
rect 21833 22389 21867 22423
rect 25053 22389 25087 22423
rect 34345 22389 34379 22423
rect 34713 22389 34747 22423
rect 40233 22389 40267 22423
rect 42901 22389 42935 22423
rect 43361 22389 43395 22423
rect 10136 22185 10170 22219
rect 11621 22185 11655 22219
rect 13645 22185 13679 22219
rect 17601 22185 17635 22219
rect 21268 22185 21302 22219
rect 25329 22185 25363 22219
rect 25697 22185 25731 22219
rect 26525 22185 26559 22219
rect 26801 22185 26835 22219
rect 29929 22185 29963 22219
rect 40417 22185 40451 22219
rect 25881 22117 25915 22151
rect 40509 22117 40543 22151
rect 9873 22049 9907 22083
rect 11897 22049 11931 22083
rect 15393 22049 15427 22083
rect 18061 22049 18095 22083
rect 18245 22049 18279 22083
rect 22753 22049 22787 22083
rect 25605 22049 25639 22083
rect 35449 22049 35483 22083
rect 40325 22049 40359 22083
rect 41061 22049 41095 22083
rect 41153 22049 41187 22083
rect 41245 22049 41279 22083
rect 44097 22049 44131 22083
rect 17969 21981 18003 22015
rect 21005 21981 21039 22015
rect 24961 21981 24995 22015
rect 25421 21981 25455 22015
rect 25697 21981 25731 22015
rect 26341 21981 26375 22015
rect 28549 21981 28583 22015
rect 28733 21981 28767 22015
rect 29837 21981 29871 22015
rect 30113 21981 30147 22015
rect 30849 21981 30883 22015
rect 34713 21981 34747 22015
rect 34989 21981 35023 22015
rect 35081 21981 35115 22015
rect 35541 21981 35575 22015
rect 40417 21981 40451 22015
rect 40693 21981 40727 22015
rect 40785 21981 40819 22015
rect 41337 21981 41371 22015
rect 41521 21981 41555 22015
rect 41705 21981 41739 22015
rect 41797 21981 41831 22015
rect 42349 21981 42383 22015
rect 42625 21981 42659 22015
rect 42809 21981 42843 22015
rect 43177 21981 43211 22015
rect 43361 21981 43395 22015
rect 12173 21913 12207 21947
rect 15669 21913 15703 21947
rect 25145 21913 25179 21947
rect 28273 21913 28307 21947
rect 30941 21913 30975 21947
rect 34897 21913 34931 21947
rect 40509 21913 40543 21947
rect 17141 21845 17175 21879
rect 29009 21845 29043 21879
rect 35265 21845 35299 21879
rect 40049 21845 40083 21879
rect 40877 21845 40911 21879
rect 41619 21845 41653 21879
rect 42441 21845 42475 21879
rect 43453 21845 43487 21879
rect 12449 21641 12483 21675
rect 15853 21641 15887 21675
rect 17509 21641 17543 21675
rect 21925 21641 21959 21675
rect 22293 21641 22327 21675
rect 28365 21641 28399 21675
rect 43453 21641 43487 21675
rect 21649 21573 21683 21607
rect 33793 21573 33827 21607
rect 39865 21573 39899 21607
rect 39957 21573 39991 21607
rect 8125 21505 8159 21539
rect 12633 21505 12667 21539
rect 13093 21505 13127 21539
rect 13369 21505 13403 21539
rect 16037 21505 16071 21539
rect 18797 21505 18831 21539
rect 19625 21505 19659 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 25881 21505 25915 21539
rect 26065 21505 26099 21539
rect 27721 21505 27755 21539
rect 28549 21505 28583 21539
rect 28641 21505 28675 21539
rect 28733 21505 28767 21539
rect 28917 21505 28951 21539
rect 31953 21505 31987 21539
rect 34253 21505 34287 21539
rect 34437 21505 34471 21539
rect 38669 21505 38703 21539
rect 38761 21505 38795 21539
rect 38945 21505 38979 21539
rect 39773 21505 39807 21539
rect 40141 21505 40175 21539
rect 40233 21505 40267 21539
rect 40601 21505 40635 21539
rect 40785 21505 40819 21539
rect 41245 21505 41279 21539
rect 41613 21505 41647 21539
rect 42809 21505 42843 21539
rect 42901 21505 42935 21539
rect 43269 21505 43303 21539
rect 43545 21505 43579 21539
rect 13645 21437 13679 21471
rect 15393 21437 15427 21471
rect 19901 21437 19935 21471
rect 22569 21437 22603 21471
rect 28273 21437 28307 21471
rect 38853 21437 38887 21471
rect 39681 21437 39715 21471
rect 40877 21437 40911 21471
rect 41337 21437 41371 21471
rect 41521 21437 41555 21471
rect 42073 21437 42107 21471
rect 42717 21437 42751 21471
rect 42993 21437 43027 21471
rect 13277 21369 13311 21403
rect 34069 21369 34103 21403
rect 41981 21369 42015 21403
rect 6837 21301 6871 21335
rect 23121 21301 23155 21335
rect 25973 21301 26007 21335
rect 30665 21301 30699 21335
rect 34345 21301 34379 21335
rect 39129 21301 39163 21335
rect 40417 21301 40451 21335
rect 43177 21301 43211 21335
rect 43269 21301 43303 21335
rect 14105 21097 14139 21131
rect 16681 21097 16715 21131
rect 20453 21097 20487 21131
rect 24225 21097 24259 21131
rect 29101 21097 29135 21131
rect 29193 21097 29227 21131
rect 33241 21097 33275 21131
rect 40233 21097 40267 21131
rect 41337 21097 41371 21131
rect 43177 21097 43211 21131
rect 20729 21029 20763 21063
rect 28365 21029 28399 21063
rect 32413 21029 32447 21063
rect 38485 21029 38519 21063
rect 43361 21029 43395 21063
rect 8953 20961 8987 20995
rect 14749 20961 14783 20995
rect 17325 20961 17359 20995
rect 21281 20961 21315 20995
rect 22477 20961 22511 20995
rect 22753 20961 22787 20995
rect 25881 20961 25915 20995
rect 26157 20961 26191 20995
rect 29009 20961 29043 20995
rect 31769 20961 31803 20995
rect 32137 20961 32171 20995
rect 39405 20961 39439 20995
rect 42257 20961 42291 20995
rect 43269 20961 43303 20995
rect 14473 20893 14507 20927
rect 17049 20893 17083 20927
rect 18521 20893 18555 20927
rect 20637 20893 20671 20927
rect 21097 20893 21131 20927
rect 25789 20893 25823 20927
rect 28549 20893 28583 20927
rect 28641 20893 28675 20927
rect 28733 20893 28767 20927
rect 28825 20893 28859 20927
rect 29285 20893 29319 20927
rect 30205 20893 30239 20927
rect 30389 20893 30423 20927
rect 31125 20893 31159 20927
rect 31309 20893 31343 20927
rect 31585 20893 31619 20927
rect 32045 20893 32079 20927
rect 32505 20893 32539 20927
rect 32781 20893 32815 20927
rect 33149 20893 33183 20927
rect 33333 20893 33367 20927
rect 33425 20893 33459 20927
rect 33609 20893 33643 20927
rect 33701 20893 33735 20927
rect 33885 20893 33919 20927
rect 34529 20893 34563 20927
rect 34897 20893 34931 20927
rect 34989 20893 35023 20927
rect 35357 20893 35391 20927
rect 36001 20893 36035 20927
rect 36645 20893 36679 20927
rect 38209 20893 38243 20927
rect 38301 20893 38335 20927
rect 38761 20893 38795 20927
rect 38945 20893 38979 20927
rect 39497 20893 39531 20927
rect 39865 20893 39899 20927
rect 40233 20893 40267 20927
rect 40417 20893 40451 20927
rect 41429 20893 41463 20927
rect 41705 20893 41739 20927
rect 42165 20893 42199 20927
rect 42533 20893 42567 20927
rect 42625 20893 42659 20927
rect 42993 20893 43027 20927
rect 43361 20893 43395 20927
rect 43637 20893 43671 20927
rect 29561 20825 29595 20859
rect 29745 20825 29779 20859
rect 29929 20825 29963 20859
rect 30021 20825 30055 20859
rect 32597 20825 32631 20859
rect 33517 20825 33551 20859
rect 34161 20825 34195 20859
rect 34345 20825 34379 20859
rect 35081 20825 35115 20859
rect 35199 20825 35233 20859
rect 38485 20825 38519 20859
rect 41889 20825 41923 20859
rect 43545 20825 43579 20859
rect 9597 20757 9631 20791
rect 14565 20757 14599 20791
rect 17141 20757 17175 20791
rect 18337 20757 18371 20791
rect 21189 20757 21223 20791
rect 32965 20757 32999 20791
rect 34069 20757 34103 20791
rect 34713 20757 34747 20791
rect 40049 20757 40083 20791
rect 42809 20757 42843 20791
rect 11529 20553 11563 20587
rect 11897 20553 11931 20587
rect 14933 20553 14967 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 19717 20553 19751 20587
rect 23121 20553 23155 20587
rect 23489 20553 23523 20587
rect 28825 20553 28859 20587
rect 36645 20553 36679 20587
rect 37289 20553 37323 20587
rect 37749 20553 37783 20587
rect 39589 20553 39623 20587
rect 42625 20553 42659 20587
rect 18245 20485 18279 20519
rect 30573 20485 30607 20519
rect 33517 20485 33551 20519
rect 35173 20485 35207 20519
rect 39405 20485 39439 20519
rect 42809 20485 42843 20519
rect 10885 20417 10919 20451
rect 11989 20417 12023 20451
rect 13277 20417 13311 20451
rect 15301 20417 15335 20451
rect 17969 20417 18003 20451
rect 21005 20417 21039 20451
rect 28457 20417 28491 20451
rect 28733 20417 28767 20451
rect 28917 20417 28951 20451
rect 29009 20417 29043 20451
rect 29561 20417 29595 20451
rect 30113 20417 30147 20451
rect 30205 20417 30239 20451
rect 30389 20417 30423 20451
rect 30849 20417 30883 20451
rect 31309 20417 31343 20451
rect 33425 20417 33459 20451
rect 33609 20417 33643 20451
rect 33701 20417 33735 20451
rect 33885 20417 33919 20451
rect 33977 20417 34011 20451
rect 34069 20417 34103 20451
rect 34437 20417 34471 20451
rect 34621 20417 34655 20451
rect 36921 20417 36955 20451
rect 37657 20417 37691 20451
rect 38117 20417 38151 20451
rect 38669 20417 38703 20451
rect 39037 20417 39071 20451
rect 39221 20417 39255 20451
rect 39681 20417 39715 20451
rect 42533 20417 42567 20451
rect 12081 20349 12115 20383
rect 14289 20349 14323 20383
rect 16037 20349 16071 20383
rect 16221 20349 16255 20383
rect 23581 20349 23615 20383
rect 23765 20349 23799 20383
rect 28273 20349 28307 20383
rect 30573 20349 30607 20383
rect 31401 20349 31435 20383
rect 34897 20349 34931 20383
rect 37841 20349 37875 20383
rect 39313 20349 39347 20383
rect 28641 20281 28675 20315
rect 31677 20281 31711 20315
rect 36737 20281 36771 20315
rect 39405 20281 39439 20315
rect 10701 20213 10735 20247
rect 13093 20213 13127 20247
rect 15485 20213 15519 20247
rect 20821 20213 20855 20247
rect 30757 20213 30791 20247
rect 34345 20213 34379 20247
rect 34529 20213 34563 20247
rect 38853 20213 38887 20247
rect 42809 20213 42843 20247
rect 10412 20009 10446 20043
rect 11897 20009 11931 20043
rect 13921 20009 13955 20043
rect 15472 20009 15506 20043
rect 17509 20009 17543 20043
rect 18153 20009 18187 20043
rect 19257 20009 19291 20043
rect 25513 20009 25547 20043
rect 30021 20009 30055 20043
rect 30205 20009 30239 20043
rect 31033 20009 31067 20043
rect 37933 20009 37967 20043
rect 38853 20009 38887 20043
rect 6193 19941 6227 19975
rect 14105 19941 14139 19975
rect 29193 19941 29227 19975
rect 29929 19941 29963 19975
rect 39405 19941 39439 19975
rect 10149 19873 10183 19907
rect 12173 19873 12207 19907
rect 12449 19873 12483 19907
rect 14749 19873 14783 19907
rect 15209 19873 15243 19907
rect 19809 19873 19843 19907
rect 25237 19873 25271 19907
rect 26065 19873 26099 19907
rect 27905 19873 27939 19907
rect 28273 19873 28307 19907
rect 28641 19873 28675 19907
rect 29561 19873 29595 19907
rect 32321 19873 32355 19907
rect 36461 19873 36495 19907
rect 38577 19873 38611 19907
rect 6377 19805 6411 19839
rect 14565 19805 14599 19839
rect 18613 19805 18647 19839
rect 19625 19805 19659 19839
rect 20545 19805 20579 19839
rect 25145 19805 25179 19839
rect 25605 19805 25639 19839
rect 25789 19805 25823 19839
rect 25973 19805 26007 19839
rect 27997 19805 28031 19839
rect 28457 19805 28491 19839
rect 28733 19805 28767 19839
rect 29193 19805 29227 19839
rect 29377 19805 29411 19839
rect 30113 19805 30147 19839
rect 31125 19805 31159 19839
rect 33609 19805 33643 19839
rect 33701 19805 33735 19839
rect 33977 19805 34011 19839
rect 34161 19805 34195 19839
rect 36185 19805 36219 19839
rect 38761 19805 38795 19839
rect 38945 19805 38979 19839
rect 39957 19805 39991 19839
rect 40141 19805 40175 19839
rect 40417 19805 40451 19839
rect 42901 19805 42935 19839
rect 6561 19737 6595 19771
rect 6929 19737 6963 19771
rect 7389 19737 7423 19771
rect 17233 19737 17267 19771
rect 17417 19737 17451 19771
rect 18245 19737 18279 19771
rect 20821 19737 20855 19771
rect 28365 19737 28399 19771
rect 32045 19737 32079 19771
rect 39037 19737 39071 19771
rect 42717 19737 42751 19771
rect 7113 19669 7147 19703
rect 14473 19669 14507 19703
rect 18429 19669 18463 19703
rect 19717 19669 19751 19703
rect 22293 19669 22327 19703
rect 27721 19669 27755 19703
rect 29101 19669 29135 19703
rect 33885 19669 33919 19703
rect 34069 19669 34103 19703
rect 38025 19669 38059 19703
rect 39497 19669 39531 19703
rect 42533 19669 42567 19703
rect 11253 19465 11287 19499
rect 16681 19465 16715 19499
rect 20913 19465 20947 19499
rect 21281 19465 21315 19499
rect 28733 19465 28767 19499
rect 28825 19465 28859 19499
rect 29929 19465 29963 19499
rect 39681 19465 39715 19499
rect 13461 19397 13495 19431
rect 18153 19397 18187 19431
rect 19901 19397 19935 19431
rect 24593 19397 24627 19431
rect 25697 19397 25731 19431
rect 29745 19397 29779 19431
rect 31401 19397 31435 19431
rect 32137 19397 32171 19431
rect 42625 19397 42659 19431
rect 2881 19329 2915 19363
rect 7297 19329 7331 19363
rect 9505 19329 9539 19363
rect 13185 19329 13219 19363
rect 14749 19329 14783 19363
rect 17877 19329 17911 19363
rect 21373 19329 21407 19363
rect 22201 19329 22235 19363
rect 22569 19329 22603 19363
rect 25881 19329 25915 19363
rect 25973 19329 26007 19363
rect 26985 19329 27019 19363
rect 29377 19329 29411 19363
rect 29561 19329 29595 19363
rect 31309 19329 31343 19363
rect 31493 19329 31527 19363
rect 31677 19329 31711 19363
rect 32689 19329 32723 19363
rect 33885 19329 33919 19363
rect 34253 19329 34287 19363
rect 34437 19329 34471 19363
rect 34529 19329 34563 19363
rect 34713 19329 34747 19363
rect 39497 19329 39531 19363
rect 42441 19329 42475 19363
rect 42717 19329 42751 19363
rect 42809 19329 42843 19363
rect 43269 19329 43303 19363
rect 43361 19329 43395 19363
rect 43545 19329 43579 19363
rect 43637 19329 43671 19363
rect 3157 19261 3191 19295
rect 4629 19261 4663 19295
rect 6653 19261 6687 19295
rect 7941 19261 7975 19295
rect 9781 19261 9815 19295
rect 15025 19261 15059 19295
rect 16497 19261 16531 19295
rect 17233 19261 17267 19295
rect 21557 19261 21591 19295
rect 22845 19261 22879 19295
rect 27261 19261 27295 19295
rect 34161 19261 34195 19295
rect 43085 19261 43119 19295
rect 22385 19193 22419 19227
rect 34069 19193 34103 19227
rect 34437 19193 34471 19227
rect 7389 19125 7423 19159
rect 25973 19125 26007 19159
rect 26157 19125 26191 19159
rect 31125 19125 31159 19159
rect 33701 19125 33735 19159
rect 34621 19125 34655 19159
rect 42993 19125 43027 19159
rect 6515 18921 6549 18955
rect 10885 18921 10919 18955
rect 15301 18921 15335 18955
rect 19257 18921 19291 18955
rect 22385 18921 22419 18955
rect 23765 18921 23799 18955
rect 25881 18921 25915 18955
rect 26341 18921 26375 18955
rect 32597 18921 32631 18955
rect 43361 18921 43395 18955
rect 1593 18853 1627 18887
rect 2053 18853 2087 18887
rect 35449 18853 35483 18887
rect 1777 18785 1811 18819
rect 8493 18785 8527 18819
rect 10333 18785 10367 18819
rect 16129 18785 16163 18819
rect 17325 18785 17359 18819
rect 19073 18785 19107 18819
rect 19809 18785 19843 18819
rect 21741 18785 21775 18819
rect 30849 18785 30883 18819
rect 31125 18785 31159 18819
rect 37473 18785 37507 18819
rect 37933 18785 37967 18819
rect 38301 18785 38335 18819
rect 41153 18785 41187 18819
rect 42165 18785 42199 18819
rect 42533 18785 42567 18819
rect 42625 18785 42659 18819
rect 1409 18717 1443 18751
rect 4721 18717 4755 18751
rect 5089 18717 5123 18751
rect 8125 18717 8159 18751
rect 8953 18717 8987 18751
rect 9505 18717 9539 18751
rect 10977 18717 11011 18751
rect 13001 18717 13035 18751
rect 15485 18717 15519 18751
rect 15945 18717 15979 18751
rect 16405 18717 16439 18751
rect 20729 18717 20763 18751
rect 22017 18717 22051 18751
rect 24409 18717 24443 18751
rect 26065 18717 26099 18751
rect 26157 18717 26191 18751
rect 34713 18717 34747 18751
rect 35633 18717 35667 18751
rect 35817 18717 35851 18751
rect 36001 18717 36035 18751
rect 38117 18717 38151 18751
rect 39129 18717 39163 18751
rect 39313 18717 39347 18751
rect 39497 18717 39531 18751
rect 40969 18717 41003 18751
rect 41245 18717 41279 18751
rect 41337 18717 41371 18751
rect 41521 18717 41555 18751
rect 41613 18717 41647 18751
rect 41981 18717 42015 18751
rect 42349 18717 42383 18751
rect 42717 18717 42751 18751
rect 42901 18717 42935 18751
rect 43085 18717 43119 18751
rect 10425 18649 10459 18683
rect 16681 18649 16715 18683
rect 17601 18649 17635 18683
rect 19625 18649 19659 18683
rect 22477 18649 22511 18683
rect 26341 18649 26375 18683
rect 35357 18649 35391 18683
rect 35725 18649 35759 18683
rect 37657 18649 37691 18683
rect 37841 18649 37875 18683
rect 38853 18649 38887 18683
rect 39037 18649 39071 18683
rect 39405 18649 39439 18683
rect 41797 18649 41831 18683
rect 43361 18649 43395 18683
rect 2237 18581 2271 18615
rect 6699 18581 6733 18615
rect 10517 18581 10551 18615
rect 12449 18581 12483 18615
rect 12817 18581 12851 18615
rect 15577 18581 15611 18615
rect 16037 18581 16071 18615
rect 19717 18581 19751 18615
rect 20085 18581 20119 18615
rect 21925 18581 21959 18615
rect 24593 18581 24627 18615
rect 38669 18581 38703 18615
rect 39681 18581 39715 18615
rect 40785 18581 40819 18615
rect 43177 18581 43211 18615
rect 2789 18377 2823 18411
rect 8125 18377 8159 18411
rect 10517 18377 10551 18411
rect 12357 18377 12391 18411
rect 18337 18377 18371 18411
rect 18889 18377 18923 18411
rect 19257 18377 19291 18411
rect 23121 18377 23155 18411
rect 23305 18377 23339 18411
rect 41337 18377 41371 18411
rect 43637 18377 43671 18411
rect 6653 18309 6687 18343
rect 8585 18309 8619 18343
rect 10333 18309 10367 18343
rect 12725 18309 12759 18343
rect 14473 18309 14507 18343
rect 22753 18309 22787 18343
rect 24777 18309 24811 18343
rect 25697 18309 25731 18343
rect 41705 18309 41739 18343
rect 2605 18241 2639 18275
rect 8309 18241 8343 18275
rect 10701 18241 10735 18275
rect 12449 18241 12483 18275
rect 16497 18241 16531 18275
rect 18521 18241 18555 18275
rect 25053 18241 25087 18275
rect 25513 18241 25547 18275
rect 26157 18241 26191 18275
rect 29653 18241 29687 18275
rect 29837 18241 29871 18275
rect 30113 18241 30147 18275
rect 36277 18241 36311 18275
rect 36829 18241 36863 18275
rect 37657 18241 37691 18275
rect 38025 18241 38059 18275
rect 38761 18241 38795 18275
rect 38945 18241 38979 18275
rect 39129 18241 39163 18275
rect 39313 18241 39347 18275
rect 39589 18241 39623 18275
rect 39773 18241 39807 18275
rect 41521 18241 41555 18275
rect 41613 18241 41647 18275
rect 41889 18241 41923 18275
rect 43361 18241 43395 18275
rect 3341 18173 3375 18207
rect 3709 18173 3743 18207
rect 5135 18173 5169 18207
rect 5549 18173 5583 18207
rect 6377 18173 6411 18207
rect 11805 18173 11839 18207
rect 19349 18173 19383 18207
rect 19441 18173 19475 18207
rect 19901 18173 19935 18207
rect 20177 18173 20211 18207
rect 22569 18173 22603 18207
rect 22661 18173 22695 18207
rect 26433 18173 26467 18207
rect 30205 18173 30239 18207
rect 30481 18173 30515 18207
rect 35817 18173 35851 18207
rect 36093 18173 36127 18207
rect 37749 18173 37783 18207
rect 38669 18173 38703 18207
rect 39037 18173 39071 18207
rect 44189 18173 44223 18207
rect 36553 18105 36587 18139
rect 6193 18037 6227 18071
rect 16313 18037 16347 18071
rect 21649 18037 21683 18071
rect 25881 18037 25915 18071
rect 25973 18037 26007 18071
rect 26341 18037 26375 18071
rect 29837 18037 29871 18071
rect 34345 18037 34379 18071
rect 37013 18037 37047 18071
rect 37381 18037 37415 18071
rect 39497 18037 39531 18071
rect 39681 18037 39715 18071
rect 42809 18037 42843 18071
rect 3617 17833 3651 17867
rect 11897 17833 11931 17867
rect 12633 17833 12667 17867
rect 20729 17833 20763 17867
rect 22477 17833 22511 17867
rect 27261 17833 27295 17867
rect 30757 17833 30791 17867
rect 38761 17833 38795 17867
rect 41613 17833 41647 17867
rect 22569 17765 22603 17799
rect 26065 17765 26099 17799
rect 26157 17765 26191 17799
rect 30205 17765 30239 17799
rect 33057 17765 33091 17799
rect 6101 17697 6135 17731
rect 6193 17697 6227 17731
rect 7941 17697 7975 17731
rect 9505 17697 9539 17731
rect 10057 17697 10091 17731
rect 13277 17697 13311 17731
rect 15945 17697 15979 17731
rect 17969 17697 18003 17731
rect 21557 17697 21591 17731
rect 21833 17697 21867 17731
rect 26433 17697 26467 17731
rect 26617 17697 26651 17731
rect 27169 17697 27203 17731
rect 29009 17697 29043 17731
rect 29377 17697 29411 17731
rect 29745 17697 29779 17731
rect 29837 17697 29871 17731
rect 29929 17697 29963 17731
rect 37289 17697 37323 17731
rect 44281 17697 44315 17731
rect 2973 17629 3007 17663
rect 8585 17629 8619 17663
rect 12449 17629 12483 17663
rect 13001 17629 13035 17663
rect 14565 17629 14599 17663
rect 20913 17629 20947 17663
rect 21373 17629 21407 17663
rect 23121 17629 23155 17663
rect 25973 17629 26007 17663
rect 26249 17629 26283 17663
rect 26709 17629 26743 17663
rect 27445 17629 27479 17663
rect 27711 17629 27745 17663
rect 27905 17629 27939 17663
rect 29193 17629 29227 17663
rect 29561 17629 29595 17663
rect 30021 17629 30055 17663
rect 30573 17629 30607 17663
rect 32781 17629 32815 17663
rect 32873 17629 32907 17663
rect 33149 17629 33183 17663
rect 37013 17629 37047 17663
rect 39589 17629 39623 17663
rect 39865 17629 39899 17663
rect 42257 17629 42291 17663
rect 42441 17629 42475 17663
rect 42533 17629 42567 17663
rect 5825 17561 5859 17595
rect 6469 17561 6503 17595
rect 10333 17561 10367 17595
rect 13829 17561 13863 17595
rect 16221 17561 16255 17595
rect 30389 17561 30423 17595
rect 35173 17561 35207 17595
rect 40141 17561 40175 17595
rect 42349 17561 42383 17595
rect 42809 17561 42843 17595
rect 4353 17493 4387 17527
rect 8033 17493 8067 17527
rect 8953 17493 8987 17527
rect 11805 17493 11839 17527
rect 13093 17493 13127 17527
rect 13553 17493 13587 17527
rect 14381 17493 14415 17527
rect 21005 17493 21039 17527
rect 21465 17493 21499 17527
rect 27077 17493 27111 17527
rect 27629 17493 27663 17527
rect 27813 17493 27847 17527
rect 32597 17493 32631 17527
rect 36461 17493 36495 17527
rect 39037 17493 39071 17527
rect 5365 17289 5399 17323
rect 6929 17289 6963 17323
rect 10701 17289 10735 17323
rect 11529 17289 11563 17323
rect 11897 17289 11931 17323
rect 16681 17289 16715 17323
rect 17049 17289 17083 17323
rect 29561 17289 29595 17323
rect 30113 17289 30147 17323
rect 39037 17289 39071 17323
rect 39221 17289 39255 17323
rect 39503 17289 39537 17323
rect 39589 17289 39623 17323
rect 43269 17289 43303 17323
rect 43437 17289 43471 17323
rect 7941 17221 7975 17255
rect 16405 17221 16439 17255
rect 20453 17221 20487 17255
rect 28089 17221 28123 17255
rect 37565 17221 37599 17255
rect 40017 17221 40051 17255
rect 40233 17221 40267 17255
rect 43637 17221 43671 17255
rect 4721 17153 4755 17187
rect 5825 17153 5859 17187
rect 7665 17153 7699 17187
rect 10885 17153 10919 17187
rect 17141 17153 17175 17187
rect 17509 17153 17543 17187
rect 21833 17153 21867 17187
rect 25973 17153 26007 17187
rect 27077 17153 27111 17187
rect 29745 17153 29779 17187
rect 30297 17153 30331 17187
rect 32137 17153 32171 17187
rect 32229 17153 32263 17187
rect 32413 17153 32447 17187
rect 32965 17153 32999 17187
rect 33241 17153 33275 17187
rect 33425 17153 33459 17187
rect 33517 17153 33551 17187
rect 33701 17153 33735 17187
rect 33977 17153 34011 17187
rect 34161 17153 34195 17187
rect 34253 17153 34287 17187
rect 34437 17153 34471 17187
rect 34713 17153 34747 17187
rect 37289 17153 37323 17187
rect 39129 17153 39163 17187
rect 39313 17153 39347 17187
rect 39405 17153 39439 17187
rect 39681 17153 39715 17187
rect 41797 17153 41831 17187
rect 42073 17153 42107 17187
rect 42257 17153 42291 17187
rect 42533 17153 42567 17187
rect 7573 17085 7607 17119
rect 9413 17085 9447 17119
rect 9965 17085 9999 17119
rect 11989 17085 12023 17119
rect 12173 17085 12207 17119
rect 14105 17085 14139 17119
rect 14381 17085 14415 17119
rect 15853 17085 15887 17119
rect 17233 17085 17267 17119
rect 18061 17085 18095 17119
rect 18429 17085 18463 17119
rect 18705 17085 18739 17119
rect 22109 17085 22143 17119
rect 23581 17085 23615 17119
rect 24225 17085 24259 17119
rect 26065 17085 26099 17119
rect 26801 17085 26835 17119
rect 29929 17085 29963 17119
rect 30021 17085 30055 17119
rect 30573 17085 30607 17119
rect 32597 17085 32631 17119
rect 34621 17085 34655 17119
rect 40601 17085 40635 17119
rect 41153 17085 41187 17119
rect 41981 17085 42015 17119
rect 43085 17085 43119 17119
rect 33149 17017 33183 17051
rect 34069 17017 34103 17051
rect 39865 17017 39899 17051
rect 5917 16949 5951 16983
rect 10609 16949 10643 16983
rect 16313 16949 16347 16983
rect 23673 16949 23707 16983
rect 30481 16949 30515 16983
rect 32689 16949 32723 16983
rect 33057 16949 33091 16983
rect 33885 16949 33919 16983
rect 34437 16949 34471 16983
rect 40049 16949 40083 16983
rect 41613 16949 41647 16983
rect 42073 16949 42107 16983
rect 43453 16949 43487 16983
rect 8953 16745 8987 16779
rect 13277 16745 13311 16779
rect 14565 16745 14599 16779
rect 17693 16745 17727 16779
rect 18705 16745 18739 16779
rect 21741 16745 21775 16779
rect 30389 16745 30423 16779
rect 32689 16745 32723 16779
rect 33241 16745 33275 16779
rect 39313 16745 39347 16779
rect 40509 16745 40543 16779
rect 42717 16745 42751 16779
rect 10425 16609 10459 16643
rect 10701 16609 10735 16643
rect 11437 16609 11471 16643
rect 13829 16609 13863 16643
rect 15209 16609 15243 16643
rect 15945 16609 15979 16643
rect 19809 16609 19843 16643
rect 22385 16609 22419 16643
rect 25053 16609 25087 16643
rect 27353 16609 27387 16643
rect 32321 16609 32355 16643
rect 34805 16609 34839 16643
rect 40969 16609 41003 16643
rect 14933 16541 14967 16575
rect 18889 16541 18923 16575
rect 19625 16541 19659 16575
rect 21557 16541 21591 16575
rect 22201 16541 22235 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 27261 16541 27295 16575
rect 29837 16541 29871 16575
rect 30021 16541 30055 16575
rect 30297 16541 30331 16575
rect 30573 16541 30607 16575
rect 30757 16541 30791 16575
rect 32413 16541 32447 16575
rect 33149 16541 33183 16575
rect 33333 16541 33367 16575
rect 34345 16541 34379 16575
rect 34529 16541 34563 16575
rect 34897 16541 34931 16575
rect 35541 16541 35575 16575
rect 39129 16541 39163 16575
rect 39313 16541 39347 16575
rect 6377 16473 6411 16507
rect 11713 16473 11747 16507
rect 16221 16473 16255 16507
rect 24869 16473 24903 16507
rect 30205 16473 30239 16507
rect 35357 16473 35391 16507
rect 40417 16473 40451 16507
rect 41245 16473 41279 16507
rect 7665 16405 7699 16439
rect 13185 16405 13219 16439
rect 15025 16405 15059 16439
rect 19257 16405 19291 16439
rect 19717 16405 19751 16439
rect 21833 16405 21867 16439
rect 22293 16405 22327 16439
rect 23673 16405 23707 16439
rect 24409 16405 24443 16439
rect 27629 16405 27663 16439
rect 30665 16405 30699 16439
rect 34345 16405 34379 16439
rect 35265 16405 35299 16439
rect 35725 16405 35759 16439
rect 2605 16201 2639 16235
rect 11897 16201 11931 16235
rect 12265 16201 12299 16235
rect 12633 16201 12667 16235
rect 16681 16201 16715 16235
rect 17141 16201 17175 16235
rect 17509 16201 17543 16235
rect 19441 16201 19475 16235
rect 19993 16201 20027 16235
rect 31401 16201 31435 16235
rect 4077 16133 4111 16167
rect 4813 16133 4847 16167
rect 9229 16133 9263 16167
rect 17601 16133 17635 16167
rect 25513 16133 25547 16167
rect 29653 16133 29687 16167
rect 30941 16133 30975 16167
rect 33149 16133 33183 16167
rect 42257 16133 42291 16167
rect 5917 16065 5951 16099
rect 8861 16065 8895 16099
rect 8953 16065 8987 16099
rect 12081 16065 12115 16099
rect 13277 16065 13311 16099
rect 16865 16065 16899 16099
rect 18153 16065 18187 16099
rect 23489 16065 23523 16099
rect 26985 16065 27019 16099
rect 29469 16065 29503 16099
rect 29561 16065 29595 16099
rect 29791 16065 29825 16099
rect 31106 16065 31140 16099
rect 31207 16065 31241 16099
rect 31401 16065 31435 16099
rect 31493 16063 31527 16097
rect 31677 16065 31711 16099
rect 31953 16065 31987 16099
rect 32137 16065 32171 16099
rect 33031 16065 33065 16099
rect 33241 16065 33275 16099
rect 33333 16065 33367 16099
rect 33793 16065 33827 16099
rect 33885 16065 33919 16099
rect 33977 16065 34011 16099
rect 34095 16065 34129 16099
rect 39865 16065 39899 16099
rect 40509 16065 40543 16099
rect 42441 16065 42475 16099
rect 44005 16065 44039 16099
rect 4353 15997 4387 16031
rect 5365 15997 5399 16031
rect 6009 15997 6043 16031
rect 7067 15997 7101 16031
rect 8493 15997 8527 16031
rect 12725 15997 12759 16031
rect 12909 15997 12943 16031
rect 13553 15997 13587 16031
rect 15025 15997 15059 16031
rect 15669 15997 15703 16031
rect 17693 15997 17727 16031
rect 20545 15997 20579 16031
rect 23765 15997 23799 16031
rect 29929 15997 29963 16031
rect 30021 15997 30055 16031
rect 30573 15997 30607 16031
rect 30757 15997 30791 16031
rect 32781 15997 32815 16031
rect 32873 15997 32907 16031
rect 34253 15997 34287 16031
rect 34345 15997 34379 16031
rect 34897 15997 34931 16031
rect 39957 15997 39991 16031
rect 42993 15997 43027 16031
rect 31861 15929 31895 15963
rect 5549 15861 5583 15895
rect 10701 15861 10735 15895
rect 15117 15861 15151 15895
rect 27169 15861 27203 15895
rect 29285 15861 29319 15895
rect 31585 15861 31619 15895
rect 33517 15861 33551 15895
rect 33609 15861 33643 15895
rect 40233 15861 40267 15895
rect 44189 15861 44223 15895
rect 5411 15657 5445 15691
rect 11989 15657 12023 15691
rect 13737 15657 13771 15691
rect 26709 15657 26743 15691
rect 29377 15657 29411 15691
rect 30573 15657 30607 15691
rect 32873 15657 32907 15691
rect 33517 15657 33551 15691
rect 34253 15657 34287 15691
rect 41981 15657 42015 15691
rect 21833 15589 21867 15623
rect 26801 15589 26835 15623
rect 36277 15589 36311 15623
rect 41705 15589 41739 15623
rect 1869 15521 1903 15555
rect 3617 15521 3651 15555
rect 4353 15521 4387 15555
rect 5273 15521 5307 15555
rect 7205 15521 7239 15555
rect 10241 15521 10275 15555
rect 12725 15521 12759 15555
rect 14657 15521 14691 15555
rect 19901 15521 19935 15555
rect 22477 15521 22511 15555
rect 24225 15521 24259 15555
rect 24409 15521 24443 15555
rect 26157 15521 26191 15555
rect 27629 15521 27663 15555
rect 27905 15521 27939 15555
rect 32045 15521 32079 15555
rect 37749 15521 37783 15555
rect 38025 15521 38059 15555
rect 39221 15521 39255 15555
rect 39957 15521 39991 15555
rect 40233 15521 40267 15555
rect 42533 15521 42567 15555
rect 6837 15453 6871 15487
rect 12449 15453 12483 15487
rect 13921 15453 13955 15487
rect 14473 15453 14507 15487
rect 18705 15453 18739 15487
rect 20085 15453 20119 15487
rect 22201 15453 22235 15487
rect 26341 15453 26375 15487
rect 27353 15453 27387 15487
rect 32321 15453 32355 15487
rect 33057 15453 33091 15487
rect 33333 15453 33367 15487
rect 33609 15453 33643 15487
rect 33701 15453 33735 15487
rect 34345 15453 34379 15487
rect 35357 15453 35391 15487
rect 35541 15453 35575 15487
rect 38853 15453 38887 15487
rect 39313 15453 39347 15487
rect 41797 15453 41831 15487
rect 41981 15453 42015 15487
rect 2145 15385 2179 15419
rect 10517 15385 10551 15419
rect 19625 15385 19659 15419
rect 20361 15385 20395 15419
rect 22753 15385 22787 15419
rect 33425 15385 33459 15419
rect 42809 15385 42843 15419
rect 3801 15317 3835 15351
rect 4629 15317 4663 15351
rect 12081 15317 12115 15351
rect 12541 15317 12575 15351
rect 14105 15317 14139 15351
rect 14565 15317 14599 15351
rect 18521 15317 18555 15351
rect 19257 15317 19291 15351
rect 19717 15317 19751 15351
rect 22385 15317 22419 15351
rect 25053 15317 25087 15351
rect 26249 15317 26283 15351
rect 33241 15317 33275 15351
rect 35449 15317 35483 15351
rect 38209 15317 38243 15351
rect 38945 15317 38979 15351
rect 44281 15317 44315 15351
rect 5917 15113 5951 15147
rect 10885 15113 10919 15147
rect 19625 15113 19659 15147
rect 20545 15113 20579 15147
rect 20913 15113 20947 15147
rect 21925 15113 21959 15147
rect 22753 15113 22787 15147
rect 39589 15113 39623 15147
rect 43545 15113 43579 15147
rect 3709 15045 3743 15079
rect 9045 15045 9079 15079
rect 22109 15045 22143 15079
rect 35357 15045 35391 15079
rect 38117 15045 38151 15079
rect 43637 15045 43671 15079
rect 3433 14977 3467 15011
rect 5549 14977 5583 15011
rect 8769 14977 8803 15011
rect 11069 14977 11103 15011
rect 17877 14977 17911 15011
rect 20361 14977 20395 15011
rect 20729 14977 20763 15011
rect 21281 14977 21315 15011
rect 21833 14977 21867 15011
rect 24961 14977 24995 15011
rect 32781 14977 32815 15011
rect 35081 14977 35115 15011
rect 37841 14977 37875 15011
rect 42993 14977 43027 15011
rect 43361 14977 43395 15011
rect 44281 14977 44315 15011
rect 5641 14909 5675 14943
rect 10517 14909 10551 14943
rect 18153 14909 18187 14943
rect 20177 14909 20211 14943
rect 21373 14909 21407 14943
rect 21557 14909 21591 14943
rect 22845 14909 22879 14943
rect 22937 14909 22971 14943
rect 25237 14909 25271 14943
rect 26709 14909 26743 14943
rect 27537 14909 27571 14943
rect 33057 14909 33091 14943
rect 42625 14909 42659 14943
rect 43085 14909 43119 14943
rect 22109 14841 22143 14875
rect 22385 14841 22419 14875
rect 26985 14841 27019 14875
rect 34529 14841 34563 14875
rect 5181 14773 5215 14807
rect 36829 14773 36863 14807
rect 12725 14569 12759 14603
rect 14197 14569 14231 14603
rect 16497 14569 16531 14603
rect 25237 14569 25271 14603
rect 34897 14569 34931 14603
rect 43269 14569 43303 14603
rect 11989 14501 12023 14535
rect 25697 14501 25731 14535
rect 26065 14501 26099 14535
rect 43085 14501 43119 14535
rect 43361 14501 43395 14535
rect 5365 14433 5399 14467
rect 14841 14433 14875 14467
rect 16313 14433 16347 14467
rect 16405 14433 16439 14467
rect 16589 14433 16623 14467
rect 27813 14433 27847 14467
rect 35173 14433 35207 14467
rect 37013 14433 37047 14467
rect 41337 14433 41371 14467
rect 43729 14433 43763 14467
rect 11897 14365 11931 14399
rect 12633 14365 12667 14399
rect 12909 14365 12943 14399
rect 13185 14365 13219 14399
rect 14565 14365 14599 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 16037 14365 16071 14399
rect 16129 14365 16163 14399
rect 16681 14365 16715 14399
rect 25421 14365 25455 14399
rect 25513 14365 25547 14399
rect 25789 14365 25823 14399
rect 31217 14365 31251 14399
rect 31401 14365 31435 14399
rect 34713 14365 34747 14399
rect 34897 14365 34931 14399
rect 35449 14365 35483 14399
rect 35725 14365 35759 14399
rect 36001 14365 36035 14399
rect 36369 14365 36403 14399
rect 14657 14297 14691 14331
rect 27537 14297 27571 14331
rect 36461 14297 36495 14331
rect 41613 14297 41647 14331
rect 6009 14229 6043 14263
rect 13093 14229 13127 14263
rect 31309 14229 31343 14263
rect 7849 14025 7883 14059
rect 12265 14025 12299 14059
rect 14565 14025 14599 14059
rect 15570 14025 15604 14059
rect 16681 14025 16715 14059
rect 18521 14025 18555 14059
rect 18797 14025 18831 14059
rect 21931 14025 21965 14059
rect 22017 14025 22051 14059
rect 22753 14025 22787 14059
rect 22845 14025 22879 14059
rect 36277 14025 36311 14059
rect 42441 14025 42475 14059
rect 15669 13957 15703 13991
rect 21833 13957 21867 13991
rect 23213 13957 23247 13991
rect 28089 13957 28123 13991
rect 31493 13957 31527 13991
rect 36429 13957 36463 13991
rect 36645 13957 36679 13991
rect 5733 13889 5767 13923
rect 7113 13889 7147 13923
rect 7297 13889 7331 13923
rect 7665 13889 7699 13923
rect 11989 13889 12023 13923
rect 12449 13889 12483 13923
rect 12541 13889 12575 13923
rect 12633 13889 12667 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 15393 13889 15427 13923
rect 15485 13889 15519 13923
rect 18061 13889 18095 13923
rect 18337 13889 18371 13923
rect 19073 13889 19107 13923
rect 19165 13889 19199 13923
rect 19258 13889 19292 13923
rect 22093 13889 22127 13923
rect 22477 13889 22511 13923
rect 23305 13889 23339 13923
rect 23949 13889 23983 13923
rect 29929 13889 29963 13923
rect 30159 13889 30193 13923
rect 30941 13889 30975 13923
rect 31217 13889 31251 13923
rect 31401 13889 31435 13923
rect 31769 13889 31803 13923
rect 34713 13889 34747 13923
rect 34897 13889 34931 13923
rect 34989 13889 35023 13923
rect 35817 13889 35851 13923
rect 40417 13889 40451 13923
rect 40509 13889 40543 13923
rect 43361 13889 43395 13923
rect 44189 13889 44223 13923
rect 4629 13821 4663 13855
rect 5365 13821 5399 13855
rect 5641 13821 5675 13855
rect 12265 13821 12299 13855
rect 14197 13821 14231 13855
rect 14381 13821 14415 13855
rect 16865 13821 16899 13855
rect 16957 13821 16991 13855
rect 17049 13821 17083 13855
rect 17141 13821 17175 13855
rect 18245 13821 18279 13855
rect 18977 13821 19011 13855
rect 22293 13821 22327 13855
rect 22385 13821 22419 13855
rect 22569 13821 22603 13855
rect 23397 13821 23431 13855
rect 29837 13821 29871 13855
rect 30297 13821 30331 13855
rect 30665 13821 30699 13855
rect 30757 13821 30791 13855
rect 31585 13821 31619 13855
rect 35633 13821 35667 13855
rect 40141 13821 40175 13855
rect 40785 13821 40819 13855
rect 42257 13821 42291 13855
rect 42993 13821 43027 13855
rect 7481 13753 7515 13787
rect 30067 13753 30101 13787
rect 44005 13753 44039 13787
rect 4077 13685 4111 13719
rect 6837 13685 6871 13719
rect 12081 13685 12115 13719
rect 18061 13685 18095 13719
rect 23765 13685 23799 13719
rect 31493 13685 31527 13719
rect 31953 13685 31987 13719
rect 34713 13685 34747 13719
rect 35909 13685 35943 13719
rect 36461 13685 36495 13719
rect 38669 13685 38703 13719
rect 43269 13685 43303 13719
rect 7435 13481 7469 13515
rect 11621 13481 11655 13515
rect 13737 13481 13771 13515
rect 14289 13481 14323 13515
rect 17141 13481 17175 13515
rect 17969 13481 18003 13515
rect 23489 13481 23523 13515
rect 25053 13481 25087 13515
rect 31033 13481 31067 13515
rect 34437 13481 34471 13515
rect 40693 13481 40727 13515
rect 40877 13481 40911 13515
rect 44097 13481 44131 13515
rect 18153 13413 18187 13447
rect 20729 13413 20763 13447
rect 20913 13413 20947 13447
rect 38393 13413 38427 13447
rect 3801 13345 3835 13379
rect 5641 13345 5675 13379
rect 7941 13345 7975 13379
rect 10885 13345 10919 13379
rect 11529 13345 11563 13379
rect 11621 13345 11655 13379
rect 16773 13345 16807 13379
rect 16957 13345 16991 13379
rect 17509 13345 17543 13379
rect 21833 13345 21867 13379
rect 22569 13345 22603 13379
rect 24133 13345 24167 13379
rect 27445 13345 27479 13379
rect 32505 13345 32539 13379
rect 34713 13345 34747 13379
rect 36185 13345 36219 13379
rect 36461 13345 36495 13379
rect 38301 13345 38335 13379
rect 39037 13345 39071 13379
rect 39129 13345 39163 13379
rect 39865 13345 39899 13379
rect 40509 13345 40543 13379
rect 42625 13345 42659 13379
rect 6009 13277 6043 13311
rect 8769 13277 8803 13311
rect 10149 13277 10183 13311
rect 11437 13277 11471 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 13553 13277 13587 13311
rect 14473 13277 14507 13311
rect 14657 13277 14691 13311
rect 14841 13277 14875 13311
rect 14933 13277 14967 13311
rect 16681 13277 16715 13311
rect 16865 13277 16899 13311
rect 17233 13277 17267 13311
rect 17417 13277 17451 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 18061 13277 18095 13311
rect 18245 13277 18279 13311
rect 20453 13277 20487 13311
rect 20913 13277 20947 13311
rect 21097 13277 21131 13311
rect 21649 13277 21683 13311
rect 22477 13277 22511 13311
rect 23029 13277 23063 13311
rect 23121 13277 23155 13311
rect 23213 13277 23247 13311
rect 23305 13277 23339 13311
rect 23765 13277 23799 13311
rect 23857 13277 23891 13311
rect 24225 13277 24259 13311
rect 24409 13277 24443 13311
rect 24593 13277 24627 13311
rect 24685 13277 24719 13311
rect 24777 13277 24811 13311
rect 29745 13277 29779 13311
rect 30021 13277 30055 13311
rect 30205 13277 30239 13311
rect 30297 13277 30331 13311
rect 30389 13277 30423 13311
rect 30573 13277 30607 13311
rect 30665 13277 30699 13311
rect 31217 13277 31251 13311
rect 31493 13277 31527 13311
rect 31677 13277 31711 13311
rect 32229 13277 32263 13311
rect 34161 13277 34195 13311
rect 39313 13277 39347 13311
rect 40601 13277 40635 13311
rect 40785 13277 40819 13311
rect 41061 13277 41095 13311
rect 42349 13277 42383 13311
rect 4077 13209 4111 13243
rect 10609 13209 10643 13243
rect 11805 13209 11839 13243
rect 14565 13209 14599 13243
rect 21557 13209 21591 13243
rect 23581 13209 23615 13243
rect 27721 13209 27755 13243
rect 38025 13209 38059 13243
rect 38552 13209 38586 13243
rect 5549 13141 5583 13175
rect 8033 13141 8067 13175
rect 8125 13141 8159 13175
rect 8493 13141 8527 13175
rect 8585 13141 8619 13175
rect 10333 13141 10367 13175
rect 21189 13141 21223 13175
rect 22017 13141 22051 13175
rect 22385 13141 22419 13175
rect 23949 13141 23983 13175
rect 29193 13141 29227 13175
rect 29561 13141 29595 13175
rect 30849 13141 30883 13175
rect 33977 13141 34011 13175
rect 36553 13141 36587 13175
rect 38669 13141 38703 13175
rect 38761 13141 38795 13175
rect 39497 13141 39531 13175
rect 4031 12937 4065 12971
rect 6377 12937 6411 12971
rect 10517 12937 10551 12971
rect 11621 12937 11655 12971
rect 15669 12937 15703 12971
rect 16221 12937 16255 12971
rect 19993 12937 20027 12971
rect 23857 12937 23891 12971
rect 24409 12937 24443 12971
rect 25513 12937 25547 12971
rect 26985 12937 27019 12971
rect 30849 12937 30883 12971
rect 32597 12937 32631 12971
rect 35081 12937 35115 12971
rect 39037 12937 39071 12971
rect 39773 12937 39807 12971
rect 10149 12869 10183 12903
rect 10365 12869 10399 12903
rect 17785 12869 17819 12903
rect 19165 12869 19199 12903
rect 25973 12869 26007 12903
rect 32689 12869 32723 12903
rect 35357 12869 35391 12903
rect 39129 12869 39163 12903
rect 5457 12801 5491 12835
rect 5825 12801 5859 12835
rect 6929 12801 6963 12835
rect 7389 12801 7423 12835
rect 7941 12801 7975 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11069 12801 11103 12835
rect 11161 12801 11195 12835
rect 11621 12801 11655 12835
rect 11989 12801 12023 12835
rect 14749 12801 14783 12835
rect 14841 12801 14875 12835
rect 15025 12801 15059 12835
rect 15393 12801 15427 12835
rect 15853 12801 15887 12835
rect 16037 12801 16071 12835
rect 16957 12801 16991 12835
rect 17233 12801 17267 12835
rect 17509 12801 17543 12835
rect 17969 12801 18003 12835
rect 18061 12801 18095 12835
rect 18153 12801 18187 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 18613 12801 18647 12835
rect 18981 12801 19015 12835
rect 19625 12801 19659 12835
rect 22017 12801 22051 12835
rect 22109 12801 22143 12835
rect 22293 12801 22327 12835
rect 22385 12801 22419 12835
rect 22477 12801 22511 12835
rect 22661 12801 22695 12835
rect 23567 12801 23601 12835
rect 24317 12801 24351 12835
rect 25881 12801 25915 12835
rect 26433 12801 26467 12835
rect 26617 12801 26651 12835
rect 27261 12801 27295 12835
rect 27629 12801 27663 12835
rect 28825 12801 28859 12835
rect 29193 12801 29227 12835
rect 29653 12801 29687 12835
rect 30481 12801 30515 12835
rect 31033 12801 31067 12835
rect 31125 12801 31159 12835
rect 31309 12801 31343 12835
rect 31401 12801 31435 12835
rect 32137 12801 32171 12835
rect 32413 12801 32447 12835
rect 32965 12801 32999 12835
rect 34989 12801 35023 12835
rect 35173 12801 35207 12835
rect 35817 12801 35851 12835
rect 35998 12801 36032 12835
rect 36093 12801 36127 12835
rect 37289 12801 37323 12835
rect 39313 12801 39347 12835
rect 39589 12801 39623 12835
rect 7297 12733 7331 12767
rect 7757 12733 7791 12767
rect 8309 12733 8343 12767
rect 9735 12733 9769 12767
rect 11253 12733 11287 12767
rect 11713 12733 11747 12767
rect 13001 12733 13035 12767
rect 15669 12733 15703 12767
rect 16681 12733 16715 12767
rect 18705 12733 18739 12767
rect 19349 12733 19383 12767
rect 19533 12733 19567 12767
rect 23489 12733 23523 12767
rect 24593 12733 24627 12767
rect 26065 12733 26099 12767
rect 26985 12733 27019 12767
rect 27353 12733 27387 12767
rect 28641 12733 28675 12767
rect 32229 12733 32263 12767
rect 32873 12733 32907 12767
rect 37565 12733 37599 12767
rect 39497 12733 39531 12767
rect 10609 12665 10643 12699
rect 17693 12665 17727 12699
rect 18797 12665 18831 12699
rect 21833 12665 21867 12699
rect 26801 12665 26835 12699
rect 35633 12665 35667 12699
rect 10333 12597 10367 12631
rect 11897 12597 11931 12631
rect 15025 12597 15059 12631
rect 15485 12597 15519 12631
rect 16773 12597 16807 12631
rect 17141 12597 17175 12631
rect 17325 12597 17359 12631
rect 17785 12597 17819 12631
rect 22661 12597 22695 12631
rect 23949 12597 23983 12631
rect 26433 12597 26467 12631
rect 27169 12597 27203 12631
rect 27445 12597 27479 12631
rect 27537 12597 27571 12631
rect 29009 12597 29043 12631
rect 30297 12597 30331 12631
rect 32137 12597 32171 12631
rect 32689 12597 32723 12631
rect 33149 12597 33183 12631
rect 10241 12393 10275 12427
rect 10885 12393 10919 12427
rect 11989 12393 12023 12427
rect 14105 12393 14139 12427
rect 14933 12393 14967 12427
rect 15761 12393 15795 12427
rect 17141 12393 17175 12427
rect 19257 12393 19291 12427
rect 19993 12393 20027 12427
rect 25881 12393 25915 12427
rect 29193 12393 29227 12427
rect 15209 12325 15243 12359
rect 19809 12325 19843 12359
rect 22201 12325 22235 12359
rect 24409 12325 24443 12359
rect 11805 12257 11839 12291
rect 22293 12257 22327 12291
rect 25053 12257 25087 12291
rect 26433 12257 26467 12291
rect 27169 12257 27203 12291
rect 27353 12257 27387 12291
rect 27905 12257 27939 12291
rect 27997 12257 28031 12291
rect 35449 12257 35483 12291
rect 10977 12189 11011 12223
rect 11345 12189 11379 12223
rect 11713 12189 11747 12223
rect 14289 12189 14323 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 16865 12189 16899 12223
rect 17141 12189 17175 12223
rect 19533 12189 19567 12223
rect 19901 12189 19935 12223
rect 20085 12189 20119 12223
rect 22017 12189 22051 12223
rect 26341 12189 26375 12223
rect 28181 12189 28215 12223
rect 28273 12189 28307 12223
rect 29193 12189 29227 12223
rect 29377 12189 29411 12223
rect 34897 12189 34931 12223
rect 35081 12189 35115 12223
rect 7205 12121 7239 12155
rect 9965 12121 9999 12155
rect 11437 12121 11471 12155
rect 26249 12121 26283 12155
rect 27537 12121 27571 12155
rect 27721 12121 27755 12155
rect 27997 12121 28031 12155
rect 37933 12121 37967 12155
rect 5733 12053 5767 12087
rect 11621 12053 11655 12087
rect 16957 12053 16991 12087
rect 19441 12053 19475 12087
rect 19625 12053 19659 12087
rect 21833 12053 21867 12087
rect 24777 12053 24811 12087
rect 24869 12053 24903 12087
rect 26709 12053 26743 12087
rect 27077 12053 27111 12087
rect 34989 12053 35023 12087
rect 36093 12053 36127 12087
rect 39221 12053 39255 12087
rect 9965 11849 9999 11883
rect 10701 11849 10735 11883
rect 11713 11849 11747 11883
rect 11897 11849 11931 11883
rect 13001 11849 13035 11883
rect 17325 11849 17359 11883
rect 17969 11849 18003 11883
rect 22109 11849 22143 11883
rect 24501 11849 24535 11883
rect 34437 11849 34471 11883
rect 34605 11849 34639 11883
rect 35633 11849 35667 11883
rect 37841 11849 37875 11883
rect 34805 11781 34839 11815
rect 9689 11713 9723 11747
rect 10333 11713 10367 11747
rect 10880 11713 10914 11747
rect 10977 11713 11011 11747
rect 11069 11713 11103 11747
rect 11252 11713 11286 11747
rect 11345 11713 11379 11747
rect 11529 11713 11563 11747
rect 12357 11713 12391 11747
rect 12909 11713 12943 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 15853 11713 15887 11747
rect 16037 11713 16071 11747
rect 16129 11713 16163 11747
rect 16681 11713 16715 11747
rect 16865 11713 16899 11747
rect 16957 11713 16991 11747
rect 17049 11713 17083 11747
rect 18153 11713 18187 11747
rect 18337 11713 18371 11747
rect 18429 11713 18463 11747
rect 22385 11713 22419 11747
rect 22477 11713 22511 11747
rect 22569 11713 22603 11747
rect 22753 11713 22787 11747
rect 23213 11713 23247 11747
rect 23397 11713 23431 11747
rect 23581 11713 23615 11747
rect 24685 11713 24719 11747
rect 24961 11713 24995 11747
rect 27353 11713 27387 11747
rect 31769 11713 31803 11747
rect 35449 11713 35483 11747
rect 37933 11713 37967 11747
rect 38853 11713 38887 11747
rect 7573 11645 7607 11679
rect 7849 11645 7883 11679
rect 9321 11645 9355 11679
rect 10609 11645 10643 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 12265 11645 12299 11679
rect 13461 11645 13495 11679
rect 13645 11645 13679 11679
rect 14381 11645 14415 11679
rect 14519 11645 14553 11679
rect 14657 11645 14691 11679
rect 23489 11645 23523 11679
rect 27445 11645 27479 11679
rect 27537 11645 27571 11679
rect 36185 11645 36219 11679
rect 38393 11645 38427 11679
rect 10517 11577 10551 11611
rect 14105 11577 14139 11611
rect 15853 11577 15887 11611
rect 24869 11577 24903 11611
rect 26985 11577 27019 11611
rect 10425 11509 10459 11543
rect 15301 11509 15335 11543
rect 22937 11509 22971 11543
rect 31677 11509 31711 11543
rect 34621 11509 34655 11543
rect 34897 11509 34931 11543
rect 38761 11509 38795 11543
rect 7573 11305 7607 11339
rect 10609 11305 10643 11339
rect 10793 11305 10827 11339
rect 11805 11305 11839 11339
rect 12081 11305 12115 11339
rect 13185 11305 13219 11339
rect 14565 11305 14599 11339
rect 14933 11305 14967 11339
rect 18521 11305 18555 11339
rect 18705 11305 18739 11339
rect 22201 11305 22235 11339
rect 24961 11305 24995 11339
rect 27997 11305 28031 11339
rect 29561 11305 29595 11339
rect 34970 11305 35004 11339
rect 36461 11305 36495 11339
rect 38945 11305 38979 11339
rect 12449 11237 12483 11271
rect 31769 11237 31803 11271
rect 32781 11237 32815 11271
rect 42533 11237 42567 11271
rect 7665 11169 7699 11203
rect 7849 11169 7883 11203
rect 9873 11169 9907 11203
rect 11713 11169 11747 11203
rect 12265 11169 12299 11203
rect 13185 11169 13219 11203
rect 13277 11169 13311 11203
rect 15117 11169 15151 11203
rect 15283 11169 15317 11203
rect 15393 11169 15427 11203
rect 18613 11169 18647 11203
rect 22937 11169 22971 11203
rect 31309 11169 31343 11203
rect 32597 11169 32631 11203
rect 33149 11169 33183 11203
rect 33977 11169 34011 11203
rect 34437 11169 34471 11203
rect 34713 11169 34747 11203
rect 37105 11169 37139 11203
rect 38025 11169 38059 11203
rect 38761 11169 38795 11203
rect 44005 11169 44039 11203
rect 7389 11101 7423 11135
rect 7481 11101 7515 11135
rect 7757 11101 7791 11135
rect 7941 11101 7975 11135
rect 9781 11101 9815 11135
rect 10425 11101 10459 11135
rect 10609 11101 10643 11135
rect 10885 11101 10919 11135
rect 11161 11101 11195 11135
rect 11621 11101 11655 11135
rect 12173 11101 12207 11135
rect 12541 11101 12575 11135
rect 13369 11101 13403 11135
rect 14095 11101 14129 11135
rect 14381 11101 14415 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 15198 11101 15232 11135
rect 17877 11101 17911 11135
rect 17969 11101 18003 11135
rect 18245 11101 18279 11135
rect 18337 11101 18371 11135
rect 18889 11101 18923 11135
rect 19533 11101 19567 11135
rect 19717 11101 19751 11135
rect 21649 11101 21683 11135
rect 21833 11101 21867 11135
rect 22017 11101 22051 11135
rect 22293 11101 22327 11135
rect 22661 11101 22695 11135
rect 22845 11101 22879 11135
rect 23029 11101 23063 11135
rect 24869 11101 24903 11135
rect 25053 11101 25087 11135
rect 27905 11101 27939 11135
rect 28089 11101 28123 11135
rect 29745 11101 29779 11135
rect 29837 11101 29871 11135
rect 31125 11101 31159 11135
rect 31585 11101 31619 11135
rect 31677 11101 31711 11135
rect 31861 11101 31895 11135
rect 32137 11101 32171 11135
rect 34345 11101 34379 11135
rect 38117 11101 38151 11135
rect 38393 11101 38427 11135
rect 38577 11101 38611 11135
rect 39497 11101 39531 11135
rect 44281 11101 44315 11135
rect 13001 11033 13035 11067
rect 14197 11033 14231 11067
rect 14749 11033 14783 11067
rect 18153 11033 18187 11067
rect 21925 11033 21959 11067
rect 31401 11033 31435 11067
rect 10977 10965 11011 10999
rect 11989 10965 12023 10999
rect 19073 10965 19107 10999
rect 19625 10965 19659 10999
rect 30941 10965 30975 10999
rect 32137 10965 32171 10999
rect 32689 10965 32723 10999
rect 36553 10965 36587 10999
rect 37381 10965 37415 10999
rect 6101 10761 6135 10795
rect 6929 10761 6963 10795
rect 12265 10761 12299 10795
rect 12725 10761 12759 10795
rect 15485 10761 15519 10795
rect 17141 10761 17175 10795
rect 17509 10761 17543 10795
rect 18613 10761 18647 10795
rect 19441 10761 19475 10795
rect 20177 10761 20211 10795
rect 22385 10761 22419 10795
rect 22575 10761 22609 10795
rect 24133 10761 24167 10795
rect 25145 10761 25179 10795
rect 25605 10761 25639 10795
rect 26065 10761 26099 10795
rect 26433 10761 26467 10795
rect 27905 10761 27939 10795
rect 29653 10761 29687 10795
rect 30297 10761 30331 10795
rect 35265 10761 35299 10795
rect 35449 10761 35483 10795
rect 37105 10761 37139 10795
rect 39037 10761 39071 10795
rect 19257 10693 19291 10727
rect 21557 10693 21591 10727
rect 22017 10693 22051 10727
rect 26525 10693 26559 10727
rect 27445 10693 27479 10727
rect 28089 10693 28123 10727
rect 28825 10693 28859 10727
rect 29285 10693 29319 10727
rect 29469 10693 29503 10727
rect 30573 10693 30607 10727
rect 30665 10693 30699 10727
rect 33793 10693 33827 10727
rect 35633 10693 35667 10727
rect 37565 10693 37599 10727
rect 6561 10625 6595 10659
rect 7205 10625 7239 10659
rect 8033 10625 8067 10659
rect 11621 10625 11655 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12081 10625 12115 10659
rect 12357 10625 12391 10659
rect 12541 10625 12575 10659
rect 15393 10625 15427 10659
rect 15577 10625 15611 10659
rect 17325 10625 17359 10659
rect 17417 10625 17451 10659
rect 18061 10625 18095 10659
rect 18429 10625 18463 10659
rect 19533 10625 19567 10659
rect 19625 10625 19659 10659
rect 19901 10625 19935 10659
rect 20361 10625 20395 10659
rect 20821 10625 20855 10659
rect 21465 10625 21499 10659
rect 21649 10625 21683 10659
rect 22201 10625 22235 10659
rect 22477 10625 22511 10659
rect 22661 10625 22695 10659
rect 22753 10625 22787 10659
rect 23949 10625 23983 10659
rect 24133 10625 24167 10659
rect 24685 10625 24719 10659
rect 25513 10625 25547 10659
rect 27353 10625 27387 10659
rect 27813 10625 27847 10659
rect 28365 10625 28399 10659
rect 28733 10625 28767 10659
rect 28917 10625 28951 10659
rect 29837 10625 29871 10659
rect 30481 10625 30515 10659
rect 30849 10625 30883 10659
rect 30941 10625 30975 10659
rect 31217 10625 31251 10659
rect 31585 10625 31619 10659
rect 31677 10625 31711 10659
rect 31953 10625 31987 10659
rect 32137 10625 32171 10659
rect 32321 10625 32355 10659
rect 32505 10625 32539 10659
rect 32689 10625 32723 10659
rect 35357 10625 35391 10659
rect 36829 10625 36863 10659
rect 37289 10625 37323 10659
rect 4353 10557 4387 10591
rect 4629 10557 4663 10591
rect 6653 10557 6687 10591
rect 7297 10557 7331 10591
rect 7941 10557 7975 10591
rect 17693 10557 17727 10591
rect 17785 10557 17819 10591
rect 20545 10557 20579 10591
rect 20637 10557 20671 10591
rect 24777 10557 24811 10591
rect 24961 10557 24995 10591
rect 25697 10557 25731 10591
rect 26709 10557 26743 10591
rect 27537 10557 27571 10591
rect 28089 10557 28123 10591
rect 29101 10557 29135 10591
rect 29929 10557 29963 10591
rect 30021 10557 30055 10591
rect 30113 10557 30147 10591
rect 31033 10557 31067 10591
rect 31493 10557 31527 10591
rect 32413 10557 32447 10591
rect 33517 10557 33551 10591
rect 36737 10557 36771 10591
rect 36921 10557 36955 10591
rect 39129 10557 39163 10591
rect 39681 10557 39715 10591
rect 7573 10489 7607 10523
rect 19257 10489 19291 10523
rect 20085 10489 20119 10523
rect 20453 10489 20487 10523
rect 24317 10489 24351 10523
rect 26985 10489 27019 10523
rect 7757 10421 7791 10455
rect 18153 10421 18187 10455
rect 19717 10421 19751 10455
rect 28273 10421 28307 10455
rect 31401 10421 31435 10455
rect 32873 10421 32907 10455
rect 35633 10421 35667 10455
rect 4629 10217 4663 10251
rect 10977 10217 11011 10251
rect 19257 10217 19291 10251
rect 22017 10217 22051 10251
rect 28181 10217 28215 10251
rect 28457 10217 28491 10251
rect 28825 10217 28859 10251
rect 29561 10217 29595 10251
rect 31493 10217 31527 10251
rect 37657 10217 37691 10251
rect 10701 10149 10735 10183
rect 15669 10149 15703 10183
rect 18981 10149 19015 10183
rect 19809 10149 19843 10183
rect 9965 10081 9999 10115
rect 16129 10081 16163 10115
rect 16221 10081 16255 10115
rect 19073 10081 19107 10115
rect 39405 10081 39439 10115
rect 5181 10013 5215 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10333 10013 10367 10047
rect 10517 10013 10551 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 15577 10013 15611 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16037 10013 16071 10047
rect 18798 9991 18832 10025
rect 18889 10013 18923 10047
rect 19438 10013 19472 10047
rect 19901 10013 19935 10047
rect 22201 10013 22235 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 27905 10013 27939 10047
rect 28089 10013 28123 10047
rect 28641 10013 28675 10047
rect 28917 10013 28951 10047
rect 30021 10013 30055 10047
rect 30205 10013 30239 10047
rect 32965 10013 32999 10047
rect 9965 9945 9999 9979
rect 22385 9945 22419 9979
rect 28365 9945 28399 9979
rect 29745 9945 29779 9979
rect 29929 9945 29963 9979
rect 39129 9945 39163 9979
rect 10425 9877 10459 9911
rect 16405 9877 16439 9911
rect 19441 9877 19475 9911
rect 27721 9877 27755 9911
rect 30113 9877 30147 9911
rect 2697 9673 2731 9707
rect 4537 9673 4571 9707
rect 23213 9673 23247 9707
rect 23581 9673 23615 9707
rect 24317 9673 24351 9707
rect 24777 9673 24811 9707
rect 26249 9673 26283 9707
rect 40877 9673 40911 9707
rect 3065 9605 3099 9639
rect 14289 9605 14323 9639
rect 21833 9605 21867 9639
rect 42533 9605 42567 9639
rect 2513 9537 2547 9571
rect 10308 9537 10342 9571
rect 13369 9537 13403 9571
rect 13553 9537 13587 9571
rect 13829 9537 13863 9571
rect 14105 9537 14139 9571
rect 16129 9537 16163 9571
rect 16221 9537 16255 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 17325 9537 17359 9571
rect 22109 9537 22143 9571
rect 24685 9537 24719 9571
rect 26157 9537 26191 9571
rect 28641 9537 28675 9571
rect 28733 9537 28767 9571
rect 28917 9537 28951 9571
rect 29009 9537 29043 9571
rect 29193 9537 29227 9571
rect 29285 9537 29319 9571
rect 29469 9537 29503 9571
rect 30665 9537 30699 9571
rect 30849 9537 30883 9571
rect 31493 9537 31527 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 2789 9469 2823 9503
rect 10149 9469 10183 9503
rect 10425 9469 10459 9503
rect 11161 9469 11195 9503
rect 11345 9469 11379 9503
rect 13737 9469 13771 9503
rect 14013 9469 14047 9503
rect 16037 9469 16071 9503
rect 16313 9469 16347 9503
rect 21833 9469 21867 9503
rect 23673 9469 23707 9503
rect 23765 9469 23799 9503
rect 24961 9469 24995 9503
rect 26433 9469 26467 9503
rect 28549 9469 28583 9503
rect 31309 9469 31343 9503
rect 31677 9469 31711 9503
rect 31769 9469 31803 9503
rect 33701 9469 33735 9503
rect 41521 9469 41555 9503
rect 10701 9401 10735 9435
rect 13645 9401 13679 9435
rect 16681 9401 16715 9435
rect 28273 9401 28307 9435
rect 30757 9401 30791 9435
rect 33977 9401 34011 9435
rect 9505 9333 9539 9367
rect 14473 9333 14507 9367
rect 16497 9333 16531 9367
rect 22017 9333 22051 9367
rect 25789 9333 25823 9367
rect 28457 9333 28491 9367
rect 28733 9333 28767 9367
rect 29101 9333 29135 9367
rect 29561 9333 29595 9367
rect 32229 9333 32263 9367
rect 34161 9333 34195 9367
rect 43821 9333 43855 9367
rect 2237 9129 2271 9163
rect 9781 9129 9815 9163
rect 10701 9129 10735 9163
rect 11253 9129 11287 9163
rect 11529 9129 11563 9163
rect 12081 9129 12115 9163
rect 13921 9129 13955 9163
rect 14105 9129 14139 9163
rect 14657 9129 14691 9163
rect 16865 9129 16899 9163
rect 19901 9129 19935 9163
rect 22201 9129 22235 9163
rect 22753 9129 22787 9163
rect 24409 9129 24443 9163
rect 25697 9129 25731 9163
rect 30389 9129 30423 9163
rect 31493 9129 31527 9163
rect 33044 9129 33078 9163
rect 1593 9061 1627 9095
rect 2053 9061 2087 9095
rect 13369 9061 13403 9095
rect 16957 9061 16991 9095
rect 17969 9061 18003 9095
rect 18061 9061 18095 9095
rect 20453 9061 20487 9095
rect 26525 9061 26559 9095
rect 1777 8993 1811 9027
rect 6745 8993 6779 9027
rect 7021 8993 7055 9027
rect 7297 8993 7331 9027
rect 10793 8993 10827 9027
rect 12909 8993 12943 9027
rect 13553 8993 13587 9027
rect 16221 8993 16255 9027
rect 18981 8993 19015 9027
rect 20545 8993 20579 9027
rect 21557 8993 21591 9027
rect 22569 8993 22603 9027
rect 24869 8993 24903 9027
rect 25053 8993 25087 9027
rect 26341 8993 26375 9027
rect 26985 8993 27019 9027
rect 27169 8993 27203 9027
rect 31125 8993 31159 9027
rect 32781 8993 32815 9027
rect 35081 8993 35115 9027
rect 1409 8925 1443 8959
rect 6653 8925 6687 8959
rect 7481 8925 7515 8959
rect 8125 8925 8159 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10885 8925 10919 8959
rect 11069 8925 11103 8959
rect 11529 8925 11563 8959
rect 11707 8925 11741 8959
rect 11989 8925 12023 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 13461 8925 13495 8959
rect 13737 8925 13771 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 14657 8925 14691 8959
rect 14749 8925 14783 8959
rect 15945 8925 15979 8959
rect 16129 8925 16163 8959
rect 16313 8925 16347 8959
rect 16740 8925 16774 8959
rect 17141 8925 17175 8959
rect 17233 8925 17267 8959
rect 17417 8925 17451 8959
rect 17509 8925 17543 8959
rect 17693 8925 17727 8959
rect 17969 8925 18003 8959
rect 18337 8925 18371 8959
rect 18429 8925 18463 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 18797 8925 18831 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 19533 8925 19567 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 21741 8925 21775 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 22109 8925 22143 8959
rect 22385 8925 22419 8959
rect 22661 8925 22695 8959
rect 22845 8925 22879 8959
rect 26157 8925 26191 8959
rect 27629 8925 27663 8959
rect 27813 8925 27847 8959
rect 27905 8925 27939 8959
rect 30113 8925 30147 8959
rect 30297 8925 30331 8959
rect 30573 8925 30607 8959
rect 30941 8925 30975 8959
rect 31033 8919 31067 8953
rect 31585 8925 31619 8959
rect 36921 8925 36955 8959
rect 37565 8925 37599 8959
rect 37657 8925 37691 8959
rect 37841 8925 37875 8959
rect 7389 8857 7423 8891
rect 9781 8857 9815 8891
rect 10333 8857 10367 8891
rect 10517 8857 10551 8891
rect 18061 8857 18095 8891
rect 24777 8857 24811 8891
rect 28181 8857 28215 8891
rect 30205 8857 30239 8891
rect 30665 8857 30699 8891
rect 30757 8857 30791 8891
rect 35357 8857 35391 8891
rect 7849 8789 7883 8823
rect 7941 8789 7975 8823
rect 11345 8789 11379 8823
rect 15025 8789 15059 8823
rect 16037 8789 16071 8823
rect 16681 8789 16715 8823
rect 17785 8789 17819 8823
rect 18245 8789 18279 8823
rect 26065 8789 26099 8823
rect 26893 8789 26927 8823
rect 27997 8789 28031 8823
rect 34529 8789 34563 8823
rect 36829 8789 36863 8823
rect 37749 8789 37783 8823
rect 10425 8585 10459 8619
rect 10701 8585 10735 8619
rect 13093 8585 13127 8619
rect 13461 8585 13495 8619
rect 14381 8585 14415 8619
rect 17325 8585 17359 8619
rect 20177 8585 20211 8619
rect 21373 8585 21407 8619
rect 23305 8585 23339 8619
rect 24041 8585 24075 8619
rect 24409 8585 24443 8619
rect 26065 8585 26099 8619
rect 27353 8585 27387 8619
rect 29009 8585 29043 8619
rect 30389 8585 30423 8619
rect 35541 8585 35575 8619
rect 42533 8585 42567 8619
rect 34437 8517 34471 8551
rect 7849 8449 7883 8483
rect 9275 8449 9309 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 13277 8449 13311 8483
rect 13553 8449 13587 8483
rect 14105 8449 14139 8483
rect 14289 8449 14323 8483
rect 14381 8449 14415 8483
rect 17233 8449 17267 8483
rect 17417 8449 17451 8483
rect 19533 8449 19567 8483
rect 21649 8449 21683 8483
rect 21925 8449 21959 8483
rect 22109 8449 22143 8483
rect 23581 8449 23615 8483
rect 23673 8449 23707 8483
rect 23765 8449 23799 8483
rect 23949 8449 23983 8483
rect 24501 8449 24535 8483
rect 27537 8449 27571 8483
rect 28549 8449 28583 8483
rect 28825 8449 28859 8483
rect 29101 8449 29135 8483
rect 30297 8449 30331 8483
rect 30481 8449 30515 8483
rect 30757 8449 30791 8483
rect 31033 8449 31067 8483
rect 31493 8449 31527 8483
rect 31780 8449 31814 8483
rect 32137 8449 32171 8483
rect 32321 8449 32355 8483
rect 33885 8449 33919 8483
rect 34713 8449 34747 8483
rect 35449 8449 35483 8483
rect 35633 8449 35667 8483
rect 35909 8449 35943 8483
rect 36093 8449 36127 8483
rect 36921 8449 36955 8483
rect 37105 8449 37139 8483
rect 37289 8449 37323 8483
rect 38025 8449 38059 8483
rect 38209 8449 38243 8483
rect 38301 8449 38335 8483
rect 44281 8449 44315 8483
rect 7481 8381 7515 8415
rect 12173 8381 12207 8415
rect 12357 8381 12391 8415
rect 18337 8381 18371 8415
rect 18521 8381 18555 8415
rect 19257 8381 19291 8415
rect 19395 8381 19429 8415
rect 21373 8381 21407 8415
rect 24593 8381 24627 8415
rect 26157 8381 26191 8415
rect 26249 8381 26283 8415
rect 27721 8381 27755 8415
rect 30849 8381 30883 8415
rect 30941 8381 30975 8415
rect 33977 8381 34011 8415
rect 35725 8381 35759 8415
rect 36829 8381 36863 8415
rect 37013 8381 37047 8415
rect 37933 8381 37967 8415
rect 44005 8381 44039 8415
rect 18981 8313 19015 8347
rect 21557 8313 21591 8347
rect 28273 8313 28307 8347
rect 30573 8313 30607 8347
rect 31217 8313 31251 8347
rect 32229 8313 32263 8347
rect 33701 8313 33735 8347
rect 34069 8313 34103 8347
rect 34529 8313 34563 8347
rect 38025 8313 38059 8347
rect 11897 8245 11931 8279
rect 22109 8245 22143 8279
rect 25697 8245 25731 8279
rect 28733 8245 28767 8279
rect 31585 8245 31619 8279
rect 36185 8245 36219 8279
rect 11161 8041 11195 8075
rect 13369 8041 13403 8075
rect 15577 8041 15611 8075
rect 16313 8041 16347 8075
rect 17785 8041 17819 8075
rect 18613 8041 18647 8075
rect 19257 8041 19291 8075
rect 21465 8041 21499 8075
rect 22293 8041 22327 8075
rect 23489 8041 23523 8075
rect 25881 8041 25915 8075
rect 28089 8041 28123 8075
rect 28273 8041 28307 8075
rect 31125 8041 31159 8075
rect 31585 8041 31619 8075
rect 38117 8041 38151 8075
rect 38393 8041 38427 8075
rect 43545 8041 43579 8075
rect 10793 7973 10827 8007
rect 19073 7973 19107 8007
rect 30205 7973 30239 8007
rect 38209 7973 38243 8007
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 11989 7905 12023 7939
rect 12725 7905 12759 7939
rect 16037 7905 16071 7939
rect 16865 7905 16899 7939
rect 18521 7905 18555 7939
rect 19901 7905 19935 7939
rect 21925 7905 21959 7939
rect 22845 7905 22879 7939
rect 24133 7905 24167 7939
rect 24961 7905 24995 7939
rect 26525 7905 26559 7939
rect 29561 7905 29595 7939
rect 31217 7905 31251 7939
rect 31677 7905 31711 7939
rect 6745 7837 6779 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 10517 7837 10551 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 11562 7837 11596 7871
rect 12081 7837 12115 7871
rect 12633 7837 12667 7871
rect 12817 7837 12851 7871
rect 15117 7837 15151 7871
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 15669 7837 15703 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16681 7837 16715 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17969 7837 18003 7871
rect 18061 7837 18095 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 19073 7837 19107 7871
rect 19625 7837 19659 7871
rect 19717 7837 19751 7871
rect 21649 7837 21683 7871
rect 21741 7837 21775 7871
rect 22017 7837 22051 7871
rect 23857 7837 23891 7871
rect 24777 7837 24811 7871
rect 26341 7837 26375 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 31309 7837 31343 7871
rect 31769 7847 31803 7881
rect 34529 7837 34563 7871
rect 37473 7837 37507 7871
rect 43361 7837 43395 7871
rect 13093 7769 13127 7803
rect 15761 7769 15795 7803
rect 17785 7769 17819 7803
rect 22661 7769 22695 7803
rect 24869 7769 24903 7803
rect 26249 7769 26283 7803
rect 28457 7769 28491 7803
rect 34253 7769 34287 7803
rect 37105 7769 37139 7803
rect 38361 7769 38395 7803
rect 38577 7769 38611 7803
rect 9965 7701 9999 7735
rect 11437 7701 11471 7735
rect 11621 7701 11655 7735
rect 15853 7701 15887 7735
rect 16497 7701 16531 7735
rect 17049 7701 17083 7735
rect 22753 7701 22787 7735
rect 23949 7701 23983 7735
rect 24409 7701 24443 7735
rect 28257 7701 28291 7735
rect 30941 7701 30975 7735
rect 31401 7701 31435 7735
rect 32781 7701 32815 7735
rect 35817 7701 35851 7735
rect 7297 7497 7331 7531
rect 10977 7497 11011 7531
rect 11161 7497 11195 7531
rect 12357 7497 12391 7531
rect 12725 7497 12759 7531
rect 19073 7497 19107 7531
rect 21373 7497 21407 7531
rect 22569 7497 22603 7531
rect 23949 7497 23983 7531
rect 25329 7497 25363 7531
rect 25789 7497 25823 7531
rect 27445 7497 27479 7531
rect 28089 7497 28123 7531
rect 29653 7497 29687 7531
rect 33149 7497 33183 7531
rect 37105 7497 37139 7531
rect 37473 7497 37507 7531
rect 43361 7497 43395 7531
rect 7389 7429 7423 7463
rect 15577 7429 15611 7463
rect 16037 7429 16071 7463
rect 22385 7429 22419 7463
rect 24409 7429 24443 7463
rect 26249 7429 26283 7463
rect 28625 7429 28659 7463
rect 28825 7429 28859 7463
rect 31217 7429 31251 7463
rect 31401 7429 31435 7463
rect 34621 7429 34655 7463
rect 43821 7429 43855 7463
rect 5825 7361 5859 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11069 7361 11103 7395
rect 11253 7361 11287 7395
rect 15393 7361 15427 7395
rect 15669 7361 15703 7395
rect 15945 7361 15979 7395
rect 18613 7361 18647 7395
rect 18705 7361 18739 7395
rect 18889 7361 18923 7395
rect 21005 7361 21039 7395
rect 21189 7361 21223 7395
rect 22844 7361 22878 7395
rect 24317 7361 24351 7395
rect 24869 7361 24903 7395
rect 25697 7361 25731 7395
rect 26433 7361 26467 7395
rect 26525 7361 26559 7395
rect 26709 7361 26743 7395
rect 26801 7361 26835 7395
rect 27353 7361 27387 7395
rect 27813 7361 27847 7395
rect 28181 7361 28215 7395
rect 28905 7361 28939 7395
rect 29101 7361 29135 7395
rect 29193 7361 29227 7395
rect 29331 7361 29365 7395
rect 29930 7361 29964 7395
rect 30113 7361 30147 7395
rect 30941 7361 30975 7395
rect 39221 7361 39255 7395
rect 44281 7361 44315 7395
rect 5917 7293 5951 7327
rect 7481 7293 7515 7327
rect 10701 7293 10735 7327
rect 10793 7293 10827 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 15209 7293 15243 7327
rect 22569 7293 22603 7327
rect 24593 7293 24627 7327
rect 25881 7293 25915 7327
rect 27537 7293 27571 7327
rect 27997 7293 28031 7327
rect 29837 7293 29871 7327
rect 30021 7293 30055 7327
rect 30849 7293 30883 7327
rect 35357 7293 35391 7327
rect 35633 7293 35667 7327
rect 38945 7293 38979 7327
rect 6193 7225 6227 7259
rect 22201 7225 22235 7259
rect 27813 7225 27847 7259
rect 29561 7225 29595 7259
rect 43545 7225 43579 7259
rect 44097 7225 44131 7259
rect 6929 7157 6963 7191
rect 22753 7157 22787 7191
rect 25145 7157 25179 7191
rect 26985 7157 27019 7191
rect 28457 7157 28491 7191
rect 28641 7157 28675 7191
rect 30573 7157 30607 7191
rect 30757 7157 30791 7191
rect 31033 7157 31067 7191
rect 10977 6953 11011 6987
rect 11437 6953 11471 6987
rect 14749 6953 14783 6987
rect 14933 6953 14967 6987
rect 18061 6953 18095 6987
rect 25053 6953 25087 6987
rect 29561 6953 29595 6987
rect 29745 6953 29779 6987
rect 31585 6953 31619 6987
rect 2237 6885 2271 6919
rect 7021 6885 7055 6919
rect 18153 6885 18187 6919
rect 30849 6885 30883 6919
rect 33793 6885 33827 6919
rect 1961 6817 1995 6851
rect 2421 6817 2455 6851
rect 7573 6817 7607 6851
rect 8401 6817 8435 6851
rect 11345 6817 11379 6851
rect 25605 6817 25639 6851
rect 26525 6817 26559 6851
rect 26684 6817 26718 6851
rect 26801 6817 26835 6851
rect 27077 6817 27111 6851
rect 27537 6817 27571 6851
rect 28181 6817 28215 6851
rect 30481 6817 30515 6851
rect 33425 6817 33459 6851
rect 33885 6817 33919 6851
rect 34805 6817 34839 6851
rect 36553 6817 36587 6851
rect 37473 6817 37507 6851
rect 38025 6817 38059 6851
rect 2973 6749 3007 6783
rect 6745 6749 6779 6783
rect 7389 6749 7423 6783
rect 8217 6749 8251 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 11437 6749 11471 6783
rect 11621 6749 11655 6783
rect 11805 6749 11839 6783
rect 11989 6749 12023 6783
rect 12725 6749 12759 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 16129 6749 16163 6783
rect 16313 6749 16347 6783
rect 17785 6749 17819 6783
rect 18061 6749 18095 6783
rect 18429 6749 18463 6783
rect 25881 6749 25915 6783
rect 27721 6749 27755 6783
rect 28089 6749 28123 6783
rect 28365 6749 28399 6783
rect 28641 6749 28675 6783
rect 28917 6749 28951 6783
rect 29009 6749 29043 6783
rect 30113 6749 30147 6783
rect 30665 6749 30699 6783
rect 31033 6749 31067 6783
rect 31217 6749 31251 6783
rect 31401 6749 31435 6783
rect 31493 6749 31527 6783
rect 31677 6749 31711 6783
rect 33333 6749 33367 6783
rect 37289 6749 37323 6783
rect 7481 6681 7515 6715
rect 8309 6681 8343 6715
rect 12173 6681 12207 6715
rect 13369 6681 13403 6715
rect 13737 6681 13771 6715
rect 18153 6681 18187 6715
rect 18337 6681 18371 6715
rect 25421 6681 25455 6715
rect 29929 6681 29963 6715
rect 30297 6681 30331 6715
rect 35081 6681 35115 6715
rect 3157 6613 3191 6647
rect 6929 6613 6963 6647
rect 7849 6613 7883 6647
rect 12909 6613 12943 6647
rect 14105 6613 14139 6647
rect 16221 6613 16255 6647
rect 17877 6613 17911 6647
rect 25513 6613 25547 6647
rect 29719 6613 29753 6647
rect 31309 6613 31343 6647
rect 33149 6613 33183 6647
rect 37105 6613 37139 6647
rect 5273 6409 5307 6443
rect 14933 6409 14967 6443
rect 15117 6409 15151 6443
rect 16313 6409 16347 6443
rect 16865 6409 16899 6443
rect 20177 6409 20211 6443
rect 22477 6409 22511 6443
rect 35725 6409 35759 6443
rect 3801 6341 3835 6375
rect 10517 6341 10551 6375
rect 13921 6341 13955 6375
rect 14298 6341 14332 6375
rect 17509 6341 17543 6375
rect 27445 6341 27479 6375
rect 9413 6273 9447 6307
rect 10333 6273 10367 6307
rect 10977 6273 11011 6307
rect 11713 6273 11747 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 14841 6273 14875 6307
rect 15025 6273 15059 6307
rect 15393 6273 15427 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 16681 6273 16715 6307
rect 16865 6273 16899 6307
rect 17060 6273 17094 6307
rect 17325 6273 17359 6307
rect 17601 6273 17635 6307
rect 17785 6273 17819 6307
rect 17877 6273 17911 6307
rect 18061 6273 18095 6307
rect 18337 6273 18371 6307
rect 19257 6273 19291 6307
rect 22385 6273 22419 6307
rect 22477 6273 22511 6307
rect 22661 6273 22695 6307
rect 27077 6273 27111 6307
rect 28824 6273 28858 6307
rect 28917 6273 28951 6307
rect 29009 6273 29043 6307
rect 29193 6273 29227 6307
rect 35817 6273 35851 6307
rect 37473 6273 37507 6307
rect 3525 6205 3559 6239
rect 7389 6205 7423 6239
rect 7665 6205 7699 6239
rect 10149 6205 10183 6239
rect 10701 6205 10735 6239
rect 11805 6205 11839 6239
rect 12909 6205 12943 6239
rect 15301 6205 15335 6239
rect 15485 6205 15519 6239
rect 15577 6205 15611 6239
rect 17233 6205 17267 6239
rect 18521 6205 18555 6239
rect 19374 6205 19408 6239
rect 19533 6205 19567 6239
rect 22109 6205 22143 6239
rect 37381 6205 37415 6239
rect 37841 6205 37875 6239
rect 17141 6137 17175 6171
rect 17969 6137 18003 6171
rect 18245 6137 18279 6171
rect 18981 6137 19015 6171
rect 21833 6137 21867 6171
rect 28549 6137 28583 6171
rect 12725 6069 12759 6103
rect 13553 6069 13587 6103
rect 14289 6069 14323 6103
rect 14473 6069 14507 6103
rect 22293 6069 22327 6103
rect 12909 5865 12943 5899
rect 16221 5865 16255 5899
rect 16405 5865 16439 5899
rect 17877 5865 17911 5899
rect 18337 5865 18371 5899
rect 19717 5865 19751 5899
rect 21925 5865 21959 5899
rect 24225 5865 24259 5899
rect 32676 5865 32710 5899
rect 12541 5797 12575 5831
rect 15577 5797 15611 5831
rect 24593 5797 24627 5831
rect 13645 5729 13679 5763
rect 19257 5729 19291 5763
rect 20453 5729 20487 5763
rect 22109 5729 22143 5763
rect 25237 5729 25271 5763
rect 32413 5729 32447 5763
rect 6745 5661 6779 5695
rect 6837 5661 6871 5695
rect 12541 5661 12575 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 13829 5661 13863 5695
rect 13921 5661 13955 5695
rect 15485 5661 15519 5695
rect 15577 5661 15611 5695
rect 16313 5661 16347 5695
rect 16497 5661 16531 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 18153 5661 18187 5695
rect 19349 5661 19383 5695
rect 19533 5661 19567 5695
rect 20177 5661 20211 5695
rect 22293 5661 22327 5695
rect 22477 5661 22511 5695
rect 22569 5661 22603 5695
rect 23765 5661 23799 5695
rect 24041 5661 24075 5695
rect 24409 5661 24443 5695
rect 25145 5661 25179 5695
rect 13185 5593 13219 5627
rect 13415 5593 13449 5627
rect 15853 5593 15887 5627
rect 16037 5593 16071 5627
rect 23857 5593 23891 5627
rect 6561 5525 6595 5559
rect 8125 5525 8159 5559
rect 12725 5525 12759 5559
rect 13645 5525 13679 5559
rect 22753 5525 22787 5559
rect 34161 5525 34195 5559
rect 8171 5321 8205 5355
rect 10609 5321 10643 5355
rect 11069 5321 11103 5355
rect 12909 5321 12943 5355
rect 15025 5321 15059 5355
rect 31769 5321 31803 5355
rect 8677 5253 8711 5287
rect 9045 5253 9079 5287
rect 10057 5253 10091 5287
rect 13369 5253 13403 5287
rect 26157 5253 26191 5287
rect 32229 5253 32263 5287
rect 33149 5253 33183 5287
rect 6377 5185 6411 5219
rect 9505 5185 9539 5219
rect 9689 5185 9723 5219
rect 9965 5185 9999 5219
rect 10517 5185 10551 5219
rect 10793 5185 10827 5219
rect 11253 5185 11287 5219
rect 11713 5185 11747 5219
rect 11891 5185 11925 5219
rect 14749 5185 14783 5219
rect 14933 5185 14967 5219
rect 22385 5185 22419 5219
rect 22569 5185 22603 5219
rect 26249 5185 26283 5219
rect 26609 5185 26643 5219
rect 31033 5185 31067 5219
rect 31217 5185 31251 5219
rect 31309 5185 31343 5219
rect 31401 5185 31435 5219
rect 31585 5185 31619 5219
rect 32137 5185 32171 5219
rect 32873 5185 32907 5219
rect 6745 5117 6779 5151
rect 29009 5117 29043 5151
rect 11897 5049 11931 5083
rect 13001 5049 13035 5083
rect 25789 5049 25823 5083
rect 31033 5049 31067 5083
rect 9873 4981 9907 5015
rect 22569 4981 22603 5015
rect 26525 4981 26559 5015
rect 28365 4981 28399 5015
rect 34621 4981 34655 5015
rect 11069 4777 11103 4811
rect 11253 4777 11287 4811
rect 11713 4777 11747 4811
rect 13277 4777 13311 4811
rect 13737 4777 13771 4811
rect 15853 4777 15887 4811
rect 19257 4777 19291 4811
rect 22753 4777 22787 4811
rect 29377 4777 29411 4811
rect 30665 4777 30699 4811
rect 34805 4777 34839 4811
rect 10701 4709 10735 4743
rect 19533 4709 19567 4743
rect 33241 4709 33275 4743
rect 33425 4709 33459 4743
rect 12449 4641 12483 4675
rect 15025 4641 15059 4675
rect 15669 4641 15703 4675
rect 18889 4641 18923 4675
rect 19625 4641 19659 4675
rect 19717 4641 19751 4675
rect 27905 4641 27939 4675
rect 32413 4641 32447 4675
rect 7021 4573 7055 4607
rect 9873 4573 9907 4607
rect 10057 4573 10091 4607
rect 10609 4573 10643 4607
rect 12081 4573 12115 4607
rect 12357 4573 12391 4607
rect 12633 4573 12667 4607
rect 12817 4573 12851 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 15117 4573 15151 4607
rect 15485 4573 15519 4607
rect 15945 4573 15979 4607
rect 18797 4573 18831 4607
rect 18981 4573 19015 4607
rect 19441 4573 19475 4607
rect 19901 4573 19935 4607
rect 22385 4573 22419 4607
rect 23029 4573 23063 4607
rect 23213 4573 23247 4607
rect 23397 4573 23431 4607
rect 23673 4573 23707 4607
rect 23765 4573 23799 4607
rect 24409 4573 24443 4607
rect 26433 4573 26467 4607
rect 27629 4573 27663 4607
rect 33701 4573 33735 4607
rect 34437 4573 34471 4607
rect 34713 4573 34747 4607
rect 10885 4505 10919 4539
rect 11090 4505 11124 4539
rect 11437 4505 11471 4539
rect 15669 4505 15703 4539
rect 23581 4505 23615 4539
rect 24685 4505 24719 4539
rect 32137 4505 32171 4539
rect 33793 4505 33827 4539
rect 7205 4437 7239 4471
rect 22753 4437 22787 4471
rect 22937 4437 22971 4471
rect 23121 4437 23155 4471
rect 23949 4437 23983 4471
rect 35173 4437 35207 4471
rect 22477 4233 22511 4267
rect 35357 4233 35391 4267
rect 9321 4165 9355 4199
rect 10057 4165 10091 4199
rect 14749 4165 14783 4199
rect 15209 4165 15243 4199
rect 17785 4165 17819 4199
rect 21649 4165 21683 4199
rect 28733 4165 28767 4199
rect 7021 4097 7055 4131
rect 9137 4097 9171 4131
rect 9413 4097 9447 4131
rect 11253 4097 11287 4131
rect 11713 4097 11747 4131
rect 12081 4097 12115 4131
rect 14197 4097 14231 4131
rect 14933 4097 14967 4131
rect 15025 4097 15059 4131
rect 15669 4097 15703 4131
rect 16313 4097 16347 4131
rect 16497 4097 16531 4131
rect 16865 4097 16899 4131
rect 17141 4097 17175 4131
rect 17233 4097 17267 4131
rect 17509 4097 17543 4131
rect 17601 4097 17635 4131
rect 17877 4097 17911 4131
rect 18061 4097 18095 4131
rect 18245 4097 18279 4131
rect 18337 4097 18371 4131
rect 18429 4097 18463 4131
rect 19073 4097 19107 4131
rect 20085 4097 20119 4131
rect 22569 4097 22603 4131
rect 23489 4097 23523 4131
rect 23765 4097 23799 4131
rect 24133 4097 24167 4131
rect 24317 4097 24351 4131
rect 24593 4097 24627 4131
rect 24685 4097 24719 4131
rect 24869 4097 24903 4131
rect 37105 4097 37139 4131
rect 7389 4029 7423 4063
rect 8861 4029 8895 4063
rect 9873 4029 9907 4063
rect 10977 4029 11011 4063
rect 11529 4029 11563 4063
rect 12357 4029 12391 4063
rect 12541 4029 12575 4063
rect 13277 4029 13311 4063
rect 13415 4029 13449 4063
rect 13553 4029 13587 4063
rect 18521 4029 18555 4063
rect 18797 4029 18831 4063
rect 22385 4029 22419 4063
rect 23949 4029 23983 4063
rect 24409 4029 24443 4063
rect 24777 4029 24811 4063
rect 29193 4029 29227 4063
rect 29469 4029 29503 4063
rect 30941 4029 30975 4063
rect 36829 4029 36863 4063
rect 11989 3961 12023 3995
rect 13001 3961 13035 3995
rect 16313 3961 16347 3995
rect 17509 3961 17543 3995
rect 17969 3961 18003 3995
rect 18705 3961 18739 3995
rect 18981 3961 19015 3995
rect 23581 3961 23615 3995
rect 23673 3961 23707 3995
rect 24225 3961 24259 3995
rect 10333 3893 10367 3927
rect 14749 3893 14783 3927
rect 15485 3893 15519 3927
rect 15761 3893 15795 3927
rect 16957 3893 16991 3927
rect 17417 3893 17451 3927
rect 18889 3893 18923 3927
rect 22937 3893 22971 3927
rect 23305 3893 23339 3927
rect 27445 3893 27479 3927
rect 10333 3689 10367 3723
rect 13185 3689 13219 3723
rect 14841 3689 14875 3723
rect 15761 3689 15795 3723
rect 18705 3689 18739 3723
rect 22109 3689 22143 3723
rect 23949 3689 23983 3723
rect 26157 3689 26191 3723
rect 28733 3689 28767 3723
rect 36277 3689 36311 3723
rect 9597 3621 9631 3655
rect 11437 3621 11471 3655
rect 12265 3621 12299 3655
rect 13461 3621 13495 3655
rect 14657 3621 14691 3655
rect 16313 3621 16347 3655
rect 22753 3621 22787 3655
rect 23581 3621 23615 3655
rect 10701 3553 10735 3587
rect 12633 3553 12667 3587
rect 15209 3553 15243 3587
rect 15393 3553 15427 3587
rect 16129 3553 16163 3587
rect 16405 3553 16439 3587
rect 17049 3553 17083 3587
rect 17325 3553 17359 3587
rect 17463 3553 17497 3587
rect 20361 3553 20395 3587
rect 20729 3553 20763 3587
rect 22293 3553 22327 3587
rect 26985 3553 27019 3587
rect 9229 3485 9263 3519
rect 9781 3485 9815 3519
rect 10241 3485 10275 3519
rect 11437 3485 11471 3519
rect 11621 3485 11655 3519
rect 12449 3485 12483 3519
rect 12909 3485 12943 3519
rect 13006 3495 13040 3529
rect 13357 3463 13391 3497
rect 13553 3485 13587 3519
rect 13645 3485 13679 3519
rect 13829 3485 13863 3519
rect 14749 3485 14783 3519
rect 15577 3485 15611 3519
rect 15945 3485 15979 3519
rect 16313 3485 16347 3519
rect 16589 3485 16623 3519
rect 17601 3485 17635 3519
rect 18337 3485 18371 3519
rect 18521 3485 18555 3519
rect 19257 3485 19291 3519
rect 22477 3485 22511 3519
rect 22569 3485 22603 3519
rect 22845 3485 22879 3519
rect 23121 3485 23155 3519
rect 23305 3485 23339 3519
rect 23397 3485 23431 3519
rect 24041 3485 24075 3519
rect 25513 3485 25547 3519
rect 26709 3485 26743 3519
rect 36093 3485 36127 3519
rect 9413 3417 9447 3451
rect 10149 3417 10183 3451
rect 11161 3417 11195 3451
rect 12633 3417 12667 3451
rect 12817 3417 12851 3451
rect 14289 3417 14323 3451
rect 14473 3417 14507 3451
rect 27261 3417 27295 3451
rect 11069 3349 11103 3383
rect 16037 3349 16071 3383
rect 18245 3349 18279 3383
rect 19441 3349 19475 3383
rect 22937 3349 22971 3383
rect 26893 3349 26927 3383
rect 8217 3145 8251 3179
rect 12725 3145 12759 3179
rect 15669 3145 15703 3179
rect 16865 3145 16899 3179
rect 19165 3145 19199 3179
rect 21465 3145 21499 3179
rect 30297 3145 30331 3179
rect 36553 3145 36587 3179
rect 8769 3077 8803 3111
rect 9229 3077 9263 3111
rect 11161 3077 11195 3111
rect 14841 3077 14875 3111
rect 15025 3077 15059 3111
rect 23029 3077 23063 3111
rect 26525 3077 26559 3111
rect 36093 3077 36127 3111
rect 8033 3009 8067 3043
rect 8953 3009 8987 3043
rect 10793 3009 10827 3043
rect 10977 3009 11011 3043
rect 12725 3009 12759 3043
rect 12909 3009 12943 3043
rect 15577 3009 15611 3043
rect 15761 3009 15795 3043
rect 17049 3009 17083 3043
rect 17233 3009 17267 3043
rect 17325 3009 17359 3043
rect 18705 3009 18739 3043
rect 19717 3009 19751 3043
rect 22201 3007 22235 3041
rect 22753 3009 22787 3043
rect 22845 3009 22879 3043
rect 23397 3009 23431 3043
rect 24501 3009 24535 3043
rect 28549 3009 28583 3043
rect 8309 2941 8343 2975
rect 15209 2941 15243 2975
rect 17141 2941 17175 2975
rect 19993 2941 20027 2975
rect 22661 2941 22695 2975
rect 23489 2941 23523 2975
rect 24777 2941 24811 2975
rect 28825 2941 28859 2975
rect 8493 2873 8527 2907
rect 18981 2873 19015 2907
rect 23029 2873 23063 2907
rect 23765 2873 23799 2907
rect 36461 2873 36495 2907
rect 10701 2805 10735 2839
rect 22293 2805 22327 2839
rect 1593 2601 1627 2635
rect 8677 2601 8711 2635
rect 17693 2601 17727 2635
rect 26065 2601 26099 2635
rect 43269 2601 43303 2635
rect 25973 2533 26007 2567
rect 26157 2533 26191 2567
rect 19809 2465 19843 2499
rect 20453 2465 20487 2499
rect 1409 2397 1443 2431
rect 8493 2397 8527 2431
rect 17509 2397 17543 2431
rect 25605 2397 25639 2431
rect 26341 2397 26375 2431
rect 43453 2397 43487 2431
<< metal1 >>
rect 1104 45722 44620 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 44620 45722
rect 1104 45648 44620 45670
rect 14826 45500 14832 45552
rect 14884 45500 14890 45552
rect 32214 45500 32220 45552
rect 32272 45500 32278 45552
rect 1394 45432 1400 45484
rect 1452 45432 1458 45484
rect 6454 45432 6460 45484
rect 6512 45472 6518 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 6512 45444 6561 45472
rect 6512 45432 6518 45444
rect 6549 45441 6561 45444
rect 6595 45441 6607 45475
rect 14844 45472 14872 45500
rect 14921 45475 14979 45481
rect 14921 45472 14933 45475
rect 14844 45444 14933 45472
rect 6549 45435 6607 45441
rect 14921 45441 14933 45444
rect 14967 45441 14979 45475
rect 14921 45435 14979 45441
rect 23934 45432 23940 45484
rect 23992 45432 23998 45484
rect 32232 45472 32260 45500
rect 32493 45475 32551 45481
rect 32493 45472 32505 45475
rect 32232 45444 32505 45472
rect 32493 45441 32505 45444
rect 32539 45441 32551 45475
rect 32493 45435 32551 45441
rect 41230 45432 41236 45484
rect 41288 45472 41294 45484
rect 41509 45475 41567 45481
rect 41509 45472 41521 45475
rect 41288 45444 41521 45472
rect 41288 45432 41294 45444
rect 41509 45441 41521 45444
rect 41555 45441 41567 45475
rect 41509 45435 41567 45441
rect 1581 45271 1639 45277
rect 1581 45237 1593 45271
rect 1627 45268 1639 45271
rect 5902 45268 5908 45280
rect 1627 45240 5908 45268
rect 1627 45237 1639 45240
rect 1581 45231 1639 45237
rect 5902 45228 5908 45240
rect 5960 45228 5966 45280
rect 6733 45271 6791 45277
rect 6733 45237 6745 45271
rect 6779 45268 6791 45271
rect 7282 45268 7288 45280
rect 6779 45240 7288 45268
rect 6779 45237 6791 45240
rect 6733 45231 6791 45237
rect 7282 45228 7288 45240
rect 7340 45228 7346 45280
rect 15102 45228 15108 45280
rect 15160 45228 15166 45280
rect 24121 45271 24179 45277
rect 24121 45237 24133 45271
rect 24167 45268 24179 45271
rect 24302 45268 24308 45280
rect 24167 45240 24308 45268
rect 24167 45237 24179 45240
rect 24121 45231 24179 45237
rect 24302 45228 24308 45240
rect 24360 45228 24366 45280
rect 32306 45228 32312 45280
rect 32364 45228 32370 45280
rect 41322 45228 41328 45280
rect 41380 45228 41386 45280
rect 1104 45178 44620 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 44620 45178
rect 1104 45104 44620 45126
rect 15102 45024 15108 45076
rect 15160 45064 15166 45076
rect 15160 45036 18736 45064
rect 15160 45024 15166 45036
rect 5902 44956 5908 45008
rect 5960 44956 5966 45008
rect 16114 44996 16120 45008
rect 11900 44968 16120 44996
rect 5629 44931 5687 44937
rect 5629 44897 5641 44931
rect 5675 44928 5687 44931
rect 6638 44928 6644 44940
rect 5675 44900 6644 44928
rect 5675 44897 5687 44900
rect 5629 44891 5687 44897
rect 6638 44888 6644 44900
rect 6696 44928 6702 44940
rect 11900 44928 11928 44968
rect 16114 44956 16120 44968
rect 16172 44956 16178 45008
rect 18708 45005 18736 45036
rect 32306 45024 32312 45076
rect 32364 45024 32370 45076
rect 41322 45024 41328 45076
rect 41380 45024 41386 45076
rect 18693 44999 18751 45005
rect 18693 44965 18705 44999
rect 18739 44965 18751 44999
rect 18693 44959 18751 44965
rect 31941 44999 31999 45005
rect 31941 44965 31953 44999
rect 31987 44996 31999 44999
rect 32324 44996 32352 45024
rect 31987 44968 32352 44996
rect 36817 44999 36875 45005
rect 31987 44965 31999 44968
rect 31941 44959 31999 44965
rect 36817 44965 36829 44999
rect 36863 44996 36875 44999
rect 41340 44996 41368 45024
rect 36863 44968 41368 44996
rect 36863 44965 36875 44968
rect 36817 44959 36875 44965
rect 6696 44900 11928 44928
rect 11977 44931 12035 44937
rect 6696 44888 6702 44900
rect 11977 44897 11989 44931
rect 12023 44928 12035 44931
rect 16393 44931 16451 44937
rect 16393 44928 16405 44931
rect 12023 44900 12434 44928
rect 12023 44897 12035 44900
rect 11977 44891 12035 44897
rect 12406 44872 12434 44900
rect 16040 44900 16405 44928
rect 16040 44872 16068 44900
rect 16393 44897 16405 44900
rect 16439 44897 16451 44931
rect 16393 44891 16451 44897
rect 16482 44888 16488 44940
rect 16540 44928 16546 44940
rect 18417 44931 18475 44937
rect 18417 44928 18429 44931
rect 16540 44900 18429 44928
rect 16540 44888 16546 44900
rect 18417 44897 18429 44900
rect 18463 44897 18475 44931
rect 18417 44891 18475 44897
rect 18877 44931 18935 44937
rect 18877 44897 18889 44931
rect 18923 44928 18935 44931
rect 18923 44900 19564 44928
rect 18923 44897 18935 44900
rect 18877 44891 18935 44897
rect 9858 44820 9864 44872
rect 9916 44860 9922 44872
rect 10229 44863 10287 44869
rect 10229 44860 10241 44863
rect 9916 44832 10241 44860
rect 9916 44820 9922 44832
rect 10229 44829 10241 44832
rect 10275 44829 10287 44863
rect 12406 44832 12440 44872
rect 10229 44823 10287 44829
rect 12434 44820 12440 44832
rect 12492 44860 12498 44872
rect 12621 44863 12679 44869
rect 12621 44860 12633 44863
rect 12492 44832 12633 44860
rect 12492 44820 12498 44832
rect 12621 44829 12633 44832
rect 12667 44829 12679 44863
rect 12621 44823 12679 44829
rect 13633 44863 13691 44869
rect 13633 44829 13645 44863
rect 13679 44860 13691 44863
rect 14090 44860 14096 44872
rect 13679 44832 14096 44860
rect 13679 44829 13691 44832
rect 13633 44823 13691 44829
rect 14090 44820 14096 44832
rect 14148 44820 14154 44872
rect 15838 44820 15844 44872
rect 15896 44820 15902 44872
rect 16022 44820 16028 44872
rect 16080 44820 16086 44872
rect 16114 44820 16120 44872
rect 16172 44820 16178 44872
rect 10502 44752 10508 44804
rect 10560 44752 10566 44804
rect 11790 44792 11796 44804
rect 11730 44764 11796 44792
rect 11790 44752 11796 44764
rect 11848 44792 11854 44804
rect 14461 44795 14519 44801
rect 14461 44792 14473 44795
rect 11848 44764 14473 44792
rect 11848 44752 11854 44764
rect 14461 44761 14473 44764
rect 14507 44792 14519 44795
rect 14507 44764 16160 44792
rect 14507 44761 14519 44764
rect 14461 44755 14519 44761
rect 6086 44684 6092 44736
rect 6144 44684 6150 44736
rect 12066 44684 12072 44736
rect 12124 44684 12130 44736
rect 13446 44684 13452 44736
rect 13504 44684 13510 44736
rect 14369 44727 14427 44733
rect 14369 44693 14381 44727
rect 14415 44724 14427 44727
rect 14642 44724 14648 44736
rect 14415 44696 14648 44724
rect 14415 44693 14427 44696
rect 14369 44687 14427 44693
rect 14642 44684 14648 44696
rect 14700 44684 14706 44736
rect 16022 44684 16028 44736
rect 16080 44684 16086 44736
rect 16132 44724 16160 44764
rect 16850 44752 16856 44804
rect 16908 44752 16914 44804
rect 18432 44792 18460 44891
rect 19536 44869 19564 44900
rect 19521 44863 19579 44869
rect 19521 44829 19533 44863
rect 19567 44829 19579 44863
rect 19521 44823 19579 44829
rect 31573 44795 31631 44801
rect 31573 44792 31585 44795
rect 17696 44764 18000 44792
rect 18432 44764 31585 44792
rect 17696 44724 17724 44764
rect 16132 44696 17724 44724
rect 17862 44684 17868 44736
rect 17920 44684 17926 44736
rect 17972 44724 18000 44764
rect 31573 44761 31585 44764
rect 31619 44792 31631 44795
rect 36449 44795 36507 44801
rect 36449 44792 36461 44795
rect 31619 44764 36461 44792
rect 31619 44761 31631 44764
rect 31573 44755 31631 44761
rect 36449 44761 36461 44764
rect 36495 44792 36507 44795
rect 36998 44792 37004 44804
rect 36495 44764 37004 44792
rect 36495 44761 36507 44764
rect 36449 44755 36507 44761
rect 36998 44752 37004 44764
rect 37056 44752 37062 44804
rect 19150 44724 19156 44736
rect 17972 44696 19156 44724
rect 19150 44684 19156 44696
rect 19208 44684 19214 44736
rect 19705 44727 19763 44733
rect 19705 44693 19717 44727
rect 19751 44724 19763 44727
rect 19978 44724 19984 44736
rect 19751 44696 19984 44724
rect 19751 44693 19763 44696
rect 19705 44687 19763 44693
rect 19978 44684 19984 44696
rect 20036 44684 20042 44736
rect 32030 44684 32036 44736
rect 32088 44684 32094 44736
rect 36906 44684 36912 44736
rect 36964 44684 36970 44736
rect 1104 44634 44620 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 44620 44634
rect 1104 44560 44620 44582
rect 6086 44480 6092 44532
rect 6144 44480 6150 44532
rect 10502 44480 10508 44532
rect 10560 44520 10566 44532
rect 10781 44523 10839 44529
rect 10781 44520 10793 44523
rect 10560 44492 10793 44520
rect 10560 44480 10566 44492
rect 10781 44489 10793 44492
rect 10827 44489 10839 44523
rect 10781 44483 10839 44489
rect 11885 44523 11943 44529
rect 11885 44489 11897 44523
rect 11931 44520 11943 44523
rect 12066 44520 12072 44532
rect 11931 44492 12072 44520
rect 11931 44489 11943 44492
rect 11885 44483 11943 44489
rect 12066 44480 12072 44492
rect 12124 44480 12130 44532
rect 13446 44520 13452 44532
rect 13372 44492 13452 44520
rect 6104 44384 6132 44480
rect 13372 44461 13400 44492
rect 13446 44480 13452 44492
rect 13504 44480 13510 44532
rect 15838 44480 15844 44532
rect 15896 44520 15902 44532
rect 16669 44523 16727 44529
rect 16669 44520 16681 44523
rect 15896 44492 16681 44520
rect 15896 44480 15902 44492
rect 16669 44489 16681 44492
rect 16715 44489 16727 44523
rect 16669 44483 16727 44489
rect 19978 44480 19984 44532
rect 20036 44520 20042 44532
rect 20036 44492 20208 44520
rect 20036 44480 20042 44492
rect 8573 44455 8631 44461
rect 8573 44452 8585 44455
rect 7300 44424 8585 44452
rect 7300 44396 7328 44424
rect 8573 44421 8585 44424
rect 8619 44452 8631 44455
rect 13357 44455 13415 44461
rect 8619 44424 11928 44452
rect 8619 44421 8631 44424
rect 8573 44415 8631 44421
rect 6365 44387 6423 44393
rect 6365 44384 6377 44387
rect 6104 44356 6377 44384
rect 6365 44353 6377 44356
rect 6411 44353 6423 44387
rect 6365 44347 6423 44353
rect 7282 44344 7288 44396
rect 7340 44344 7346 44396
rect 8297 44387 8355 44393
rect 8297 44353 8309 44387
rect 8343 44353 8355 44387
rect 8297 44347 8355 44353
rect 10965 44387 11023 44393
rect 10965 44353 10977 44387
rect 11011 44384 11023 44387
rect 11011 44356 11560 44384
rect 11011 44353 11023 44356
rect 10965 44347 11023 44353
rect 6549 44183 6607 44189
rect 6549 44149 6561 44183
rect 6595 44180 6607 44183
rect 6914 44180 6920 44192
rect 6595 44152 6920 44180
rect 6595 44149 6607 44152
rect 6549 44143 6607 44149
rect 6914 44140 6920 44152
rect 6972 44140 6978 44192
rect 8202 44140 8208 44192
rect 8260 44140 8266 44192
rect 8312 44180 8340 44347
rect 11532 44257 11560 44356
rect 11517 44251 11575 44257
rect 11517 44217 11529 44251
rect 11563 44217 11575 44251
rect 11517 44211 11575 44217
rect 8849 44183 8907 44189
rect 8849 44180 8861 44183
rect 8312 44152 8861 44180
rect 8849 44149 8861 44152
rect 8895 44180 8907 44183
rect 11790 44180 11796 44192
rect 8895 44152 11796 44180
rect 8895 44149 8907 44152
rect 8849 44143 8907 44149
rect 11790 44140 11796 44152
rect 11848 44140 11854 44192
rect 11900 44180 11928 44424
rect 13357 44421 13369 44455
rect 13403 44421 13415 44455
rect 13357 44415 13415 44421
rect 18969 44455 19027 44461
rect 18969 44421 18981 44455
rect 19015 44452 19027 44455
rect 20070 44452 20076 44464
rect 19015 44424 20076 44452
rect 19015 44421 19027 44424
rect 18969 44415 19027 44421
rect 20070 44412 20076 44424
rect 20128 44412 20134 44464
rect 20180 44461 20208 44492
rect 32030 44480 32036 44532
rect 32088 44480 32094 44532
rect 36906 44480 36912 44532
rect 36964 44480 36970 44532
rect 20165 44455 20223 44461
rect 20165 44421 20177 44455
rect 20211 44421 20223 44455
rect 20165 44415 20223 44421
rect 20622 44412 20628 44464
rect 20680 44412 20686 44464
rect 14642 44384 14648 44396
rect 14490 44356 14648 44384
rect 14642 44344 14648 44356
rect 14700 44344 14706 44396
rect 17037 44387 17095 44393
rect 17037 44353 17049 44387
rect 17083 44384 17095 44387
rect 17862 44384 17868 44396
rect 17083 44356 17868 44384
rect 17083 44353 17095 44356
rect 17037 44347 17095 44353
rect 17862 44344 17868 44356
rect 17920 44344 17926 44396
rect 18506 44344 18512 44396
rect 18564 44384 18570 44396
rect 18785 44387 18843 44393
rect 18785 44384 18797 44387
rect 18564 44356 18797 44384
rect 18564 44344 18570 44356
rect 18785 44353 18797 44356
rect 18831 44353 18843 44387
rect 18785 44347 18843 44353
rect 19061 44387 19119 44393
rect 19061 44353 19073 44387
rect 19107 44353 19119 44387
rect 19061 44347 19119 44353
rect 11974 44276 11980 44328
rect 12032 44276 12038 44328
rect 12066 44276 12072 44328
rect 12124 44276 12130 44328
rect 12894 44276 12900 44328
rect 12952 44276 12958 44328
rect 13078 44276 13084 44328
rect 13136 44276 13142 44328
rect 14829 44319 14887 44325
rect 14829 44285 14841 44319
rect 14875 44316 14887 44319
rect 14918 44316 14924 44328
rect 14875 44288 14924 44316
rect 14875 44285 14887 44288
rect 14829 44279 14887 44285
rect 14918 44276 14924 44288
rect 14976 44316 14982 44328
rect 15473 44319 15531 44325
rect 15473 44316 15485 44319
rect 14976 44288 15485 44316
rect 14976 44276 14982 44288
rect 15473 44285 15485 44288
rect 15519 44285 15531 44319
rect 15473 44279 15531 44285
rect 17126 44276 17132 44328
rect 17184 44276 17190 44328
rect 17310 44276 17316 44328
rect 17368 44276 17374 44328
rect 17954 44276 17960 44328
rect 18012 44316 18018 44328
rect 19076 44316 19104 44347
rect 19150 44344 19156 44396
rect 19208 44384 19214 44396
rect 19337 44387 19395 44393
rect 19337 44384 19349 44387
rect 19208 44356 19349 44384
rect 19208 44344 19214 44356
rect 19337 44353 19349 44356
rect 19383 44353 19395 44387
rect 19337 44347 19395 44353
rect 31849 44387 31907 44393
rect 31849 44353 31861 44387
rect 31895 44384 31907 44387
rect 32048 44384 32076 44480
rect 31895 44356 32076 44384
rect 36449 44387 36507 44393
rect 31895 44353 31907 44356
rect 31849 44347 31907 44353
rect 36449 44353 36461 44387
rect 36495 44384 36507 44387
rect 36924 44384 36952 44480
rect 36495 44356 36952 44384
rect 36495 44353 36507 44356
rect 36449 44347 36507 44353
rect 18012 44288 19104 44316
rect 18012 44276 18018 44288
rect 19426 44276 19432 44328
rect 19484 44316 19490 44328
rect 19889 44319 19947 44325
rect 19889 44316 19901 44319
rect 19484 44288 19901 44316
rect 19484 44276 19490 44288
rect 19889 44285 19901 44288
rect 19935 44285 19947 44319
rect 27338 44316 27344 44328
rect 19889 44279 19947 44285
rect 19996 44288 27344 44316
rect 11992 44248 12020 44276
rect 12345 44251 12403 44257
rect 12345 44248 12357 44251
rect 11992 44220 12357 44248
rect 12345 44217 12357 44220
rect 12391 44217 12403 44251
rect 19996 44248 20024 44288
rect 27338 44276 27344 44288
rect 27396 44276 27402 44328
rect 12345 44211 12403 44217
rect 14384 44220 20024 44248
rect 14384 44180 14412 44220
rect 11900 44152 14412 44180
rect 14458 44140 14464 44192
rect 14516 44180 14522 44192
rect 14921 44183 14979 44189
rect 14921 44180 14933 44183
rect 14516 44152 14933 44180
rect 14516 44140 14522 44152
rect 14921 44149 14933 44152
rect 14967 44149 14979 44183
rect 14921 44143 14979 44149
rect 18598 44140 18604 44192
rect 18656 44140 18662 44192
rect 19521 44183 19579 44189
rect 19521 44149 19533 44183
rect 19567 44180 19579 44183
rect 20622 44180 20628 44192
rect 19567 44152 20628 44180
rect 19567 44149 19579 44152
rect 19521 44143 19579 44149
rect 20622 44140 20628 44152
rect 20680 44140 20686 44192
rect 21637 44183 21695 44189
rect 21637 44149 21649 44183
rect 21683 44180 21695 44183
rect 25406 44180 25412 44192
rect 21683 44152 25412 44180
rect 21683 44149 21695 44152
rect 21637 44143 21695 44149
rect 25406 44140 25412 44152
rect 25464 44140 25470 44192
rect 31662 44140 31668 44192
rect 31720 44140 31726 44192
rect 36265 44183 36323 44189
rect 36265 44149 36277 44183
rect 36311 44180 36323 44183
rect 36354 44180 36360 44192
rect 36311 44152 36360 44180
rect 36311 44149 36323 44152
rect 36265 44143 36323 44149
rect 36354 44140 36360 44152
rect 36412 44140 36418 44192
rect 1104 44090 44620 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 44620 44090
rect 1104 44016 44620 44038
rect 12345 43979 12403 43985
rect 12345 43945 12357 43979
rect 12391 43976 12403 43979
rect 12894 43976 12900 43988
rect 12391 43948 12900 43976
rect 12391 43945 12403 43948
rect 12345 43939 12403 43945
rect 12894 43936 12900 43948
rect 12952 43936 12958 43988
rect 14090 43936 14096 43988
rect 14148 43936 14154 43988
rect 15212 43948 16620 43976
rect 14182 43868 14188 43920
rect 14240 43908 14246 43920
rect 15013 43911 15071 43917
rect 15013 43908 15025 43911
rect 14240 43880 15025 43908
rect 14240 43868 14246 43880
rect 15013 43877 15025 43880
rect 15059 43877 15071 43911
rect 15013 43871 15071 43877
rect 6733 43843 6791 43849
rect 6733 43809 6745 43843
rect 6779 43840 6791 43843
rect 7006 43840 7012 43852
rect 6779 43812 7012 43840
rect 6779 43809 6791 43812
rect 6733 43803 6791 43809
rect 7006 43800 7012 43812
rect 7064 43800 7070 43852
rect 8202 43800 8208 43852
rect 8260 43840 8266 43852
rect 8260 43812 8340 43840
rect 8260 43800 8266 43812
rect 6914 43664 6920 43716
rect 6972 43704 6978 43716
rect 7009 43707 7067 43713
rect 7009 43704 7021 43707
rect 6972 43676 7021 43704
rect 6972 43664 6978 43676
rect 7009 43673 7021 43676
rect 7055 43673 7067 43707
rect 8312 43704 8340 43812
rect 12066 43800 12072 43852
rect 12124 43840 12130 43852
rect 14737 43843 14795 43849
rect 14737 43840 14749 43843
rect 12124 43812 14749 43840
rect 12124 43800 12130 43812
rect 14737 43809 14749 43812
rect 14783 43840 14795 43843
rect 15212 43840 15240 43948
rect 16592 43908 16620 43948
rect 17126 43936 17132 43988
rect 17184 43976 17190 43988
rect 17770 43976 17776 43988
rect 17184 43948 17776 43976
rect 17184 43936 17190 43948
rect 17770 43936 17776 43948
rect 17828 43936 17834 43988
rect 20530 43976 20536 43988
rect 17880 43948 20536 43976
rect 17310 43908 17316 43920
rect 16592 43880 17316 43908
rect 17310 43868 17316 43880
rect 17368 43908 17374 43920
rect 17880 43908 17908 43948
rect 20530 43936 20536 43948
rect 20588 43936 20594 43988
rect 17368 43880 17908 43908
rect 17368 43868 17374 43880
rect 14783 43812 15240 43840
rect 15289 43843 15347 43849
rect 14783 43809 14795 43812
rect 14737 43803 14795 43809
rect 15289 43809 15301 43843
rect 15335 43840 15347 43843
rect 16114 43840 16120 43852
rect 15335 43812 16120 43840
rect 15335 43809 15347 43812
rect 15289 43803 15347 43809
rect 16114 43800 16120 43812
rect 16172 43800 16178 43852
rect 17037 43843 17095 43849
rect 17037 43809 17049 43843
rect 17083 43840 17095 43843
rect 17129 43843 17187 43849
rect 17129 43840 17141 43843
rect 17083 43812 17141 43840
rect 17083 43809 17095 43812
rect 17037 43803 17095 43809
rect 17129 43809 17141 43812
rect 17175 43809 17187 43843
rect 17129 43803 17187 43809
rect 18598 43800 18604 43852
rect 18656 43840 18662 43852
rect 18969 43843 19027 43849
rect 18969 43840 18981 43843
rect 18656 43812 18981 43840
rect 18656 43800 18662 43812
rect 18969 43809 18981 43812
rect 19015 43809 19027 43843
rect 18969 43803 19027 43809
rect 20070 43800 20076 43852
rect 20128 43840 20134 43852
rect 21085 43843 21143 43849
rect 21085 43840 21097 43843
rect 20128 43812 21097 43840
rect 20128 43800 20134 43812
rect 21085 43809 21097 43812
rect 21131 43809 21143 43843
rect 21085 43803 21143 43809
rect 25406 43800 25412 43852
rect 25464 43800 25470 43852
rect 31573 43843 31631 43849
rect 31573 43809 31585 43843
rect 31619 43840 31631 43843
rect 31662 43840 31668 43852
rect 31619 43812 31668 43840
rect 31619 43809 31631 43812
rect 31573 43803 31631 43809
rect 31662 43800 31668 43812
rect 31720 43800 31726 43852
rect 36354 43800 36360 43852
rect 36412 43800 36418 43852
rect 9858 43732 9864 43784
rect 9916 43772 9922 43784
rect 10597 43775 10655 43781
rect 10597 43772 10609 43775
rect 9916 43744 10609 43772
rect 9916 43732 9922 43744
rect 10597 43741 10609 43744
rect 10643 43741 10655 43775
rect 10597 43735 10655 43741
rect 13170 43732 13176 43784
rect 13228 43732 13234 43784
rect 13906 43732 13912 43784
rect 13964 43732 13970 43784
rect 14458 43732 14464 43784
rect 14516 43732 14522 43784
rect 14918 43732 14924 43784
rect 14976 43732 14982 43784
rect 16850 43772 16856 43784
rect 16698 43744 16856 43772
rect 16850 43732 16856 43744
rect 16908 43732 16914 43784
rect 18141 43775 18199 43781
rect 18141 43741 18153 43775
rect 18187 43772 18199 43775
rect 19058 43772 19064 43784
rect 18187 43744 19064 43772
rect 18187 43741 18199 43744
rect 18141 43735 18199 43741
rect 19058 43732 19064 43744
rect 19116 43732 19122 43784
rect 19242 43732 19248 43784
rect 19300 43732 19306 43784
rect 20622 43732 20628 43784
rect 20680 43732 20686 43784
rect 20806 43732 20812 43784
rect 20864 43772 20870 43784
rect 21637 43775 21695 43781
rect 21637 43772 21649 43775
rect 20864 43744 21649 43772
rect 20864 43732 20870 43744
rect 21637 43741 21649 43744
rect 21683 43741 21695 43775
rect 21637 43735 21695 43741
rect 31202 43732 31208 43784
rect 31260 43772 31266 43784
rect 31297 43775 31355 43781
rect 31297 43772 31309 43775
rect 31260 43744 31309 43772
rect 31260 43732 31266 43744
rect 31297 43741 31309 43744
rect 31343 43741 31355 43775
rect 31297 43735 31355 43741
rect 36078 43732 36084 43784
rect 36136 43732 36142 43784
rect 8234 43676 9444 43704
rect 7009 43667 7067 43673
rect 8478 43596 8484 43648
rect 8536 43596 8542 43648
rect 9416 43636 9444 43676
rect 10870 43664 10876 43716
rect 10928 43664 10934 43716
rect 10980 43676 11362 43704
rect 10980 43648 11008 43676
rect 15562 43664 15568 43716
rect 15620 43664 15626 43716
rect 19521 43707 19579 43713
rect 19521 43704 19533 43707
rect 18340 43676 19533 43704
rect 10962 43636 10968 43648
rect 9416 43608 10968 43636
rect 10962 43596 10968 43608
rect 11020 43596 11026 43648
rect 12526 43596 12532 43648
rect 12584 43596 12590 43648
rect 13265 43639 13323 43645
rect 13265 43605 13277 43639
rect 13311 43636 13323 43639
rect 13814 43636 13820 43648
rect 13311 43608 13820 43636
rect 13311 43605 13323 43608
rect 13265 43599 13323 43605
rect 13814 43596 13820 43608
rect 13872 43636 13878 43648
rect 18340 43645 18368 43676
rect 19521 43673 19533 43676
rect 19567 43673 19579 43707
rect 19521 43667 19579 43673
rect 32582 43664 32588 43716
rect 32640 43664 32646 43716
rect 36814 43664 36820 43716
rect 36872 43664 36878 43716
rect 43438 43664 43444 43716
rect 43496 43664 43502 43716
rect 44269 43707 44327 43713
rect 44269 43673 44281 43707
rect 44315 43704 44327 43707
rect 44634 43704 44640 43716
rect 44315 43676 44640 43704
rect 44315 43673 44327 43676
rect 44269 43667 44327 43673
rect 44634 43664 44640 43676
rect 44692 43664 44698 43716
rect 14553 43639 14611 43645
rect 14553 43636 14565 43639
rect 13872 43608 14565 43636
rect 13872 43596 13878 43608
rect 14553 43605 14565 43608
rect 14599 43605 14611 43639
rect 14553 43599 14611 43605
rect 18325 43639 18383 43645
rect 18325 43605 18337 43639
rect 18371 43605 18383 43639
rect 18325 43599 18383 43605
rect 18414 43596 18420 43648
rect 18472 43596 18478 43648
rect 20990 43596 20996 43648
rect 21048 43596 21054 43648
rect 26053 43639 26111 43645
rect 26053 43605 26065 43639
rect 26099 43636 26111 43639
rect 29178 43636 29184 43648
rect 26099 43608 29184 43636
rect 26099 43605 26111 43608
rect 26053 43599 26111 43605
rect 29178 43596 29184 43608
rect 29236 43596 29242 43648
rect 33042 43596 33048 43648
rect 33100 43596 33106 43648
rect 37826 43596 37832 43648
rect 37884 43596 37890 43648
rect 1104 43546 44620 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 44620 43546
rect 1104 43472 44620 43494
rect 10870 43392 10876 43444
rect 10928 43432 10934 43444
rect 11517 43435 11575 43441
rect 11517 43432 11529 43435
rect 10928 43404 11529 43432
rect 10928 43392 10934 43404
rect 11517 43401 11529 43404
rect 11563 43401 11575 43435
rect 11517 43395 11575 43401
rect 12526 43392 12532 43444
rect 12584 43392 12590 43444
rect 13906 43392 13912 43444
rect 13964 43432 13970 43444
rect 14461 43435 14519 43441
rect 14461 43432 14473 43435
rect 13964 43404 14473 43432
rect 13964 43392 13970 43404
rect 14461 43401 14473 43404
rect 14507 43401 14519 43435
rect 14461 43395 14519 43401
rect 15562 43392 15568 43444
rect 15620 43432 15626 43444
rect 15749 43435 15807 43441
rect 15749 43432 15761 43435
rect 15620 43404 15761 43432
rect 15620 43392 15626 43404
rect 15749 43401 15761 43404
rect 15795 43401 15807 43435
rect 15749 43395 15807 43401
rect 17770 43392 17776 43444
rect 17828 43432 17834 43444
rect 17865 43435 17923 43441
rect 17865 43432 17877 43435
rect 17828 43404 17877 43432
rect 17828 43392 17834 43404
rect 17865 43401 17877 43404
rect 17911 43401 17923 43435
rect 17865 43395 17923 43401
rect 19889 43435 19947 43441
rect 19889 43401 19901 43435
rect 19935 43401 19947 43435
rect 19889 43395 19947 43401
rect 20349 43435 20407 43441
rect 20349 43401 20361 43435
rect 20395 43432 20407 43435
rect 20990 43432 20996 43444
rect 20395 43404 20996 43432
rect 20395 43401 20407 43404
rect 20349 43395 20407 43401
rect 10965 43367 11023 43373
rect 10965 43333 10977 43367
rect 11011 43364 11023 43367
rect 11974 43364 11980 43376
rect 11011 43336 11980 43364
rect 11011 43333 11023 43336
rect 10965 43327 11023 43333
rect 11974 43324 11980 43336
rect 12032 43324 12038 43376
rect 12544 43364 12572 43392
rect 12989 43367 13047 43373
rect 12989 43364 13001 43367
rect 12544 43336 13001 43364
rect 12989 43333 13001 43336
rect 13035 43333 13047 43367
rect 19904 43364 19932 43395
rect 20990 43392 20996 43404
rect 21048 43392 21054 43444
rect 31202 43432 31208 43444
rect 28920 43404 31208 43432
rect 20806 43364 20812 43376
rect 19904 43336 20812 43364
rect 12989 43327 13047 43333
rect 20806 43324 20812 43336
rect 20864 43324 20870 43376
rect 10870 43256 10876 43308
rect 10928 43256 10934 43308
rect 11149 43299 11207 43305
rect 11149 43265 11161 43299
rect 11195 43296 11207 43299
rect 11195 43268 12204 43296
rect 11195 43265 11207 43268
rect 11149 43259 11207 43265
rect 11333 43231 11391 43237
rect 11333 43197 11345 43231
rect 11379 43228 11391 43231
rect 12069 43231 12127 43237
rect 12069 43228 12081 43231
rect 11379 43200 12081 43228
rect 11379 43197 11391 43200
rect 11333 43191 11391 43197
rect 12069 43197 12081 43200
rect 12115 43197 12127 43231
rect 12176 43228 12204 43268
rect 12434 43256 12440 43308
rect 12492 43256 12498 43308
rect 14642 43296 14648 43308
rect 14122 43268 14648 43296
rect 14642 43256 14648 43268
rect 14700 43256 14706 43308
rect 16114 43256 16120 43308
rect 16172 43296 16178 43308
rect 16172 43268 17632 43296
rect 16172 43256 16178 43268
rect 12618 43228 12624 43240
rect 12176 43200 12624 43228
rect 12069 43191 12127 43197
rect 12618 43188 12624 43200
rect 12676 43188 12682 43240
rect 12713 43231 12771 43237
rect 12713 43197 12725 43231
rect 12759 43197 12771 43231
rect 12713 43191 12771 43197
rect 12526 43052 12532 43104
rect 12584 43052 12590 43104
rect 12728 43092 12756 43191
rect 14826 43188 14832 43240
rect 14884 43228 14890 43240
rect 15565 43231 15623 43237
rect 15565 43228 15577 43231
rect 14884 43200 15577 43228
rect 14884 43188 14890 43200
rect 15565 43197 15577 43200
rect 15611 43197 15623 43231
rect 15565 43191 15623 43197
rect 16393 43231 16451 43237
rect 16393 43197 16405 43231
rect 16439 43197 16451 43231
rect 16393 43191 16451 43197
rect 16408 43160 16436 43191
rect 17310 43188 17316 43240
rect 17368 43188 17374 43240
rect 17604 43228 17632 43268
rect 17678 43256 17684 43308
rect 17736 43256 17742 43308
rect 17954 43256 17960 43308
rect 18012 43256 18018 43308
rect 20622 43296 20628 43308
rect 19550 43268 20628 43296
rect 20622 43256 20628 43268
rect 20680 43256 20686 43308
rect 21008 43305 21036 43392
rect 28920 43305 28948 43404
rect 31202 43392 31208 43404
rect 31260 43392 31266 43444
rect 33042 43392 33048 43444
rect 33100 43432 33106 43444
rect 33100 43404 33456 43432
rect 33100 43392 33106 43404
rect 29178 43324 29184 43376
rect 29236 43324 29242 43376
rect 20993 43299 21051 43305
rect 20993 43265 21005 43299
rect 21039 43265 21051 43299
rect 20993 43259 21051 43265
rect 28905 43299 28963 43305
rect 28905 43265 28917 43299
rect 28951 43265 28963 43299
rect 32582 43296 32588 43308
rect 30314 43282 32588 43296
rect 28905 43259 28963 43265
rect 30300 43268 32588 43282
rect 18138 43228 18144 43240
rect 17604 43200 18144 43228
rect 18138 43188 18144 43200
rect 18196 43188 18202 43240
rect 18414 43188 18420 43240
rect 18472 43188 18478 43240
rect 19058 43188 19064 43240
rect 19116 43228 19122 43240
rect 19116 43200 19472 43228
rect 19116 43188 19122 43200
rect 17497 43163 17555 43169
rect 17497 43160 17509 43163
rect 16408 43132 17509 43160
rect 17497 43129 17509 43132
rect 17543 43129 17555 43163
rect 19444 43160 19472 43200
rect 20070 43188 20076 43240
rect 20128 43228 20134 43240
rect 20441 43231 20499 43237
rect 20441 43228 20453 43231
rect 20128 43200 20453 43228
rect 20128 43188 20134 43200
rect 20441 43197 20453 43200
rect 20487 43197 20499 43231
rect 20441 43191 20499 43197
rect 20530 43188 20536 43240
rect 20588 43188 20594 43240
rect 24026 43228 24032 43240
rect 22066 43200 24032 43228
rect 19981 43163 20039 43169
rect 19981 43160 19993 43163
rect 19444 43132 19993 43160
rect 17497 43123 17555 43129
rect 19981 43129 19993 43132
rect 20027 43129 20039 43163
rect 22066 43160 22094 43200
rect 24026 43188 24032 43200
rect 24084 43188 24090 43240
rect 27154 43188 27160 43240
rect 27212 43228 27218 43240
rect 30300 43228 30328 43268
rect 32582 43256 32588 43268
rect 32640 43256 32646 43308
rect 33428 43305 33456 43404
rect 40586 43364 40592 43376
rect 40434 43336 40592 43364
rect 40586 43324 40592 43336
rect 40644 43324 40650 43376
rect 33413 43299 33471 43305
rect 33413 43265 33425 43299
rect 33459 43265 33471 43299
rect 33413 43259 33471 43265
rect 27212 43200 30328 43228
rect 36173 43231 36231 43237
rect 27212 43188 27218 43200
rect 36173 43197 36185 43231
rect 36219 43228 36231 43231
rect 36446 43228 36452 43240
rect 36219 43200 36452 43228
rect 36219 43197 36231 43200
rect 36173 43191 36231 43197
rect 36446 43188 36452 43200
rect 36504 43188 36510 43240
rect 38654 43188 38660 43240
rect 38712 43228 38718 43240
rect 38933 43231 38991 43237
rect 38933 43228 38945 43231
rect 38712 43200 38945 43228
rect 38712 43188 38718 43200
rect 38933 43197 38945 43200
rect 38979 43197 38991 43231
rect 38933 43191 38991 43197
rect 39206 43188 39212 43240
rect 39264 43188 39270 43240
rect 19981 43123 20039 43129
rect 20088 43132 22094 43160
rect 13078 43092 13084 43104
rect 12728 43064 13084 43092
rect 13078 43052 13084 43064
rect 13136 43052 13142 43104
rect 15010 43052 15016 43104
rect 15068 43052 15074 43104
rect 16758 43052 16764 43104
rect 16816 43052 16822 43104
rect 17218 43052 17224 43104
rect 17276 43092 17282 43104
rect 20088 43092 20116 43132
rect 24302 43120 24308 43172
rect 24360 43120 24366 43172
rect 17276 43064 20116 43092
rect 20901 43095 20959 43101
rect 17276 43052 17282 43064
rect 20901 43061 20913 43095
rect 20947 43092 20959 43095
rect 21450 43092 21456 43104
rect 20947 43064 21456 43092
rect 20947 43061 20959 43064
rect 20901 43055 20959 43061
rect 21450 43052 21456 43064
rect 21508 43052 21514 43104
rect 24489 43095 24547 43101
rect 24489 43061 24501 43095
rect 24535 43092 24547 43095
rect 24854 43092 24860 43104
rect 24535 43064 24860 43092
rect 24535 43061 24547 43064
rect 24489 43055 24547 43061
rect 24854 43052 24860 43064
rect 24912 43052 24918 43104
rect 30653 43095 30711 43101
rect 30653 43061 30665 43095
rect 30699 43092 30711 43095
rect 31294 43092 31300 43104
rect 30699 43064 31300 43092
rect 30699 43061 30711 43064
rect 30653 43055 30711 43061
rect 31294 43052 31300 43064
rect 31352 43052 31358 43104
rect 34054 43052 34060 43104
rect 34112 43052 34118 43104
rect 35526 43052 35532 43104
rect 35584 43052 35590 43104
rect 40678 43052 40684 43104
rect 40736 43052 40742 43104
rect 1104 43002 44620 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 44620 43002
rect 1104 42928 44620 42950
rect 12618 42848 12624 42900
rect 12676 42888 12682 42900
rect 12805 42891 12863 42897
rect 12805 42888 12817 42891
rect 12676 42860 12817 42888
rect 12676 42848 12682 42860
rect 12805 42857 12817 42860
rect 12851 42857 12863 42891
rect 12805 42851 12863 42857
rect 13170 42848 13176 42900
rect 13228 42888 13234 42900
rect 13449 42891 13507 42897
rect 13449 42888 13461 42891
rect 13228 42860 13461 42888
rect 13228 42848 13234 42860
rect 13449 42857 13461 42860
rect 13495 42857 13507 42891
rect 16669 42891 16727 42897
rect 13449 42851 13507 42857
rect 13556 42860 16620 42888
rect 13556 42820 13584 42860
rect 7944 42792 13584 42820
rect 16592 42820 16620 42860
rect 16669 42857 16681 42891
rect 16715 42888 16727 42891
rect 17310 42888 17316 42900
rect 16715 42860 17316 42888
rect 16715 42857 16727 42860
rect 16669 42851 16727 42857
rect 17310 42848 17316 42860
rect 17368 42848 17374 42900
rect 18138 42848 18144 42900
rect 18196 42888 18202 42900
rect 18196 42860 18644 42888
rect 18196 42848 18202 42860
rect 17218 42820 17224 42832
rect 16592 42792 17224 42820
rect 6638 42712 6644 42764
rect 6696 42712 6702 42764
rect 5534 42644 5540 42696
rect 5592 42684 5598 42696
rect 5813 42687 5871 42693
rect 5813 42684 5825 42687
rect 5592 42656 5825 42684
rect 5592 42644 5598 42656
rect 5813 42653 5825 42656
rect 5859 42684 5871 42687
rect 7944 42684 7972 42792
rect 17218 42780 17224 42792
rect 17276 42780 17282 42832
rect 18616 42764 18644 42860
rect 24026 42848 24032 42900
rect 24084 42888 24090 42900
rect 39025 42891 39083 42897
rect 24084 42860 36584 42888
rect 24084 42848 24090 42860
rect 36556 42820 36584 42860
rect 39025 42857 39037 42891
rect 39071 42888 39083 42891
rect 39206 42888 39212 42900
rect 39071 42860 39212 42888
rect 39071 42857 39083 42860
rect 39025 42851 39083 42857
rect 39206 42848 39212 42860
rect 39264 42848 39270 42900
rect 43438 42848 43444 42900
rect 43496 42848 43502 42900
rect 43456 42820 43484 42848
rect 36556 42792 43484 42820
rect 12345 42755 12403 42761
rect 12345 42721 12357 42755
rect 12391 42752 12403 42755
rect 12897 42755 12955 42761
rect 12897 42752 12909 42755
rect 12391 42724 12909 42752
rect 12391 42721 12403 42724
rect 12345 42715 12403 42721
rect 12897 42721 12909 42724
rect 12943 42721 12955 42755
rect 14550 42752 14556 42764
rect 12897 42715 12955 42721
rect 13096 42724 14556 42752
rect 5859 42656 7972 42684
rect 9585 42687 9643 42693
rect 5859 42653 5871 42656
rect 5813 42647 5871 42653
rect 9585 42653 9597 42687
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 9861 42687 9919 42693
rect 9861 42653 9873 42687
rect 9907 42684 9919 42687
rect 10134 42684 10140 42696
rect 9907 42656 10140 42684
rect 9907 42653 9919 42656
rect 9861 42647 9919 42653
rect 8846 42576 8852 42628
rect 8904 42616 8910 42628
rect 9600 42616 9628 42647
rect 10134 42644 10140 42656
rect 10192 42644 10198 42696
rect 10962 42644 10968 42696
rect 11020 42684 11026 42696
rect 11701 42687 11759 42693
rect 11701 42684 11713 42687
rect 11020 42656 11713 42684
rect 11020 42644 11026 42656
rect 11701 42653 11713 42656
rect 11747 42653 11759 42687
rect 11701 42647 11759 42653
rect 11974 42644 11980 42696
rect 12032 42684 12038 42696
rect 13096 42693 13124 42724
rect 14550 42712 14556 42724
rect 14608 42712 14614 42764
rect 14642 42712 14648 42764
rect 14700 42752 14706 42764
rect 14700 42724 16436 42752
rect 14700 42712 14706 42724
rect 12437 42687 12495 42693
rect 12437 42684 12449 42687
rect 12032 42656 12449 42684
rect 12032 42644 12038 42656
rect 12437 42653 12449 42656
rect 12483 42653 12495 42687
rect 12437 42647 12495 42653
rect 12621 42687 12679 42693
rect 12621 42653 12633 42687
rect 12667 42684 12679 42687
rect 13081 42687 13139 42693
rect 13081 42684 13093 42687
rect 12667 42656 13093 42684
rect 12667 42653 12679 42656
rect 12621 42647 12679 42653
rect 13081 42653 13093 42656
rect 13127 42653 13139 42687
rect 13081 42647 13139 42653
rect 13633 42687 13691 42693
rect 13633 42653 13645 42687
rect 13679 42653 13691 42687
rect 13633 42647 13691 42653
rect 13265 42619 13323 42625
rect 8904 42588 12940 42616
rect 8904 42576 8910 42588
rect 8938 42508 8944 42560
rect 8996 42508 9002 42560
rect 9490 42508 9496 42560
rect 9548 42548 9554 42560
rect 9677 42551 9735 42557
rect 9677 42548 9689 42551
rect 9548 42520 9689 42548
rect 9548 42508 9554 42520
rect 9677 42517 9689 42520
rect 9723 42517 9735 42551
rect 9677 42511 9735 42517
rect 10042 42508 10048 42560
rect 10100 42548 10106 42560
rect 10321 42551 10379 42557
rect 10321 42548 10333 42551
rect 10100 42520 10333 42548
rect 10100 42508 10106 42520
rect 10321 42517 10333 42520
rect 10367 42517 10379 42551
rect 12912 42548 12940 42588
rect 13265 42585 13277 42619
rect 13311 42616 13323 42619
rect 13648 42616 13676 42647
rect 13814 42644 13820 42696
rect 13872 42644 13878 42696
rect 13906 42644 13912 42696
rect 13964 42644 13970 42696
rect 13998 42644 14004 42696
rect 14056 42684 14062 42696
rect 14921 42687 14979 42693
rect 14921 42684 14933 42687
rect 14056 42656 14933 42684
rect 14056 42644 14062 42656
rect 14921 42653 14933 42656
rect 14967 42653 14979 42687
rect 14921 42647 14979 42653
rect 13311 42588 14964 42616
rect 13311 42585 13323 42588
rect 13265 42579 13323 42585
rect 14936 42560 14964 42588
rect 15194 42576 15200 42628
rect 15252 42576 15258 42628
rect 16408 42616 16436 42724
rect 18598 42712 18604 42764
rect 18656 42752 18662 42764
rect 19242 42752 19248 42764
rect 18656 42724 19248 42752
rect 18656 42712 18662 42724
rect 19242 42712 19248 42724
rect 19300 42712 19306 42764
rect 38838 42712 38844 42764
rect 38896 42712 38902 42764
rect 40497 42755 40555 42761
rect 40497 42721 40509 42755
rect 40543 42752 40555 42755
rect 40678 42752 40684 42764
rect 40543 42724 40684 42752
rect 40543 42721 40555 42724
rect 40497 42715 40555 42721
rect 40678 42712 40684 42724
rect 40736 42712 40742 42764
rect 16850 42644 16856 42696
rect 16908 42684 16914 42696
rect 21637 42687 21695 42693
rect 21637 42684 21649 42687
rect 16908 42656 17250 42684
rect 18616 42656 21649 42684
rect 16908 42644 16914 42656
rect 16868 42616 16896 42644
rect 16408 42602 16896 42616
rect 16422 42588 16896 42602
rect 18322 42576 18328 42628
rect 18380 42576 18386 42628
rect 14090 42548 14096 42560
rect 12912 42520 14096 42548
rect 10321 42511 10379 42517
rect 14090 42508 14096 42520
rect 14148 42508 14154 42560
rect 14918 42508 14924 42560
rect 14976 42508 14982 42560
rect 16853 42551 16911 42557
rect 16853 42517 16865 42551
rect 16899 42548 16911 42551
rect 17034 42548 17040 42560
rect 16899 42520 17040 42548
rect 16899 42517 16911 42520
rect 16853 42511 16911 42517
rect 17034 42508 17040 42520
rect 17092 42548 17098 42560
rect 18616 42548 18644 42656
rect 21637 42653 21649 42656
rect 21683 42653 21695 42687
rect 21637 42647 21695 42653
rect 24854 42644 24860 42696
rect 24912 42684 24918 42696
rect 24949 42687 25007 42693
rect 24949 42684 24961 42687
rect 24912 42656 24961 42684
rect 24912 42644 24918 42656
rect 24949 42653 24961 42656
rect 24995 42653 25007 42687
rect 24949 42647 25007 42653
rect 34701 42687 34759 42693
rect 34701 42653 34713 42687
rect 34747 42653 34759 42687
rect 36814 42684 36820 42696
rect 36110 42656 36820 42684
rect 34701 42647 34759 42653
rect 20990 42576 20996 42628
rect 21048 42576 21054 42628
rect 34716 42616 34744 42647
rect 36814 42644 36820 42656
rect 36872 42684 36878 42696
rect 37090 42684 37096 42696
rect 36872 42656 37096 42684
rect 36872 42644 36878 42656
rect 37090 42644 37096 42656
rect 37148 42644 37154 42696
rect 38749 42687 38807 42693
rect 38749 42653 38761 42687
rect 38795 42684 38807 42687
rect 39853 42687 39911 42693
rect 39853 42684 39865 42687
rect 38795 42656 39865 42684
rect 38795 42653 38807 42656
rect 38749 42647 38807 42653
rect 39853 42653 39865 42656
rect 39899 42653 39911 42687
rect 39853 42647 39911 42653
rect 40770 42644 40776 42696
rect 40828 42644 40834 42696
rect 34716 42588 34836 42616
rect 34808 42560 34836 42588
rect 34974 42576 34980 42628
rect 35032 42576 35038 42628
rect 17092 42520 18644 42548
rect 17092 42508 17098 42520
rect 19150 42508 19156 42560
rect 19208 42548 19214 42560
rect 21085 42551 21143 42557
rect 21085 42548 21097 42551
rect 19208 42520 21097 42548
rect 19208 42508 19214 42520
rect 21085 42517 21097 42520
rect 21131 42517 21143 42551
rect 21085 42511 21143 42517
rect 25130 42508 25136 42560
rect 25188 42508 25194 42560
rect 34790 42508 34796 42560
rect 34848 42508 34854 42560
rect 36446 42508 36452 42560
rect 36504 42548 36510 42560
rect 36906 42548 36912 42560
rect 36504 42520 36912 42548
rect 36504 42508 36510 42520
rect 36906 42508 36912 42520
rect 36964 42508 36970 42560
rect 40310 42508 40316 42560
rect 40368 42548 40374 42560
rect 40589 42551 40647 42557
rect 40589 42548 40601 42551
rect 40368 42520 40601 42548
rect 40368 42508 40374 42520
rect 40589 42517 40601 42520
rect 40635 42517 40647 42551
rect 40589 42511 40647 42517
rect 1104 42458 44620 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 44620 42458
rect 1104 42384 44620 42406
rect 9858 42344 9864 42356
rect 7116 42316 9864 42344
rect 7006 42168 7012 42220
rect 7064 42208 7070 42220
rect 7116 42217 7144 42316
rect 8846 42236 8852 42288
rect 8904 42236 8910 42288
rect 7101 42211 7159 42217
rect 7101 42208 7113 42211
rect 7064 42180 7113 42208
rect 7064 42168 7070 42180
rect 7101 42177 7113 42180
rect 7147 42177 7159 42211
rect 7101 42171 7159 42177
rect 7374 42100 7380 42152
rect 7432 42100 7438 42152
rect 8496 42072 8524 42194
rect 8864 42149 8892 42236
rect 8956 42217 8984 42316
rect 9858 42304 9864 42316
rect 9916 42304 9922 42356
rect 10689 42347 10747 42353
rect 10689 42313 10701 42347
rect 10735 42344 10747 42347
rect 10962 42344 10968 42356
rect 10735 42316 10968 42344
rect 10735 42313 10747 42316
rect 10689 42307 10747 42313
rect 10962 42304 10968 42316
rect 11020 42304 11026 42356
rect 13280 42316 14780 42344
rect 13280 42288 13308 42316
rect 9217 42279 9275 42285
rect 9217 42245 9229 42279
rect 9263 42276 9275 42279
rect 9490 42276 9496 42288
rect 9263 42248 9496 42276
rect 9263 42245 9275 42248
rect 9217 42239 9275 42245
rect 9490 42236 9496 42248
rect 9548 42236 9554 42288
rect 11790 42276 11796 42288
rect 10442 42262 11796 42276
rect 10428 42248 11796 42262
rect 8941 42211 8999 42217
rect 8941 42177 8953 42211
rect 8987 42177 8999 42211
rect 8941 42171 8999 42177
rect 8849 42143 8907 42149
rect 8849 42109 8861 42143
rect 8895 42109 8907 42143
rect 10428 42140 10456 42248
rect 11790 42236 11796 42248
rect 11848 42236 11854 42288
rect 13262 42236 13268 42288
rect 13320 42236 13326 42288
rect 14642 42276 14648 42288
rect 14582 42248 14648 42276
rect 14642 42236 14648 42248
rect 14700 42236 14706 42288
rect 14752 42276 14780 42316
rect 14826 42304 14832 42356
rect 14884 42304 14890 42356
rect 15194 42304 15200 42356
rect 15252 42344 15258 42356
rect 15565 42347 15623 42353
rect 15565 42344 15577 42347
rect 15252 42316 15577 42344
rect 15252 42304 15258 42316
rect 15565 42313 15577 42316
rect 15611 42313 15623 42347
rect 15565 42307 15623 42313
rect 16025 42347 16083 42353
rect 16025 42313 16037 42347
rect 16071 42344 16083 42347
rect 16666 42344 16672 42356
rect 16071 42316 16672 42344
rect 16071 42313 16083 42316
rect 16025 42307 16083 42313
rect 16666 42304 16672 42316
rect 16724 42344 16730 42356
rect 17678 42344 17684 42356
rect 16724 42316 17684 42344
rect 16724 42304 16730 42316
rect 17678 42304 17684 42316
rect 17736 42304 17742 42356
rect 17865 42347 17923 42353
rect 17865 42313 17877 42347
rect 17911 42344 17923 42347
rect 18322 42344 18328 42356
rect 17911 42316 18328 42344
rect 17911 42313 17923 42316
rect 17865 42307 17923 42313
rect 18322 42304 18328 42316
rect 18380 42304 18386 42356
rect 18414 42304 18420 42356
rect 18472 42304 18478 42356
rect 19150 42344 19156 42356
rect 18524 42316 19156 42344
rect 15289 42279 15347 42285
rect 14752 42248 15240 42276
rect 11885 42211 11943 42217
rect 11885 42177 11897 42211
rect 11931 42208 11943 42211
rect 12345 42211 12403 42217
rect 12345 42208 12357 42211
rect 11931 42180 12357 42208
rect 11931 42177 11943 42180
rect 11885 42171 11943 42177
rect 12345 42177 12357 42180
rect 12391 42177 12403 42211
rect 12345 42171 12403 42177
rect 14918 42168 14924 42220
rect 14976 42168 14982 42220
rect 15010 42168 15016 42220
rect 15068 42208 15074 42220
rect 15212 42217 15240 42248
rect 15289 42245 15301 42279
rect 15335 42276 15347 42279
rect 16758 42276 16764 42288
rect 15335 42248 16764 42276
rect 15335 42245 15347 42248
rect 15289 42239 15347 42245
rect 16758 42236 16764 42248
rect 16816 42236 16822 42288
rect 18432 42276 18460 42304
rect 18340 42248 18460 42276
rect 15197 42211 15255 42217
rect 15068 42180 15113 42208
rect 15068 42168 15074 42180
rect 15197 42177 15209 42211
rect 15243 42177 15255 42211
rect 15197 42171 15255 42177
rect 15427 42211 15485 42217
rect 15427 42177 15439 42211
rect 15473 42208 15485 42211
rect 15562 42208 15568 42220
rect 15473 42180 15568 42208
rect 15473 42177 15485 42180
rect 15427 42171 15485 42177
rect 15562 42168 15568 42180
rect 15620 42168 15626 42220
rect 15657 42211 15715 42217
rect 15657 42177 15669 42211
rect 15703 42177 15715 42211
rect 15657 42171 15715 42177
rect 15841 42211 15899 42217
rect 15841 42177 15853 42211
rect 15887 42177 15899 42211
rect 15841 42171 15899 42177
rect 8849 42103 8907 42109
rect 8956 42112 10456 42140
rect 8956 42072 8984 42112
rect 11238 42100 11244 42152
rect 11296 42140 11302 42152
rect 11977 42143 12035 42149
rect 11977 42140 11989 42143
rect 11296 42112 11989 42140
rect 11296 42100 11302 42112
rect 11977 42109 11989 42112
rect 12023 42109 12035 42143
rect 11977 42103 12035 42109
rect 12158 42100 12164 42152
rect 12216 42100 12222 42152
rect 12897 42143 12955 42149
rect 12897 42140 12909 42143
rect 12406 42112 12909 42140
rect 8496 42044 8984 42072
rect 11514 41964 11520 42016
rect 11572 41964 11578 42016
rect 11974 41964 11980 42016
rect 12032 42004 12038 42016
rect 12406 42004 12434 42112
rect 12897 42109 12909 42112
rect 12943 42109 12955 42143
rect 12897 42103 12955 42109
rect 13078 42100 13084 42152
rect 13136 42100 13142 42152
rect 13354 42100 13360 42152
rect 13412 42100 13418 42152
rect 14090 42100 14096 42152
rect 14148 42140 14154 42152
rect 15672 42140 15700 42171
rect 14148 42112 15700 42140
rect 14148 42100 14154 42112
rect 12032 41976 12434 42004
rect 13096 42004 13124 42100
rect 14458 42032 14464 42084
rect 14516 42032 14522 42084
rect 14550 42032 14556 42084
rect 14608 42072 14614 42084
rect 15856 42072 15884 42171
rect 17402 42168 17408 42220
rect 17460 42168 17466 42220
rect 18340 42217 18368 42248
rect 18524 42217 18552 42316
rect 19150 42304 19156 42316
rect 19208 42304 19214 42356
rect 19242 42304 19248 42356
rect 19300 42344 19306 42356
rect 20346 42344 20352 42356
rect 19300 42316 20352 42344
rect 19300 42304 19306 42316
rect 20346 42304 20352 42316
rect 20404 42344 20410 42356
rect 20404 42316 21864 42344
rect 20404 42304 20410 42316
rect 19260 42276 19288 42304
rect 19076 42248 19288 42276
rect 18325 42211 18383 42217
rect 18325 42177 18337 42211
rect 18371 42177 18383 42211
rect 18325 42171 18383 42177
rect 18473 42211 18552 42217
rect 18473 42177 18485 42211
rect 18519 42180 18552 42211
rect 18601 42211 18659 42217
rect 18519 42177 18531 42180
rect 18473 42171 18531 42177
rect 18601 42177 18613 42211
rect 18647 42177 18659 42211
rect 18601 42171 18659 42177
rect 18693 42211 18751 42217
rect 18693 42177 18705 42211
rect 18739 42177 18751 42211
rect 18693 42171 18751 42177
rect 17310 42100 17316 42152
rect 17368 42100 17374 42152
rect 17420 42140 17448 42168
rect 18616 42140 18644 42171
rect 17420 42112 18644 42140
rect 18708 42140 18736 42171
rect 18782 42168 18788 42220
rect 18840 42217 18846 42220
rect 19076 42217 19104 42248
rect 18840 42208 18848 42217
rect 19061 42211 19119 42217
rect 18840 42180 18885 42208
rect 18840 42171 18848 42180
rect 19061 42177 19073 42211
rect 19107 42177 19119 42211
rect 20622 42208 20628 42220
rect 20470 42180 20628 42208
rect 19061 42171 19119 42177
rect 18840 42168 18846 42171
rect 20622 42168 20628 42180
rect 20680 42168 20686 42220
rect 21836 42217 21864 42316
rect 25130 42304 25136 42356
rect 25188 42344 25194 42356
rect 25188 42316 25360 42344
rect 25188 42304 25194 42316
rect 22370 42236 22376 42288
rect 22428 42276 22434 42288
rect 25332 42285 25360 42316
rect 27154 42304 27160 42356
rect 27212 42304 27218 42356
rect 34054 42344 34060 42356
rect 33704 42316 34060 42344
rect 25317 42279 25375 42285
rect 22428 42248 22586 42276
rect 22428 42236 22434 42248
rect 25317 42245 25329 42279
rect 25363 42245 25375 42279
rect 27172 42276 27200 42304
rect 27430 42276 27436 42288
rect 26542 42248 27436 42276
rect 25317 42239 25375 42245
rect 27430 42236 27436 42248
rect 27488 42236 27494 42288
rect 33704 42285 33732 42316
rect 34054 42304 34060 42316
rect 34112 42304 34118 42356
rect 35526 42344 35532 42356
rect 34900 42316 35532 42344
rect 33689 42279 33747 42285
rect 33689 42245 33701 42279
rect 33735 42245 33747 42279
rect 34790 42276 34796 42288
rect 33689 42239 33747 42245
rect 33980 42248 34796 42276
rect 21821 42211 21879 42217
rect 21821 42177 21833 42211
rect 21867 42177 21879 42211
rect 21821 42171 21879 42177
rect 26973 42211 27031 42217
rect 26973 42177 26985 42211
rect 27019 42177 27031 42211
rect 26973 42171 27031 42177
rect 18708 42112 19196 42140
rect 18138 42072 18144 42084
rect 14608 42044 18144 42072
rect 14608 42032 14614 42044
rect 18138 42032 18144 42044
rect 18196 42032 18202 42084
rect 13998 42004 14004 42016
rect 13096 41976 14004 42004
rect 12032 41964 12038 41976
rect 13998 41964 14004 41976
rect 14056 41964 14062 42016
rect 14476 42004 14504 42032
rect 17954 42004 17960 42016
rect 14476 41976 17960 42004
rect 17954 41964 17960 41976
rect 18012 41964 18018 42016
rect 18966 41964 18972 42016
rect 19024 41964 19030 42016
rect 19168 42004 19196 42112
rect 19334 42100 19340 42152
rect 19392 42100 19398 42152
rect 21453 42143 21511 42149
rect 21453 42140 21465 42143
rect 20824 42112 21465 42140
rect 20824 42013 20852 42112
rect 21453 42109 21465 42112
rect 21499 42109 21511 42143
rect 21453 42103 21511 42109
rect 22094 42100 22100 42152
rect 22152 42100 22158 42152
rect 24394 42100 24400 42152
rect 24452 42140 24458 42152
rect 25041 42143 25099 42149
rect 25041 42140 25053 42143
rect 24452 42112 25053 42140
rect 24452 42100 24458 42112
rect 25041 42109 25053 42112
rect 25087 42109 25099 42143
rect 25041 42103 25099 42109
rect 26878 42100 26884 42152
rect 26936 42140 26942 42152
rect 26988 42140 27016 42171
rect 27338 42168 27344 42220
rect 27396 42168 27402 42220
rect 32582 42168 32588 42220
rect 32640 42168 32646 42220
rect 33980 42217 34008 42248
rect 34790 42236 34796 42248
rect 34848 42236 34854 42288
rect 33965 42211 34023 42217
rect 33965 42177 33977 42211
rect 34011 42177 34023 42211
rect 33965 42171 34023 42177
rect 34609 42211 34667 42217
rect 34609 42177 34621 42211
rect 34655 42208 34667 42211
rect 34900 42208 34928 42316
rect 35526 42304 35532 42316
rect 35584 42304 35590 42356
rect 38838 42304 38844 42356
rect 38896 42304 38902 42356
rect 40310 42344 40316 42356
rect 40144 42316 40316 42344
rect 35069 42279 35127 42285
rect 35069 42245 35081 42279
rect 35115 42276 35127 42279
rect 35115 42248 35756 42276
rect 35115 42245 35127 42248
rect 35069 42239 35127 42245
rect 35728 42220 35756 42248
rect 36170 42236 36176 42288
rect 36228 42276 36234 42288
rect 36693 42279 36751 42285
rect 36693 42276 36705 42279
rect 36228 42248 36705 42276
rect 36228 42236 36234 42248
rect 36693 42245 36705 42248
rect 36739 42245 36751 42279
rect 36693 42239 36751 42245
rect 36906 42236 36912 42288
rect 36964 42236 36970 42288
rect 40144 42285 40172 42316
rect 40310 42304 40316 42316
rect 40368 42304 40374 42356
rect 42245 42347 42303 42353
rect 42245 42313 42257 42347
rect 42291 42313 42303 42347
rect 42245 42307 42303 42313
rect 40129 42279 40187 42285
rect 40129 42245 40141 42279
rect 40175 42245 40187 42279
rect 40129 42239 40187 42245
rect 40586 42236 40592 42288
rect 40644 42236 40650 42288
rect 42260 42276 42288 42307
rect 42705 42279 42763 42285
rect 42705 42276 42717 42279
rect 42260 42248 42717 42276
rect 42705 42245 42717 42248
rect 42751 42245 42763 42279
rect 42705 42239 42763 42245
rect 34655 42180 34928 42208
rect 35253 42211 35311 42217
rect 34655 42177 34667 42180
rect 34609 42171 34667 42177
rect 35253 42177 35265 42211
rect 35299 42177 35311 42211
rect 35253 42171 35311 42177
rect 26936 42112 27568 42140
rect 26936 42100 26942 42112
rect 27540 42081 27568 42112
rect 31726 42112 33916 42140
rect 27525 42075 27583 42081
rect 27525 42041 27537 42075
rect 27571 42072 27583 42075
rect 31726 42072 31754 42112
rect 27571 42044 31754 42072
rect 33888 42072 33916 42112
rect 34698 42100 34704 42152
rect 34756 42100 34762 42152
rect 34974 42100 34980 42152
rect 35032 42100 35038 42152
rect 35268 42072 35296 42171
rect 35710 42168 35716 42220
rect 35768 42208 35774 42220
rect 35768 42180 36860 42208
rect 35768 42168 35774 42180
rect 35526 42100 35532 42152
rect 35584 42140 35590 42152
rect 35805 42143 35863 42149
rect 35805 42140 35817 42143
rect 35584 42112 35817 42140
rect 35584 42100 35590 42112
rect 35805 42109 35817 42112
rect 35851 42109 35863 42143
rect 35805 42103 35863 42109
rect 33888 42044 35296 42072
rect 27571 42041 27583 42044
rect 27525 42035 27583 42041
rect 35618 42032 35624 42084
rect 35676 42072 35682 42084
rect 35676 42044 36768 42072
rect 35676 42032 35682 42044
rect 36740 42016 36768 42044
rect 20809 42007 20867 42013
rect 20809 42004 20821 42007
rect 19168 41976 20821 42004
rect 20809 41973 20821 41976
rect 20855 41973 20867 42007
rect 20809 41967 20867 41973
rect 20898 41964 20904 42016
rect 20956 41964 20962 42016
rect 23566 41964 23572 42016
rect 23624 41964 23630 42016
rect 26789 42007 26847 42013
rect 26789 41973 26801 42007
rect 26835 42004 26847 42007
rect 27062 42004 27068 42016
rect 26835 41976 27068 42004
rect 26835 41973 26847 41976
rect 26789 41967 26847 41973
rect 27062 41964 27068 41976
rect 27120 41964 27126 42016
rect 30926 41964 30932 42016
rect 30984 42004 30990 42016
rect 32217 42007 32275 42013
rect 32217 42004 32229 42007
rect 30984 41976 32229 42004
rect 30984 41964 30990 41976
rect 32217 41973 32229 41976
rect 32263 41973 32275 42007
rect 32217 41967 32275 41973
rect 36446 41964 36452 42016
rect 36504 41964 36510 42016
rect 36538 41964 36544 42016
rect 36596 41964 36602 42016
rect 36722 41964 36728 42016
rect 36780 41964 36786 42016
rect 36832 42004 36860 42180
rect 38838 42168 38844 42220
rect 38896 42168 38902 42220
rect 39025 42211 39083 42217
rect 39025 42177 39037 42211
rect 39071 42208 39083 42211
rect 39390 42208 39396 42220
rect 39071 42180 39396 42208
rect 39071 42177 39083 42180
rect 39025 42171 39083 42177
rect 39390 42168 39396 42180
rect 39448 42168 39454 42220
rect 42061 42211 42119 42217
rect 42061 42177 42073 42211
rect 42107 42208 42119 42211
rect 42242 42208 42248 42220
rect 42107 42180 42248 42208
rect 42107 42177 42119 42180
rect 42061 42171 42119 42177
rect 42242 42168 42248 42180
rect 42300 42168 42306 42220
rect 38470 42100 38476 42152
rect 38528 42140 38534 42152
rect 39853 42143 39911 42149
rect 39853 42140 39865 42143
rect 38528 42112 39865 42140
rect 38528 42100 38534 42112
rect 39853 42109 39865 42112
rect 39899 42109 39911 42143
rect 39853 42103 39911 42109
rect 40586 42100 40592 42152
rect 40644 42140 40650 42152
rect 41138 42140 41144 42152
rect 40644 42112 41144 42140
rect 40644 42100 40650 42112
rect 41138 42100 41144 42112
rect 41196 42140 41202 42152
rect 41196 42112 41414 42140
rect 41196 42100 41202 42112
rect 41386 42072 41414 42112
rect 42426 42100 42432 42152
rect 42484 42100 42490 42152
rect 43824 42140 43852 42194
rect 42536 42112 43852 42140
rect 42536 42072 42564 42112
rect 41386 42044 42564 42072
rect 41230 42004 41236 42016
rect 36832 41976 41236 42004
rect 41230 41964 41236 41976
rect 41288 41964 41294 42016
rect 41598 41964 41604 42016
rect 41656 42004 41662 42016
rect 42334 42004 42340 42016
rect 41656 41976 42340 42004
rect 41656 41964 41662 41976
rect 42334 41964 42340 41976
rect 42392 41964 42398 42016
rect 44174 41964 44180 42016
rect 44232 41964 44238 42016
rect 1104 41914 44620 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 44620 41914
rect 1104 41840 44620 41862
rect 7374 41760 7380 41812
rect 7432 41800 7438 41812
rect 7745 41803 7803 41809
rect 7745 41800 7757 41803
rect 7432 41772 7757 41800
rect 7432 41760 7438 41772
rect 7745 41769 7757 41772
rect 7791 41769 7803 41803
rect 8938 41800 8944 41812
rect 7745 41763 7803 41769
rect 8404 41772 8944 41800
rect 8404 41605 8432 41772
rect 8938 41760 8944 41772
rect 8996 41760 9002 41812
rect 10134 41760 10140 41812
rect 10192 41760 10198 41812
rect 11974 41760 11980 41812
rect 12032 41760 12038 41812
rect 12158 41760 12164 41812
rect 12216 41800 12222 41812
rect 12216 41772 12434 41800
rect 12216 41760 12222 41772
rect 9600 41704 10364 41732
rect 9600 41676 9628 41704
rect 8665 41667 8723 41673
rect 8665 41633 8677 41667
rect 8711 41664 8723 41667
rect 9582 41664 9588 41676
rect 8711 41636 9588 41664
rect 8711 41633 8723 41636
rect 8665 41627 8723 41633
rect 9582 41624 9588 41636
rect 9640 41624 9646 41676
rect 9858 41624 9864 41676
rect 9916 41664 9922 41676
rect 10229 41667 10287 41673
rect 10229 41664 10241 41667
rect 9916 41636 10241 41664
rect 9916 41624 9922 41636
rect 10229 41633 10241 41636
rect 10275 41633 10287 41667
rect 10336 41664 10364 41704
rect 12176 41664 12204 41760
rect 12406 41732 12434 41772
rect 13354 41760 13360 41812
rect 13412 41800 13418 41812
rect 14093 41803 14151 41809
rect 14093 41800 14105 41803
rect 13412 41772 14105 41800
rect 13412 41760 13418 41772
rect 14093 41769 14105 41772
rect 14139 41769 14151 41803
rect 14093 41763 14151 41769
rect 15562 41760 15568 41812
rect 15620 41760 15626 41812
rect 17310 41760 17316 41812
rect 17368 41760 17374 41812
rect 17957 41803 18015 41809
rect 17957 41769 17969 41803
rect 18003 41800 18015 41803
rect 18414 41800 18420 41812
rect 18003 41772 18420 41800
rect 18003 41769 18015 41772
rect 17957 41763 18015 41769
rect 18414 41760 18420 41772
rect 18472 41760 18478 41812
rect 18966 41760 18972 41812
rect 19024 41760 19030 41812
rect 19334 41760 19340 41812
rect 19392 41800 19398 41812
rect 19889 41803 19947 41809
rect 19889 41800 19901 41803
rect 19392 41772 19901 41800
rect 19392 41760 19398 41772
rect 19889 41769 19901 41772
rect 19935 41769 19947 41803
rect 19889 41763 19947 41769
rect 20898 41760 20904 41812
rect 20956 41760 20962 41812
rect 21453 41803 21511 41809
rect 21453 41769 21465 41803
rect 21499 41800 21511 41803
rect 22094 41800 22100 41812
rect 21499 41772 22100 41800
rect 21499 41769 21511 41772
rect 21453 41763 21511 41769
rect 22094 41760 22100 41772
rect 22152 41760 22158 41812
rect 23566 41760 23572 41812
rect 23624 41760 23630 41812
rect 31202 41760 31208 41812
rect 31260 41800 31266 41812
rect 31297 41803 31355 41809
rect 31297 41800 31309 41803
rect 31260 41772 31309 41800
rect 31260 41760 31266 41772
rect 31297 41769 31309 41772
rect 31343 41769 31355 41803
rect 31297 41763 31355 41769
rect 13633 41735 13691 41741
rect 12406 41704 13584 41732
rect 10336 41636 12204 41664
rect 10229 41627 10287 41633
rect 12894 41624 12900 41676
rect 12952 41664 12958 41676
rect 12952 41636 13216 41664
rect 12952 41624 12958 41636
rect 7929 41599 7987 41605
rect 7929 41565 7941 41599
rect 7975 41596 7987 41599
rect 8389 41599 8447 41605
rect 7975 41568 8064 41596
rect 7975 41565 7987 41568
rect 7929 41559 7987 41565
rect 8036 41469 8064 41568
rect 8389 41565 8401 41599
rect 8435 41565 8447 41599
rect 8389 41559 8447 41565
rect 10042 41556 10048 41608
rect 10100 41556 10106 41608
rect 11790 41596 11796 41608
rect 11638 41568 11796 41596
rect 11790 41556 11796 41568
rect 11848 41556 11854 41608
rect 11882 41556 11888 41608
rect 11940 41596 11946 41608
rect 12253 41599 12311 41605
rect 12253 41596 12265 41599
rect 11940 41568 12265 41596
rect 11940 41556 11946 41568
rect 12253 41565 12265 41568
rect 12299 41565 12311 41599
rect 12253 41559 12311 41565
rect 12618 41556 12624 41608
rect 12676 41596 12682 41608
rect 12989 41599 13047 41605
rect 12989 41596 13001 41599
rect 12676 41568 13001 41596
rect 12676 41556 12682 41568
rect 12989 41565 13001 41568
rect 13035 41565 13047 41599
rect 12989 41559 13047 41565
rect 13082 41599 13140 41605
rect 13082 41565 13094 41599
rect 13128 41565 13140 41599
rect 13188 41596 13216 41636
rect 13454 41599 13512 41605
rect 13454 41596 13466 41599
rect 13188 41568 13466 41596
rect 13082 41559 13140 41565
rect 13454 41565 13466 41568
rect 13500 41565 13512 41599
rect 13556 41596 13584 41704
rect 13633 41701 13645 41735
rect 13679 41701 13691 41735
rect 13633 41695 13691 41701
rect 13648 41664 13676 41695
rect 14645 41667 14703 41673
rect 14645 41664 14657 41667
rect 13648 41636 14657 41664
rect 14645 41633 14657 41636
rect 14691 41633 14703 41667
rect 15580 41664 15608 41760
rect 18782 41664 18788 41676
rect 15580 41636 18788 41664
rect 14645 41627 14703 41633
rect 15470 41596 15476 41608
rect 13556 41568 15476 41596
rect 13454 41559 13512 41565
rect 8021 41463 8079 41469
rect 8021 41429 8033 41463
rect 8067 41429 8079 41463
rect 8021 41423 8079 41429
rect 8478 41420 8484 41472
rect 8536 41420 8542 41472
rect 9674 41420 9680 41472
rect 9732 41420 9738 41472
rect 9769 41463 9827 41469
rect 9769 41429 9781 41463
rect 9815 41460 9827 41463
rect 10060 41460 10088 41556
rect 10502 41488 10508 41540
rect 10560 41488 10566 41540
rect 12526 41488 12532 41540
rect 12584 41488 12590 41540
rect 12897 41531 12955 41537
rect 12897 41497 12909 41531
rect 12943 41528 12955 41531
rect 13096 41528 13124 41559
rect 15470 41556 15476 41568
rect 15528 41556 15534 41608
rect 16666 41556 16672 41608
rect 16724 41556 16730 41608
rect 16758 41556 16764 41608
rect 16816 41596 16822 41608
rect 16816 41568 16861 41596
rect 16816 41556 16822 41568
rect 17034 41556 17040 41608
rect 17092 41556 17098 41608
rect 17144 41605 17172 41636
rect 18782 41624 18788 41636
rect 18840 41624 18846 41676
rect 18984 41664 19012 41760
rect 19245 41667 19303 41673
rect 19245 41664 19257 41667
rect 18984 41636 19257 41664
rect 19245 41633 19257 41636
rect 19291 41633 19303 41667
rect 19245 41627 19303 41633
rect 17134 41599 17192 41605
rect 17134 41565 17146 41599
rect 17180 41565 17192 41599
rect 17134 41559 17192 41565
rect 17586 41556 17592 41608
rect 17644 41556 17650 41608
rect 17773 41599 17831 41605
rect 17773 41565 17785 41599
rect 17819 41565 17831 41599
rect 17773 41559 17831 41565
rect 12943 41500 13124 41528
rect 12943 41497 12955 41500
rect 12897 41491 12955 41497
rect 13262 41488 13268 41540
rect 13320 41488 13326 41540
rect 13357 41531 13415 41537
rect 13357 41497 13369 41531
rect 13403 41528 13415 41531
rect 15010 41528 15016 41540
rect 13403 41500 15016 41528
rect 13403 41497 13415 41500
rect 13357 41491 13415 41497
rect 15010 41488 15016 41500
rect 15068 41488 15074 41540
rect 16945 41531 17003 41537
rect 16945 41497 16957 41531
rect 16991 41497 17003 41531
rect 17788 41528 17816 41559
rect 18138 41528 18144 41540
rect 17788 41500 18144 41528
rect 16945 41491 17003 41497
rect 9815 41432 10088 41460
rect 12544 41460 12572 41488
rect 13280 41460 13308 41488
rect 16960 41460 16988 41491
rect 18138 41488 18144 41500
rect 18196 41488 18202 41540
rect 18800 41528 18828 41624
rect 20806 41556 20812 41608
rect 20864 41556 20870 41608
rect 20916 41605 20944 41760
rect 23584 41664 23612 41760
rect 24949 41667 25007 41673
rect 24949 41664 24961 41667
rect 23584 41636 24961 41664
rect 24949 41633 24961 41636
rect 24995 41633 25007 41667
rect 24949 41627 25007 41633
rect 20902 41599 20960 41605
rect 20902 41565 20914 41599
rect 20948 41565 20960 41599
rect 21274 41599 21332 41605
rect 21274 41596 21286 41599
rect 20902 41559 20960 41565
rect 21008 41568 21286 41596
rect 21008 41528 21036 41568
rect 21274 41565 21286 41568
rect 21320 41596 21332 41599
rect 24210 41596 24216 41608
rect 21320 41568 24216 41596
rect 21320 41565 21332 41568
rect 21274 41559 21332 41565
rect 24210 41556 24216 41568
rect 24268 41556 24274 41608
rect 18800 41500 21036 41528
rect 21085 41531 21143 41537
rect 21085 41497 21097 41531
rect 21131 41497 21143 41531
rect 21085 41491 21143 41497
rect 21177 41531 21235 41537
rect 21177 41497 21189 41531
rect 21223 41528 21235 41531
rect 23566 41528 23572 41540
rect 21223 41500 23572 41528
rect 21223 41497 21235 41500
rect 21177 41491 21235 41497
rect 17310 41460 17316 41472
rect 12544 41432 17316 41460
rect 9815 41429 9827 41432
rect 9769 41423 9827 41429
rect 17310 41420 17316 41432
rect 17368 41420 17374 41472
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 19426 41460 19432 41472
rect 18012 41432 19432 41460
rect 18012 41420 18018 41432
rect 19426 41420 19432 41432
rect 19484 41420 19490 41472
rect 21100 41460 21128 41491
rect 23566 41488 23572 41500
rect 23624 41528 23630 41540
rect 24397 41531 24455 41537
rect 24397 41528 24409 41531
rect 23624 41500 24409 41528
rect 23624 41488 23630 41500
rect 24397 41497 24409 41500
rect 24443 41497 24455 41531
rect 31312 41528 31340 41763
rect 34698 41760 34704 41812
rect 34756 41800 34762 41812
rect 35161 41803 35219 41809
rect 35161 41800 35173 41803
rect 34756 41772 35173 41800
rect 34756 41760 34762 41772
rect 35161 41769 35173 41772
rect 35207 41769 35219 41803
rect 35161 41763 35219 41769
rect 35342 41760 35348 41812
rect 35400 41800 35406 41812
rect 36078 41800 36084 41812
rect 35400 41772 36084 41800
rect 35400 41760 35406 41772
rect 36078 41760 36084 41772
rect 36136 41800 36142 41812
rect 36725 41803 36783 41809
rect 36725 41800 36737 41803
rect 36136 41772 36737 41800
rect 36136 41760 36142 41772
rect 36725 41769 36737 41772
rect 36771 41800 36783 41803
rect 37274 41800 37280 41812
rect 36771 41772 37280 41800
rect 36771 41769 36783 41772
rect 36725 41763 36783 41769
rect 37274 41760 37280 41772
rect 37332 41800 37338 41812
rect 38470 41800 38476 41812
rect 37332 41772 38476 41800
rect 37332 41760 37338 41772
rect 38470 41760 38476 41772
rect 38528 41760 38534 41812
rect 38930 41760 38936 41812
rect 38988 41800 38994 41812
rect 39301 41803 39359 41809
rect 39301 41800 39313 41803
rect 38988 41772 39313 41800
rect 38988 41760 38994 41772
rect 39301 41769 39313 41772
rect 39347 41769 39359 41803
rect 40862 41800 40868 41812
rect 39301 41763 39359 41769
rect 40236 41772 40868 41800
rect 32784 41636 38240 41664
rect 32030 41596 32036 41608
rect 31726 41568 32036 41596
rect 31726 41528 31754 41568
rect 32030 41556 32036 41568
rect 32088 41596 32094 41608
rect 32677 41599 32735 41605
rect 32677 41596 32689 41599
rect 32088 41568 32689 41596
rect 32088 41556 32094 41568
rect 32677 41565 32689 41568
rect 32723 41565 32735 41599
rect 32677 41559 32735 41565
rect 31312 41500 31754 41528
rect 32585 41531 32643 41537
rect 24397 41491 24455 41497
rect 32585 41497 32597 41531
rect 32631 41528 32643 41531
rect 32784 41528 32812 41636
rect 38212 41608 38240 41636
rect 33045 41599 33103 41605
rect 33045 41565 33057 41599
rect 33091 41596 33103 41599
rect 33134 41596 33140 41608
rect 33091 41568 33140 41596
rect 33091 41565 33103 41568
rect 33045 41559 33103 41565
rect 33134 41556 33140 41568
rect 33192 41556 33198 41608
rect 34514 41605 34520 41608
rect 34471 41599 34520 41605
rect 34471 41596 34483 41599
rect 34427 41568 34483 41596
rect 34471 41565 34483 41568
rect 34517 41565 34520 41599
rect 34471 41559 34520 41565
rect 34514 41556 34520 41559
rect 34572 41596 34578 41608
rect 35345 41599 35403 41605
rect 35345 41596 35357 41599
rect 34572 41568 35357 41596
rect 34572 41556 34578 41568
rect 35345 41565 35357 41568
rect 35391 41596 35403 41599
rect 35618 41596 35624 41608
rect 35391 41568 35624 41596
rect 35391 41565 35403 41568
rect 35345 41559 35403 41565
rect 35618 41556 35624 41568
rect 35676 41556 35682 41608
rect 36078 41556 36084 41608
rect 36136 41556 36142 41608
rect 36173 41599 36231 41605
rect 36173 41565 36185 41599
rect 36219 41565 36231 41599
rect 36173 41559 36231 41565
rect 36357 41599 36415 41605
rect 36357 41565 36369 41599
rect 36403 41596 36415 41599
rect 36446 41596 36452 41608
rect 36403 41568 36452 41596
rect 36403 41565 36415 41568
rect 36357 41559 36415 41565
rect 34882 41528 34888 41540
rect 32631 41500 32812 41528
rect 34086 41500 34888 41528
rect 32631 41497 32643 41500
rect 32585 41491 32643 41497
rect 34882 41488 34888 41500
rect 34940 41488 34946 41540
rect 35894 41488 35900 41540
rect 35952 41528 35958 41540
rect 36188 41528 36216 41559
rect 36446 41556 36452 41568
rect 36504 41556 36510 41608
rect 36538 41556 36544 41608
rect 36596 41556 36602 41608
rect 38194 41556 38200 41608
rect 38252 41556 38258 41608
rect 39942 41556 39948 41608
rect 40000 41596 40006 41608
rect 40236 41605 40264 41772
rect 40862 41760 40868 41772
rect 40920 41760 40926 41812
rect 41230 41760 41236 41812
rect 41288 41800 41294 41812
rect 41785 41803 41843 41809
rect 41288 41772 41736 41800
rect 41288 41760 41294 41772
rect 40954 41732 40960 41744
rect 40788 41704 40960 41732
rect 40681 41667 40739 41673
rect 40681 41633 40693 41667
rect 40727 41664 40739 41667
rect 40788 41664 40816 41704
rect 40954 41692 40960 41704
rect 41012 41692 41018 41744
rect 40727 41636 40816 41664
rect 41141 41667 41199 41673
rect 40727 41633 40739 41636
rect 40681 41627 40739 41633
rect 41141 41633 41153 41667
rect 41187 41664 41199 41667
rect 41598 41664 41604 41676
rect 41187 41636 41604 41664
rect 41187 41633 41199 41636
rect 41141 41627 41199 41633
rect 41598 41624 41604 41636
rect 41656 41624 41662 41676
rect 41708 41664 41736 41772
rect 41785 41769 41797 41803
rect 41831 41800 41843 41803
rect 42061 41803 42119 41809
rect 42061 41800 42073 41803
rect 41831 41772 42073 41800
rect 41831 41769 41843 41772
rect 41785 41763 41843 41769
rect 42061 41769 42073 41772
rect 42107 41769 42119 41803
rect 42061 41763 42119 41769
rect 42242 41760 42248 41812
rect 42300 41760 42306 41812
rect 41708 41636 42012 41664
rect 40221 41599 40279 41605
rect 40221 41596 40233 41599
rect 40000 41568 40233 41596
rect 40000 41556 40006 41568
rect 40221 41565 40233 41568
rect 40267 41565 40279 41599
rect 40221 41559 40279 41565
rect 40862 41556 40868 41608
rect 40920 41556 40926 41608
rect 40954 41556 40960 41608
rect 41012 41556 41018 41608
rect 41049 41599 41107 41605
rect 41049 41565 41061 41599
rect 41095 41565 41107 41599
rect 41049 41559 41107 41565
rect 41156 41568 41920 41596
rect 36556 41528 36584 41556
rect 35952 41500 36584 41528
rect 35952 41488 35958 41500
rect 39482 41488 39488 41540
rect 39540 41528 39546 41540
rect 39540 41500 40172 41528
rect 39540 41488 39546 41500
rect 22278 41460 22284 41472
rect 21100 41432 22284 41460
rect 22278 41420 22284 41432
rect 22336 41420 22342 41472
rect 35434 41420 35440 41472
rect 35492 41420 35498 41472
rect 36262 41420 36268 41472
rect 36320 41420 36326 41472
rect 39114 41420 39120 41472
rect 39172 41420 39178 41472
rect 39298 41469 39304 41472
rect 39285 41463 39304 41469
rect 39285 41429 39297 41463
rect 39285 41423 39304 41429
rect 39298 41420 39304 41423
rect 39356 41420 39362 41472
rect 39390 41420 39396 41472
rect 39448 41460 39454 41472
rect 39942 41460 39948 41472
rect 39448 41432 39948 41460
rect 39448 41420 39454 41432
rect 39942 41420 39948 41432
rect 40000 41420 40006 41472
rect 40034 41420 40040 41472
rect 40092 41420 40098 41472
rect 40144 41460 40172 41500
rect 40310 41488 40316 41540
rect 40368 41488 40374 41540
rect 40402 41488 40408 41540
rect 40460 41488 40466 41540
rect 40589 41531 40647 41537
rect 40589 41497 40601 41531
rect 40635 41528 40647 41531
rect 40678 41528 40684 41540
rect 40635 41500 40684 41528
rect 40635 41497 40647 41500
rect 40589 41491 40647 41497
rect 40678 41488 40684 41500
rect 40736 41528 40742 41540
rect 41064 41528 41092 41559
rect 40736 41500 41092 41528
rect 40736 41488 40742 41500
rect 41156 41460 41184 41568
rect 41322 41488 41328 41540
rect 41380 41528 41386 41540
rect 41417 41531 41475 41537
rect 41417 41528 41429 41531
rect 41380 41500 41429 41528
rect 41380 41488 41386 41500
rect 41417 41497 41429 41500
rect 41463 41497 41475 41531
rect 41417 41491 41475 41497
rect 41601 41531 41659 41537
rect 41601 41497 41613 41531
rect 41647 41528 41659 41531
rect 41782 41528 41788 41540
rect 41647 41500 41788 41528
rect 41647 41497 41659 41500
rect 41601 41491 41659 41497
rect 41782 41488 41788 41500
rect 41840 41488 41846 41540
rect 41892 41537 41920 41568
rect 41877 41531 41935 41537
rect 41877 41497 41889 41531
rect 41923 41497 41935 41531
rect 41984 41528 42012 41636
rect 42426 41624 42432 41676
rect 42484 41664 42490 41676
rect 42521 41667 42579 41673
rect 42521 41664 42533 41667
rect 42484 41636 42533 41664
rect 42484 41624 42490 41636
rect 42521 41633 42533 41636
rect 42567 41633 42579 41667
rect 42521 41627 42579 41633
rect 42797 41667 42855 41673
rect 42797 41633 42809 41667
rect 42843 41664 42855 41667
rect 43346 41664 43352 41676
rect 42843 41636 43352 41664
rect 42843 41633 42855 41636
rect 42797 41627 42855 41633
rect 43346 41624 43352 41636
rect 43404 41624 43410 41676
rect 43070 41528 43076 41540
rect 41984 41500 43076 41528
rect 41877 41491 41935 41497
rect 43070 41488 43076 41500
rect 43128 41528 43134 41540
rect 43128 41500 43286 41528
rect 43128 41488 43134 41500
rect 40144 41432 41184 41460
rect 42058 41420 42064 41472
rect 42116 41469 42122 41472
rect 42116 41463 42135 41469
rect 42123 41429 42135 41463
rect 42116 41423 42135 41429
rect 42116 41420 42122 41423
rect 44082 41420 44088 41472
rect 44140 41460 44146 41472
rect 44269 41463 44327 41469
rect 44269 41460 44281 41463
rect 44140 41432 44281 41460
rect 44140 41420 44146 41432
rect 44269 41429 44281 41432
rect 44315 41429 44327 41463
rect 44269 41423 44327 41429
rect 1104 41370 44620 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 44620 41370
rect 1104 41296 44620 41318
rect 10502 41216 10508 41268
rect 10560 41256 10566 41268
rect 10965 41259 11023 41265
rect 10965 41256 10977 41259
rect 10560 41228 10977 41256
rect 10560 41216 10566 41228
rect 10965 41225 10977 41228
rect 11011 41225 11023 41259
rect 10965 41219 11023 41225
rect 11882 41216 11888 41268
rect 11940 41216 11946 41268
rect 20806 41256 20812 41268
rect 19352 41228 20812 41256
rect 13357 41191 13415 41197
rect 10888 41160 12190 41188
rect 10888 41132 10916 41160
rect 13357 41157 13369 41191
rect 13403 41188 13415 41191
rect 13725 41191 13783 41197
rect 13725 41188 13737 41191
rect 13403 41160 13737 41188
rect 13403 41157 13415 41160
rect 13357 41151 13415 41157
rect 13725 41157 13737 41160
rect 13771 41157 13783 41191
rect 13725 41151 13783 41157
rect 15657 41191 15715 41197
rect 15657 41157 15669 41191
rect 15703 41188 15715 41191
rect 16669 41191 16727 41197
rect 16669 41188 16681 41191
rect 15703 41160 16681 41188
rect 15703 41157 15715 41160
rect 15657 41151 15715 41157
rect 16669 41157 16681 41160
rect 16715 41157 16727 41191
rect 16669 41151 16727 41157
rect 9125 41123 9183 41129
rect 9125 41089 9137 41123
rect 9171 41089 9183 41123
rect 9125 41083 9183 41089
rect 9140 40984 9168 41083
rect 10870 41080 10876 41132
rect 10928 41080 10934 41132
rect 11149 41123 11207 41129
rect 11149 41089 11161 41123
rect 11195 41120 11207 41123
rect 11514 41120 11520 41132
rect 11195 41092 11520 41120
rect 11195 41089 11207 41092
rect 11149 41083 11207 41089
rect 11514 41080 11520 41092
rect 11572 41080 11578 41132
rect 16301 41123 16359 41129
rect 16301 41120 16313 41123
rect 16040 41092 16313 41120
rect 13633 41055 13691 41061
rect 13633 41021 13645 41055
rect 13679 41052 13691 41055
rect 13998 41052 14004 41064
rect 13679 41024 14004 41052
rect 13679 41021 13691 41024
rect 13633 41015 13691 41021
rect 13998 41012 14004 41024
rect 14056 41012 14062 41064
rect 14274 41012 14280 41064
rect 14332 41012 14338 41064
rect 15470 41012 15476 41064
rect 15528 41012 15534 41064
rect 15562 41012 15568 41064
rect 15620 41012 15626 41064
rect 16040 40993 16068 41092
rect 16301 41089 16313 41092
rect 16347 41089 16359 41123
rect 16301 41083 16359 41089
rect 17313 41123 17371 41129
rect 17313 41089 17325 41123
rect 17359 41120 17371 41123
rect 17586 41120 17592 41132
rect 17359 41092 17592 41120
rect 17359 41089 17371 41092
rect 17313 41083 17371 41089
rect 17586 41080 17592 41092
rect 17644 41080 17650 41132
rect 18138 41080 18144 41132
rect 18196 41080 18202 41132
rect 19352 41129 19380 41228
rect 20806 41216 20812 41228
rect 20864 41216 20870 41268
rect 33134 41216 33140 41268
rect 33192 41256 33198 41268
rect 33965 41259 34023 41265
rect 33965 41256 33977 41259
rect 33192 41228 33977 41256
rect 33192 41216 33198 41228
rect 33965 41225 33977 41228
rect 34011 41225 34023 41259
rect 33965 41219 34023 41225
rect 34793 41259 34851 41265
rect 34793 41225 34805 41259
rect 34839 41256 34851 41259
rect 34882 41256 34888 41268
rect 34839 41228 34888 41256
rect 34839 41225 34851 41228
rect 34793 41219 34851 41225
rect 34882 41216 34888 41228
rect 34940 41216 34946 41268
rect 35710 41256 35716 41268
rect 35084 41228 35716 41256
rect 19426 41148 19432 41200
rect 19484 41188 19490 41200
rect 21913 41191 21971 41197
rect 19484 41160 19656 41188
rect 19484 41148 19490 41160
rect 19628 41129 19656 41160
rect 21913 41157 21925 41191
rect 21959 41188 21971 41191
rect 22186 41188 22192 41200
rect 21959 41160 22192 41188
rect 21959 41157 21971 41160
rect 21913 41151 21971 41157
rect 22186 41148 22192 41160
rect 22244 41188 22250 41200
rect 35084 41197 35112 41228
rect 35710 41216 35716 41228
rect 35768 41216 35774 41268
rect 36262 41256 36268 41268
rect 35866 41228 36268 41256
rect 22373 41191 22431 41197
rect 22373 41188 22385 41191
rect 22244 41160 22385 41188
rect 22244 41148 22250 41160
rect 22373 41157 22385 41160
rect 22419 41157 22431 41191
rect 22373 41151 22431 41157
rect 35069 41191 35127 41197
rect 35069 41157 35081 41191
rect 35115 41157 35127 41191
rect 35069 41151 35127 41157
rect 35621 41191 35679 41197
rect 35621 41157 35633 41191
rect 35667 41188 35679 41191
rect 35866 41188 35894 41228
rect 36262 41216 36268 41228
rect 36320 41216 36326 41268
rect 37090 41216 37096 41268
rect 37148 41256 37154 41268
rect 37148 41228 38700 41256
rect 37148 41216 37154 41228
rect 37108 41188 37136 41216
rect 35667 41160 35894 41188
rect 36846 41160 37228 41188
rect 35667 41157 35679 41160
rect 35621 41151 35679 41157
rect 18325 41123 18383 41129
rect 18325 41089 18337 41123
rect 18371 41120 18383 41123
rect 19337 41123 19395 41129
rect 19337 41120 19349 41123
rect 18371 41092 19349 41120
rect 18371 41089 18383 41092
rect 18325 41083 18383 41089
rect 19337 41089 19349 41092
rect 19383 41089 19395 41123
rect 19337 41083 19395 41089
rect 19521 41123 19579 41129
rect 19521 41089 19533 41123
rect 19567 41089 19579 41123
rect 19521 41083 19579 41089
rect 19613 41123 19671 41129
rect 19613 41089 19625 41123
rect 19659 41120 19671 41123
rect 21821 41123 21879 41129
rect 21821 41120 21833 41123
rect 19659 41092 21833 41120
rect 19659 41089 19671 41092
rect 19613 41083 19671 41089
rect 21821 41089 21833 41092
rect 21867 41089 21879 41123
rect 21821 41083 21879 41089
rect 17954 41012 17960 41064
rect 18012 41012 18018 41064
rect 19536 41052 19564 41083
rect 19536 41024 19932 41052
rect 16025 40987 16083 40993
rect 9140 40956 12020 40984
rect 9858 40876 9864 40928
rect 9916 40916 9922 40928
rect 10413 40919 10471 40925
rect 10413 40916 10425 40919
rect 9916 40888 10425 40916
rect 9916 40876 9922 40888
rect 10413 40885 10425 40888
rect 10459 40885 10471 40919
rect 11992 40916 12020 40956
rect 16025 40953 16037 40987
rect 16071 40953 16083 40987
rect 16025 40947 16083 40953
rect 13722 40916 13728 40928
rect 11992 40888 13728 40916
rect 10413 40879 10471 40885
rect 13722 40876 13728 40888
rect 13780 40876 13786 40928
rect 16114 40876 16120 40928
rect 16172 40876 16178 40928
rect 19150 40876 19156 40928
rect 19208 40876 19214 40928
rect 19904 40925 19932 41024
rect 20438 41012 20444 41064
rect 20496 41012 20502 41064
rect 21836 41052 21864 41083
rect 22002 41080 22008 41132
rect 22060 41120 22066 41132
rect 22097 41123 22155 41129
rect 22097 41120 22109 41123
rect 22060 41092 22109 41120
rect 22060 41080 22066 41092
rect 22097 41089 22109 41092
rect 22143 41089 22155 41123
rect 22097 41083 22155 41089
rect 22281 41123 22339 41129
rect 22281 41089 22293 41123
rect 22327 41120 22339 41123
rect 23293 41123 23351 41129
rect 23293 41120 23305 41123
rect 22327 41092 23305 41120
rect 22327 41089 22339 41092
rect 22281 41083 22339 41089
rect 23293 41089 23305 41092
rect 23339 41089 23351 41123
rect 23293 41083 23351 41089
rect 34057 41123 34115 41129
rect 34057 41089 34069 41123
rect 34103 41120 34115 41123
rect 34606 41120 34612 41132
rect 34103 41092 34612 41120
rect 34103 41089 34115 41092
rect 34057 41083 34115 41089
rect 34606 41080 34612 41092
rect 34664 41080 34670 41132
rect 22554 41052 22560 41064
rect 21836 41024 22560 41052
rect 22554 41012 22560 41024
rect 22612 41012 22618 41064
rect 22922 41012 22928 41064
rect 22980 41012 22986 41064
rect 34790 41012 34796 41064
rect 34848 41052 34854 41064
rect 35342 41052 35348 41064
rect 34848 41024 35348 41052
rect 34848 41012 34854 41024
rect 35342 41012 35348 41024
rect 35400 41012 35406 41064
rect 36170 41012 36176 41064
rect 36228 41052 36234 41064
rect 37093 41055 37151 41061
rect 37093 41052 37105 41055
rect 36228 41024 37105 41052
rect 36228 41012 36234 41024
rect 37093 41021 37105 41024
rect 37139 41021 37151 41055
rect 37093 41015 37151 41021
rect 19889 40919 19947 40925
rect 19889 40885 19901 40919
rect 19935 40916 19947 40919
rect 20070 40916 20076 40928
rect 19935 40888 20076 40916
rect 19935 40885 19947 40888
rect 19889 40879 19947 40885
rect 20070 40876 20076 40888
rect 20128 40876 20134 40928
rect 23934 40876 23940 40928
rect 23992 40876 23998 40928
rect 34882 40876 34888 40928
rect 34940 40916 34946 40928
rect 36078 40916 36084 40928
rect 34940 40888 36084 40916
rect 34940 40876 34946 40888
rect 36078 40876 36084 40888
rect 36136 40916 36142 40928
rect 37200 40916 37228 41160
rect 37274 41080 37280 41132
rect 37332 41080 37338 41132
rect 37550 41012 37556 41064
rect 37608 41012 37614 41064
rect 38672 41052 38700 41228
rect 38838 41216 38844 41268
rect 38896 41256 38902 41268
rect 39025 41259 39083 41265
rect 39025 41256 39037 41259
rect 38896 41228 39037 41256
rect 38896 41216 38902 41228
rect 39025 41225 39037 41228
rect 39071 41225 39083 41259
rect 39025 41219 39083 41225
rect 39117 41259 39175 41265
rect 39117 41225 39129 41259
rect 39163 41256 39175 41259
rect 39298 41256 39304 41268
rect 39163 41228 39304 41256
rect 39163 41225 39175 41228
rect 39117 41219 39175 41225
rect 39040 41120 39068 41219
rect 39298 41216 39304 41228
rect 39356 41216 39362 41268
rect 40497 41259 40555 41265
rect 40497 41225 40509 41259
rect 40543 41256 40555 41259
rect 40770 41256 40776 41268
rect 40543 41228 40776 41256
rect 40543 41225 40555 41228
rect 40497 41219 40555 41225
rect 40770 41216 40776 41228
rect 40828 41216 40834 41268
rect 42058 41216 42064 41268
rect 42116 41216 42122 41268
rect 39390 41148 39396 41200
rect 39448 41188 39454 41200
rect 39485 41191 39543 41197
rect 39485 41188 39497 41191
rect 39448 41160 39497 41188
rect 39448 41148 39454 41160
rect 39485 41157 39497 41160
rect 39531 41157 39543 41191
rect 40402 41188 40408 41200
rect 39485 41151 39543 41157
rect 39960 41160 40408 41188
rect 39301 41123 39359 41129
rect 39301 41120 39313 41123
rect 39040 41092 39313 41120
rect 39301 41089 39313 41092
rect 39347 41120 39359 41123
rect 39960 41120 39988 41160
rect 40402 41148 40408 41160
rect 40460 41188 40466 41200
rect 40954 41188 40960 41200
rect 40460 41160 40960 41188
rect 40460 41148 40466 41160
rect 40954 41148 40960 41160
rect 41012 41148 41018 41200
rect 42702 41188 42708 41200
rect 41984 41160 42708 41188
rect 39347 41092 39988 41120
rect 39347 41089 39359 41092
rect 39301 41083 39359 41089
rect 40034 41080 40040 41132
rect 40092 41120 40098 41132
rect 41322 41120 41328 41132
rect 40092 41092 41328 41120
rect 40092 41080 40098 41092
rect 41322 41080 41328 41092
rect 41380 41120 41386 41132
rect 41984 41129 42012 41160
rect 42702 41148 42708 41160
rect 42760 41188 42766 41200
rect 44053 41191 44111 41197
rect 44053 41188 44065 41191
rect 42760 41160 44065 41188
rect 42760 41148 42766 41160
rect 44053 41157 44065 41160
rect 44099 41157 44111 41191
rect 44269 41191 44327 41197
rect 44269 41188 44281 41191
rect 44053 41151 44111 41157
rect 44192 41160 44281 41188
rect 44192 41132 44220 41160
rect 44269 41157 44281 41160
rect 44315 41157 44327 41191
rect 44269 41151 44327 41157
rect 41969 41123 42027 41129
rect 41969 41120 41981 41123
rect 41380 41092 41981 41120
rect 41380 41080 41386 41092
rect 41969 41089 41981 41092
rect 42015 41089 42027 41123
rect 41969 41083 42027 41089
rect 42153 41123 42211 41129
rect 42153 41089 42165 41123
rect 42199 41089 42211 41123
rect 42153 41083 42211 41089
rect 41138 41052 41144 41064
rect 38672 41024 41144 41052
rect 41138 41012 41144 41024
rect 41196 41012 41202 41064
rect 41782 41012 41788 41064
rect 41840 41052 41846 41064
rect 42168 41052 42196 41083
rect 42334 41080 42340 41132
rect 42392 41120 42398 41132
rect 42613 41123 42671 41129
rect 42613 41120 42625 41123
rect 42392 41092 42625 41120
rect 42392 41080 42398 41092
rect 42613 41089 42625 41092
rect 42659 41089 42671 41123
rect 43073 41123 43131 41129
rect 43073 41120 43085 41123
rect 42613 41083 42671 41089
rect 42720 41092 43085 41120
rect 42518 41052 42524 41064
rect 41840 41024 42524 41052
rect 41840 41012 41846 41024
rect 42518 41012 42524 41024
rect 42576 41052 42582 41064
rect 42720 41052 42748 41092
rect 43073 41089 43085 41092
rect 43119 41120 43131 41123
rect 44174 41120 44180 41132
rect 43119 41092 44180 41120
rect 43119 41089 43131 41092
rect 43073 41083 43131 41089
rect 44174 41080 44180 41092
rect 44232 41080 44238 41132
rect 42576 41024 42748 41052
rect 42797 41055 42855 41061
rect 42576 41012 42582 41024
rect 42797 41021 42809 41055
rect 42843 41052 42855 41055
rect 43809 41055 43867 41061
rect 43809 41052 43821 41055
rect 42843 41024 43821 41052
rect 42843 41021 42855 41024
rect 42797 41015 42855 41021
rect 43809 41021 43821 41024
rect 43855 41052 43867 41055
rect 43855 41024 44128 41052
rect 43855 41021 43867 41024
rect 43809 41015 43867 41021
rect 40405 40987 40463 40993
rect 40405 40953 40417 40987
rect 40451 40984 40463 40987
rect 41046 40984 41052 40996
rect 40451 40956 41052 40984
rect 40451 40953 40463 40956
rect 40405 40947 40463 40953
rect 41046 40944 41052 40956
rect 41104 40944 41110 40996
rect 44100 40928 44128 41024
rect 36136 40888 37228 40916
rect 36136 40876 36142 40888
rect 41874 40876 41880 40928
rect 41932 40916 41938 40928
rect 42429 40919 42487 40925
rect 42429 40916 42441 40919
rect 41932 40888 42441 40916
rect 41932 40876 41938 40888
rect 42429 40885 42441 40888
rect 42475 40885 42487 40919
rect 42429 40879 42487 40885
rect 42794 40876 42800 40928
rect 42852 40876 42858 40928
rect 43162 40876 43168 40928
rect 43220 40876 43226 40928
rect 43254 40876 43260 40928
rect 43312 40916 43318 40928
rect 43901 40919 43959 40925
rect 43901 40916 43913 40919
rect 43312 40888 43913 40916
rect 43312 40876 43318 40888
rect 43901 40885 43913 40888
rect 43947 40885 43959 40919
rect 43901 40879 43959 40885
rect 44082 40876 44088 40928
rect 44140 40876 44146 40928
rect 1104 40826 44620 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 44620 40826
rect 1104 40752 44620 40774
rect 12897 40715 12955 40721
rect 12897 40681 12909 40715
rect 12943 40712 12955 40715
rect 14274 40712 14280 40724
rect 12943 40684 14280 40712
rect 12943 40681 12955 40684
rect 12897 40675 12955 40681
rect 14274 40672 14280 40684
rect 14332 40672 14338 40724
rect 17037 40715 17095 40721
rect 17037 40681 17049 40715
rect 17083 40712 17095 40715
rect 17586 40712 17592 40724
rect 17083 40684 17592 40712
rect 17083 40681 17095 40684
rect 17037 40675 17095 40681
rect 17586 40672 17592 40684
rect 17644 40672 17650 40724
rect 17954 40672 17960 40724
rect 18012 40712 18018 40724
rect 18233 40715 18291 40721
rect 18233 40712 18245 40715
rect 18012 40684 18245 40712
rect 18012 40672 18018 40684
rect 18233 40681 18245 40684
rect 18279 40681 18291 40715
rect 18233 40675 18291 40681
rect 19150 40672 19156 40724
rect 19208 40672 19214 40724
rect 20612 40715 20670 40721
rect 20612 40681 20624 40715
rect 20658 40712 20670 40715
rect 21082 40712 21088 40724
rect 20658 40684 21088 40712
rect 20658 40681 20670 40684
rect 20612 40675 20670 40681
rect 21082 40672 21088 40684
rect 21140 40672 21146 40724
rect 22189 40715 22247 40721
rect 22189 40681 22201 40715
rect 22235 40712 22247 40715
rect 22922 40712 22928 40724
rect 22235 40684 22928 40712
rect 22235 40681 22247 40684
rect 22189 40675 22247 40681
rect 22922 40672 22928 40684
rect 22980 40672 22986 40724
rect 23934 40672 23940 40724
rect 23992 40672 23998 40724
rect 35253 40715 35311 40721
rect 35253 40681 35265 40715
rect 35299 40712 35311 40715
rect 35526 40712 35532 40724
rect 35299 40684 35532 40712
rect 35299 40681 35311 40684
rect 35253 40675 35311 40681
rect 35526 40672 35532 40684
rect 35584 40672 35590 40724
rect 36722 40672 36728 40724
rect 36780 40672 36786 40724
rect 37550 40672 37556 40724
rect 37608 40712 37614 40724
rect 38013 40715 38071 40721
rect 38013 40712 38025 40715
rect 37608 40684 38025 40712
rect 37608 40672 37614 40684
rect 38013 40681 38025 40684
rect 38059 40681 38071 40715
rect 38013 40675 38071 40681
rect 40402 40672 40408 40724
rect 40460 40672 40466 40724
rect 40589 40715 40647 40721
rect 40589 40681 40601 40715
rect 40635 40712 40647 40715
rect 40678 40712 40684 40724
rect 40635 40684 40684 40712
rect 40635 40681 40647 40684
rect 40589 40675 40647 40681
rect 40678 40672 40684 40684
rect 40736 40672 40742 40724
rect 42702 40672 42708 40724
rect 42760 40672 42766 40724
rect 43162 40672 43168 40724
rect 43220 40672 43226 40724
rect 43346 40672 43352 40724
rect 43404 40672 43410 40724
rect 9858 40576 9864 40588
rect 9140 40548 9864 40576
rect 8205 40511 8263 40517
rect 8205 40477 8217 40511
rect 8251 40477 8263 40511
rect 8205 40471 8263 40477
rect 8220 40440 8248 40471
rect 8478 40468 8484 40520
rect 8536 40508 8542 40520
rect 9140 40517 9168 40548
rect 9858 40536 9864 40548
rect 9916 40536 9922 40588
rect 10873 40579 10931 40585
rect 10873 40545 10885 40579
rect 10919 40576 10931 40579
rect 11701 40579 11759 40585
rect 11701 40576 11713 40579
rect 10919 40548 11713 40576
rect 10919 40545 10931 40548
rect 10873 40539 10931 40545
rect 11701 40545 11713 40548
rect 11747 40545 11759 40579
rect 12989 40579 13047 40585
rect 12989 40576 13001 40579
rect 11701 40539 11759 40545
rect 12636 40548 13001 40576
rect 9125 40511 9183 40517
rect 9125 40508 9137 40511
rect 8536 40480 9137 40508
rect 8536 40468 8542 40480
rect 9125 40477 9137 40480
rect 9171 40477 9183 40511
rect 9125 40471 9183 40477
rect 12250 40468 12256 40520
rect 12308 40468 12314 40520
rect 12401 40511 12459 40517
rect 12401 40477 12413 40511
rect 12447 40508 12459 40511
rect 12636 40508 12664 40548
rect 12989 40545 13001 40548
rect 13035 40545 13047 40579
rect 12989 40539 13047 40545
rect 15565 40579 15623 40585
rect 15565 40545 15577 40579
rect 15611 40576 15623 40579
rect 16114 40576 16120 40588
rect 15611 40548 16120 40576
rect 15611 40545 15623 40548
rect 15565 40539 15623 40545
rect 16114 40536 16120 40548
rect 16172 40536 16178 40588
rect 19168 40576 19196 40672
rect 23952 40644 23980 40672
rect 20272 40616 20484 40644
rect 19797 40579 19855 40585
rect 19797 40576 19809 40579
rect 19168 40548 19809 40576
rect 19797 40545 19809 40548
rect 19843 40545 19855 40579
rect 19797 40539 19855 40545
rect 12447 40480 12664 40508
rect 12759 40511 12817 40517
rect 12447 40477 12459 40480
rect 12401 40471 12459 40477
rect 12759 40477 12771 40511
rect 12805 40508 12817 40511
rect 12894 40508 12900 40520
rect 12805 40480 12900 40508
rect 12805 40477 12817 40480
rect 12759 40471 12817 40477
rect 12894 40468 12900 40480
rect 12952 40468 12958 40520
rect 13538 40468 13544 40520
rect 13596 40468 13602 40520
rect 15102 40468 15108 40520
rect 15160 40508 15166 40520
rect 15289 40511 15347 40517
rect 15289 40508 15301 40511
rect 15160 40480 15301 40508
rect 15160 40468 15166 40480
rect 15289 40477 15301 40480
rect 15335 40477 15347 40511
rect 15289 40471 15347 40477
rect 16666 40468 16672 40520
rect 16724 40508 16730 40520
rect 17402 40508 17408 40520
rect 16724 40480 17408 40508
rect 16724 40468 16730 40480
rect 17402 40468 17408 40480
rect 17460 40468 17466 40520
rect 17678 40468 17684 40520
rect 17736 40468 17742 40520
rect 17954 40468 17960 40520
rect 18012 40508 18018 40520
rect 18049 40511 18107 40517
rect 18049 40508 18061 40511
rect 18012 40480 18061 40508
rect 18012 40468 18018 40480
rect 18049 40477 18061 40480
rect 18095 40477 18107 40511
rect 18049 40471 18107 40477
rect 18782 40468 18788 40520
rect 18840 40468 18846 40520
rect 8220 40412 8616 40440
rect 8588 40384 8616 40412
rect 9398 40400 9404 40452
rect 9456 40400 9462 40452
rect 10870 40440 10876 40452
rect 10626 40412 10876 40440
rect 10870 40400 10876 40412
rect 10928 40400 10934 40452
rect 12526 40400 12532 40452
rect 12584 40400 12590 40452
rect 12621 40443 12679 40449
rect 12621 40409 12633 40443
rect 12667 40409 12679 40443
rect 16022 40440 16028 40452
rect 12621 40403 12679 40409
rect 15948 40412 16028 40440
rect 8570 40332 8576 40384
rect 8628 40332 8634 40384
rect 8754 40332 8760 40384
rect 8812 40332 8818 40384
rect 9674 40332 9680 40384
rect 9732 40372 9738 40384
rect 10778 40372 10784 40384
rect 9732 40344 10784 40372
rect 9732 40332 9738 40344
rect 10778 40332 10784 40344
rect 10836 40332 10842 40384
rect 10962 40332 10968 40384
rect 11020 40372 11026 40384
rect 11149 40375 11207 40381
rect 11149 40372 11161 40375
rect 11020 40344 11161 40372
rect 11020 40332 11026 40344
rect 11149 40341 11161 40344
rect 11195 40341 11207 40375
rect 11149 40335 11207 40341
rect 11882 40332 11888 40384
rect 11940 40372 11946 40384
rect 12636 40372 12664 40403
rect 11940 40344 12664 40372
rect 15948 40372 15976 40412
rect 16022 40400 16028 40412
rect 16080 40400 16086 40452
rect 16684 40372 16712 40468
rect 16850 40400 16856 40452
rect 16908 40440 16914 40452
rect 17129 40443 17187 40449
rect 17129 40440 17141 40443
rect 16908 40412 17141 40440
rect 16908 40400 16914 40412
rect 17129 40409 17141 40412
rect 17175 40409 17187 40443
rect 17129 40403 17187 40409
rect 20162 40400 20168 40452
rect 20220 40440 20226 40452
rect 20272 40440 20300 40616
rect 20346 40536 20352 40588
rect 20404 40536 20410 40588
rect 20456 40576 20484 40616
rect 23860 40616 23980 40644
rect 20622 40576 20628 40588
rect 20456 40548 20628 40576
rect 20622 40536 20628 40548
rect 20680 40576 20686 40588
rect 23661 40579 23719 40585
rect 20680 40548 22094 40576
rect 20680 40536 20686 40548
rect 22066 40508 22094 40548
rect 23661 40545 23673 40579
rect 23707 40576 23719 40579
rect 23860 40576 23888 40616
rect 24394 40604 24400 40656
rect 24452 40604 24458 40656
rect 35805 40647 35863 40653
rect 35805 40644 35817 40647
rect 34716 40616 35817 40644
rect 23707 40548 23888 40576
rect 23937 40579 23995 40585
rect 23707 40545 23719 40548
rect 23661 40539 23719 40545
rect 23937 40545 23949 40579
rect 23983 40576 23995 40579
rect 24412 40576 24440 40604
rect 23983 40548 24440 40576
rect 23983 40545 23995 40548
rect 23937 40539 23995 40545
rect 22370 40508 22376 40520
rect 22066 40480 22376 40508
rect 22370 40468 22376 40480
rect 22428 40508 22434 40520
rect 22428 40480 22586 40508
rect 22428 40468 22434 40480
rect 24118 40468 24124 40520
rect 24176 40508 24182 40520
rect 24397 40511 24455 40517
rect 24397 40508 24409 40511
rect 24176 40480 24409 40508
rect 24176 40468 24182 40480
rect 24397 40477 24409 40480
rect 24443 40477 24455 40511
rect 24397 40471 24455 40477
rect 34514 40468 34520 40520
rect 34572 40468 34578 40520
rect 34716 40517 34744 40616
rect 35805 40613 35817 40616
rect 35851 40613 35863 40647
rect 35805 40607 35863 40613
rect 35713 40579 35771 40585
rect 34900 40548 35572 40576
rect 34900 40517 34928 40548
rect 35544 40517 35572 40548
rect 35713 40545 35725 40579
rect 35759 40576 35771 40579
rect 40129 40579 40187 40585
rect 35759 40548 36032 40576
rect 35759 40545 35771 40548
rect 35713 40539 35771 40545
rect 34701 40511 34759 40517
rect 34701 40477 34713 40511
rect 34747 40477 34759 40511
rect 34701 40471 34759 40477
rect 34885 40511 34943 40517
rect 34885 40477 34897 40511
rect 34931 40477 34943 40511
rect 34885 40471 34943 40477
rect 34977 40511 35035 40517
rect 34977 40477 34989 40511
rect 35023 40477 35035 40511
rect 34977 40471 35035 40477
rect 35069 40511 35127 40517
rect 35069 40477 35081 40511
rect 35115 40508 35127 40511
rect 35529 40511 35587 40517
rect 35115 40480 35480 40508
rect 35115 40477 35127 40480
rect 35069 40471 35127 40477
rect 34532 40440 34560 40468
rect 34992 40440 35020 40471
rect 20220 40412 21114 40440
rect 34532 40412 35020 40440
rect 20220 40400 20226 40412
rect 35250 40400 35256 40452
rect 35308 40400 35314 40452
rect 35452 40440 35480 40480
rect 35529 40477 35541 40511
rect 35575 40508 35587 40511
rect 35894 40508 35900 40520
rect 35575 40480 35900 40508
rect 35575 40477 35587 40480
rect 35529 40471 35587 40477
rect 35894 40468 35900 40480
rect 35952 40468 35958 40520
rect 36004 40508 36032 40548
rect 40129 40545 40141 40579
rect 40175 40576 40187 40579
rect 40420 40576 40448 40672
rect 40175 40548 40448 40576
rect 40175 40545 40187 40548
rect 40129 40539 40187 40545
rect 36357 40511 36415 40517
rect 36357 40508 36369 40511
rect 36004 40480 36369 40508
rect 36004 40452 36032 40480
rect 36357 40477 36369 40480
rect 36403 40508 36415 40511
rect 36725 40511 36783 40517
rect 36725 40508 36737 40511
rect 36403 40480 36737 40508
rect 36403 40477 36415 40480
rect 36357 40471 36415 40477
rect 36725 40477 36737 40480
rect 36771 40477 36783 40511
rect 36725 40471 36783 40477
rect 36817 40511 36875 40517
rect 36817 40477 36829 40511
rect 36863 40508 36875 40511
rect 36906 40508 36912 40520
rect 36863 40480 36912 40508
rect 36863 40477 36875 40480
rect 36817 40471 36875 40477
rect 35452 40412 35894 40440
rect 15948 40344 16712 40372
rect 11940 40332 11946 40344
rect 17218 40332 17224 40384
rect 17276 40372 17282 40384
rect 17865 40375 17923 40381
rect 17865 40372 17877 40375
rect 17276 40344 17877 40372
rect 17276 40332 17282 40344
rect 17865 40341 17877 40344
rect 17911 40341 17923 40375
rect 17865 40335 17923 40341
rect 19058 40332 19064 40384
rect 19116 40372 19122 40384
rect 19245 40375 19303 40381
rect 19245 40372 19257 40375
rect 19116 40344 19257 40372
rect 19116 40332 19122 40344
rect 19245 40341 19257 40344
rect 19291 40341 19303 40375
rect 19245 40335 19303 40341
rect 22094 40332 22100 40384
rect 22152 40332 22158 40384
rect 24946 40332 24952 40384
rect 25004 40372 25010 40384
rect 25041 40375 25099 40381
rect 25041 40372 25053 40375
rect 25004 40344 25053 40372
rect 25004 40332 25010 40344
rect 25041 40341 25053 40344
rect 25087 40341 25099 40375
rect 25041 40335 25099 40341
rect 34606 40332 34612 40384
rect 34664 40372 34670 40384
rect 34793 40375 34851 40381
rect 34793 40372 34805 40375
rect 34664 40344 34805 40372
rect 34664 40332 34670 40344
rect 34793 40341 34805 40344
rect 34839 40341 34851 40375
rect 34793 40335 34851 40341
rect 35345 40375 35403 40381
rect 35345 40341 35357 40375
rect 35391 40372 35403 40375
rect 35526 40372 35532 40384
rect 35391 40344 35532 40372
rect 35391 40341 35403 40344
rect 35345 40335 35403 40341
rect 35526 40332 35532 40344
rect 35584 40332 35590 40384
rect 35866 40372 35894 40412
rect 35986 40400 35992 40452
rect 36044 40400 36050 40452
rect 36170 40400 36176 40452
rect 36228 40440 36234 40452
rect 36541 40443 36599 40449
rect 36541 40440 36553 40443
rect 36228 40412 36553 40440
rect 36228 40400 36234 40412
rect 36541 40409 36553 40412
rect 36587 40409 36599 40443
rect 36541 40403 36599 40409
rect 36832 40372 36860 40471
rect 36906 40468 36912 40480
rect 36964 40468 36970 40520
rect 38197 40511 38255 40517
rect 38197 40477 38209 40511
rect 38243 40508 38255 40511
rect 39114 40508 39120 40520
rect 38243 40480 39120 40508
rect 38243 40477 38255 40480
rect 38197 40471 38255 40477
rect 39114 40468 39120 40480
rect 39172 40468 39178 40520
rect 40221 40511 40279 40517
rect 40221 40477 40233 40511
rect 40267 40477 40279 40511
rect 40221 40471 40279 40477
rect 40236 40440 40264 40471
rect 40586 40468 40592 40520
rect 40644 40468 40650 40520
rect 42518 40468 42524 40520
rect 42576 40468 42582 40520
rect 42720 40517 42748 40672
rect 42981 40647 43039 40653
rect 42981 40644 42993 40647
rect 42904 40616 42993 40644
rect 42705 40511 42763 40517
rect 42705 40477 42717 40511
rect 42751 40477 42763 40511
rect 42705 40471 42763 40477
rect 40144 40412 40264 40440
rect 42536 40440 42564 40468
rect 42797 40443 42855 40449
rect 42797 40440 42809 40443
rect 42536 40412 42809 40440
rect 40144 40384 40172 40412
rect 42797 40409 42809 40412
rect 42843 40409 42855 40443
rect 42904 40440 42932 40616
rect 42981 40613 42993 40616
rect 43027 40613 43039 40647
rect 42981 40607 43039 40613
rect 43180 40576 43208 40672
rect 42996 40548 43208 40576
rect 42996 40517 43024 40548
rect 42981 40511 43039 40517
rect 42981 40477 42993 40511
rect 43027 40477 43039 40511
rect 42981 40471 43039 40477
rect 43165 40511 43223 40517
rect 43165 40477 43177 40511
rect 43211 40508 43223 40511
rect 43254 40508 43260 40520
rect 43211 40480 43260 40508
rect 43211 40477 43223 40480
rect 43165 40471 43223 40477
rect 43254 40468 43260 40480
rect 43312 40468 43318 40520
rect 43349 40511 43407 40517
rect 43349 40477 43361 40511
rect 43395 40508 43407 40511
rect 43441 40511 43499 40517
rect 43441 40508 43453 40511
rect 43395 40480 43453 40508
rect 43395 40477 43407 40480
rect 43349 40471 43407 40477
rect 43441 40477 43453 40480
rect 43487 40477 43499 40511
rect 43441 40471 43499 40477
rect 43993 40511 44051 40517
rect 43993 40477 44005 40511
rect 44039 40477 44051 40511
rect 43993 40471 44051 40477
rect 44008 40440 44036 40471
rect 42904 40412 44036 40440
rect 42797 40403 42855 40409
rect 35866 40344 36860 40372
rect 37001 40375 37059 40381
rect 37001 40341 37013 40375
rect 37047 40372 37059 40375
rect 37366 40372 37372 40384
rect 37047 40344 37372 40372
rect 37047 40341 37059 40344
rect 37001 40335 37059 40341
rect 37366 40332 37372 40344
rect 37424 40332 37430 40384
rect 40126 40332 40132 40384
rect 40184 40332 40190 40384
rect 40770 40332 40776 40384
rect 40828 40332 40834 40384
rect 1104 40282 44620 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 44620 40282
rect 1104 40208 44620 40230
rect 8570 40128 8576 40180
rect 8628 40128 8634 40180
rect 8754 40128 8760 40180
rect 8812 40168 8818 40180
rect 9033 40171 9091 40177
rect 9033 40168 9045 40171
rect 8812 40140 9045 40168
rect 8812 40128 8818 40140
rect 9033 40137 9045 40140
rect 9079 40137 9091 40171
rect 9033 40131 9091 40137
rect 9398 40128 9404 40180
rect 9456 40168 9462 40180
rect 10229 40171 10287 40177
rect 10229 40168 10241 40171
rect 9456 40140 10241 40168
rect 9456 40128 9462 40140
rect 10229 40137 10241 40140
rect 10275 40137 10287 40171
rect 10229 40131 10287 40137
rect 11333 40171 11391 40177
rect 11333 40137 11345 40171
rect 11379 40168 11391 40171
rect 12250 40168 12256 40180
rect 11379 40140 12256 40168
rect 11379 40137 11391 40140
rect 11333 40131 11391 40137
rect 8588 40100 8616 40128
rect 11348 40100 11376 40131
rect 12250 40128 12256 40140
rect 12308 40128 12314 40180
rect 13722 40128 13728 40180
rect 13780 40168 13786 40180
rect 19150 40168 19156 40180
rect 13780 40140 19156 40168
rect 13780 40128 13786 40140
rect 13924 40109 13952 40140
rect 19150 40128 19156 40140
rect 19208 40168 19214 40180
rect 19208 40140 21036 40168
rect 19208 40128 19214 40140
rect 21008 40112 21036 40140
rect 21082 40128 21088 40180
rect 21140 40128 21146 40180
rect 21821 40171 21879 40177
rect 21821 40137 21833 40171
rect 21867 40137 21879 40171
rect 21821 40131 21879 40137
rect 8588 40072 9904 40100
rect 9214 40032 9220 40044
rect 8234 40004 9220 40032
rect 9214 39992 9220 40004
rect 9272 39992 9278 40044
rect 9674 39992 9680 40044
rect 9732 39992 9738 40044
rect 9769 40035 9827 40041
rect 9769 40001 9781 40035
rect 9815 40001 9827 40035
rect 9769 39995 9827 40001
rect 6825 39967 6883 39973
rect 6825 39933 6837 39967
rect 6871 39933 6883 39967
rect 6825 39927 6883 39933
rect 6840 39828 6868 39927
rect 7098 39924 7104 39976
rect 7156 39924 7162 39976
rect 9122 39924 9128 39976
rect 9180 39924 9186 39976
rect 9309 39967 9367 39973
rect 9309 39933 9321 39967
rect 9355 39964 9367 39967
rect 9490 39964 9496 39976
rect 9355 39936 9496 39964
rect 9355 39933 9367 39936
rect 9309 39927 9367 39933
rect 9490 39924 9496 39936
rect 9548 39924 9554 39976
rect 9784 39964 9812 39995
rect 9692 39936 9812 39964
rect 9876 39964 9904 40072
rect 9968 40072 11376 40100
rect 13909 40103 13967 40109
rect 9968 40041 9996 40072
rect 13909 40069 13921 40103
rect 13955 40069 13967 40103
rect 13909 40063 13967 40069
rect 16117 40103 16175 40109
rect 16117 40069 16129 40103
rect 16163 40100 16175 40103
rect 16850 40100 16856 40112
rect 16163 40072 16856 40100
rect 16163 40069 16175 40072
rect 16117 40063 16175 40069
rect 16850 40060 16856 40072
rect 16908 40060 16914 40112
rect 16945 40103 17003 40109
rect 16945 40069 16957 40103
rect 16991 40100 17003 40103
rect 17218 40100 17224 40112
rect 16991 40072 17224 40100
rect 16991 40069 17003 40072
rect 16945 40063 17003 40069
rect 17218 40060 17224 40072
rect 17276 40060 17282 40112
rect 17402 40060 17408 40112
rect 17460 40060 17466 40112
rect 18785 40103 18843 40109
rect 18785 40069 18797 40103
rect 18831 40100 18843 40103
rect 19058 40100 19064 40112
rect 18831 40072 19064 40100
rect 18831 40069 18843 40072
rect 18785 40063 18843 40069
rect 19058 40060 19064 40072
rect 19116 40060 19122 40112
rect 20162 40100 20168 40112
rect 20010 40072 20168 40100
rect 20162 40060 20168 40072
rect 20220 40060 20226 40112
rect 20438 40100 20444 40112
rect 20272 40072 20444 40100
rect 9953 40035 10011 40041
rect 9953 40001 9965 40035
rect 9999 40001 10011 40035
rect 10965 40035 11023 40041
rect 10965 40032 10977 40035
rect 9953 39995 10011 40001
rect 10060 40004 10977 40032
rect 10060 39964 10088 40004
rect 10965 40001 10977 40004
rect 11011 40001 11023 40035
rect 11149 40035 11207 40041
rect 11149 40032 11161 40035
rect 10965 39995 11023 40001
rect 11072 40004 11161 40032
rect 9876 39936 10088 39964
rect 10137 39967 10195 39973
rect 8478 39828 8484 39840
rect 6840 39800 8484 39828
rect 8478 39788 8484 39800
rect 8536 39788 8542 39840
rect 8662 39788 8668 39840
rect 8720 39788 8726 39840
rect 9692 39828 9720 39936
rect 10137 39933 10149 39967
rect 10183 39964 10195 39967
rect 10781 39967 10839 39973
rect 10781 39964 10793 39967
rect 10183 39936 10793 39964
rect 10183 39933 10195 39936
rect 10137 39927 10195 39933
rect 10781 39933 10793 39936
rect 10827 39933 10839 39967
rect 10781 39927 10839 39933
rect 11072 39908 11100 40004
rect 11149 40001 11161 40004
rect 11195 40001 11207 40035
rect 11149 39995 11207 40001
rect 15470 39992 15476 40044
rect 15528 40032 15534 40044
rect 15528 40004 16344 40032
rect 15528 39992 15534 40004
rect 16132 39976 16160 40004
rect 12066 39924 12072 39976
rect 12124 39964 12130 39976
rect 12529 39967 12587 39973
rect 12529 39964 12541 39967
rect 12124 39936 12541 39964
rect 12124 39924 12130 39936
rect 12529 39933 12541 39936
rect 12575 39933 12587 39967
rect 12529 39927 12587 39933
rect 12802 39924 12808 39976
rect 12860 39924 12866 39976
rect 16114 39924 16120 39976
rect 16172 39924 16178 39976
rect 16206 39924 16212 39976
rect 16264 39924 16270 39976
rect 16316 39973 16344 40004
rect 18506 39992 18512 40044
rect 18564 39992 18570 40044
rect 16301 39967 16359 39973
rect 16301 39933 16313 39967
rect 16347 39933 16359 39967
rect 16301 39927 16359 39933
rect 16669 39967 16727 39973
rect 16669 39933 16681 39967
rect 16715 39933 16727 39967
rect 18782 39964 18788 39976
rect 16669 39927 16727 39933
rect 18524 39936 18788 39964
rect 10962 39856 10968 39908
rect 11020 39856 11026 39908
rect 11054 39856 11060 39908
rect 11112 39856 11118 39908
rect 16684 39896 16712 39927
rect 15212 39868 16712 39896
rect 10980 39828 11008 39856
rect 9692 39800 11008 39828
rect 11882 39788 11888 39840
rect 11940 39828 11946 39840
rect 11977 39831 12035 39837
rect 11977 39828 11989 39831
rect 11940 39800 11989 39828
rect 11940 39788 11946 39800
rect 11977 39797 11989 39800
rect 12023 39797 12035 39831
rect 11977 39791 12035 39797
rect 13354 39788 13360 39840
rect 13412 39788 13418 39840
rect 13998 39788 14004 39840
rect 14056 39828 14062 39840
rect 15102 39828 15108 39840
rect 14056 39800 15108 39828
rect 14056 39788 14062 39800
rect 15102 39788 15108 39800
rect 15160 39828 15166 39840
rect 15212 39837 15240 39868
rect 18414 39856 18420 39908
rect 18472 39896 18478 39908
rect 18524 39896 18552 39936
rect 18782 39924 18788 39936
rect 18840 39924 18846 39976
rect 20272 39973 20300 40072
rect 20438 40060 20444 40072
rect 20496 40060 20502 40112
rect 20990 40060 20996 40112
rect 21048 40060 21054 40112
rect 21836 40100 21864 40131
rect 22186 40128 22192 40180
rect 22244 40168 22250 40180
rect 22281 40171 22339 40177
rect 22281 40168 22293 40171
rect 22244 40140 22293 40168
rect 22244 40128 22250 40140
rect 22281 40137 22293 40140
rect 22327 40137 22339 40171
rect 24026 40168 24032 40180
rect 22281 40131 22339 40137
rect 23768 40140 24032 40168
rect 23768 40109 23796 40140
rect 24026 40128 24032 40140
rect 24084 40128 24090 40180
rect 24118 40128 24124 40180
rect 24176 40128 24182 40180
rect 35986 40128 35992 40180
rect 36044 40128 36050 40180
rect 23753 40103 23811 40109
rect 21284 40072 21864 40100
rect 22066 40072 23520 40100
rect 21284 40041 21312 40072
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40001 21327 40035
rect 21269 39995 21327 40001
rect 22066 39976 22094 40072
rect 22186 39992 22192 40044
rect 22244 39992 22250 40044
rect 23492 40041 23520 40072
rect 23753 40069 23765 40103
rect 23799 40069 23811 40103
rect 23753 40063 23811 40069
rect 23845 40103 23903 40109
rect 23845 40069 23857 40103
rect 23891 40100 23903 40103
rect 36078 40100 36084 40112
rect 23891 40072 25912 40100
rect 35742 40072 36084 40100
rect 23891 40069 23903 40072
rect 23845 40063 23903 40069
rect 25884 40044 25912 40072
rect 36078 40060 36084 40072
rect 36136 40060 36142 40112
rect 41138 40100 41144 40112
rect 39974 40072 41144 40100
rect 41138 40060 41144 40072
rect 41196 40060 41202 40112
rect 43272 40072 43668 40100
rect 43272 40044 43300 40072
rect 23477 40035 23535 40041
rect 23477 40001 23489 40035
rect 23523 40001 23535 40035
rect 23477 39995 23535 40001
rect 23566 39992 23572 40044
rect 23624 40041 23630 40044
rect 23624 40035 23655 40041
rect 23643 40001 23655 40035
rect 23624 39995 23655 40001
rect 23942 40035 24000 40041
rect 23942 40001 23954 40035
rect 23988 40032 24000 40035
rect 23988 40004 24072 40032
rect 23988 40001 24000 40004
rect 23942 39995 24000 40001
rect 23624 39992 23630 39995
rect 20257 39967 20315 39973
rect 20257 39933 20269 39967
rect 20303 39933 20315 39967
rect 20257 39927 20315 39933
rect 20714 39924 20720 39976
rect 20772 39964 20778 39976
rect 22002 39964 22008 39976
rect 20772 39936 22008 39964
rect 20772 39924 20778 39936
rect 22002 39924 22008 39936
rect 22060 39936 22094 39976
rect 22465 39967 22523 39973
rect 22060 39924 22066 39936
rect 22465 39933 22477 39967
rect 22511 39933 22523 39967
rect 22465 39927 22523 39933
rect 18472 39868 18552 39896
rect 18472 39856 18478 39868
rect 15197 39831 15255 39837
rect 15197 39828 15209 39831
rect 15160 39800 15209 39828
rect 15160 39788 15166 39800
rect 15197 39797 15209 39800
rect 15243 39797 15255 39831
rect 15197 39791 15255 39797
rect 15746 39788 15752 39840
rect 15804 39788 15810 39840
rect 20254 39788 20260 39840
rect 20312 39828 20318 39840
rect 22370 39828 22376 39840
rect 20312 39800 22376 39828
rect 20312 39788 20318 39800
rect 22370 39788 22376 39800
rect 22428 39828 22434 39840
rect 22480 39828 22508 39927
rect 24044 39896 24072 40004
rect 25866 39992 25872 40044
rect 25924 39992 25930 40044
rect 26970 39992 26976 40044
rect 27028 40032 27034 40044
rect 27157 40035 27215 40041
rect 27157 40032 27169 40035
rect 27028 40004 27169 40032
rect 27028 39992 27034 40004
rect 27157 40001 27169 40004
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 40586 39992 40592 40044
rect 40644 39992 40650 40044
rect 40770 39992 40776 40044
rect 40828 40032 40834 40044
rect 41233 40035 41291 40041
rect 41233 40032 41245 40035
rect 40828 40004 41245 40032
rect 40828 39992 40834 40004
rect 41233 40001 41245 40004
rect 41279 40001 41291 40035
rect 41233 39995 41291 40001
rect 41417 40035 41475 40041
rect 41417 40001 41429 40035
rect 41463 40032 41475 40035
rect 41874 40032 41880 40044
rect 41463 40004 41880 40032
rect 41463 40001 41475 40004
rect 41417 39995 41475 40001
rect 41874 39992 41880 40004
rect 41932 39992 41938 40044
rect 43254 39992 43260 40044
rect 43312 39992 43318 40044
rect 43640 40041 43668 40072
rect 43349 40035 43407 40041
rect 43349 40001 43361 40035
rect 43395 40032 43407 40035
rect 43441 40035 43499 40041
rect 43441 40032 43453 40035
rect 43395 40004 43453 40032
rect 43395 40001 43407 40004
rect 43349 39995 43407 40001
rect 43441 40001 43453 40004
rect 43487 40001 43499 40035
rect 43441 39995 43499 40001
rect 43625 40035 43683 40041
rect 43625 40001 43637 40035
rect 43671 40001 43683 40035
rect 43625 39995 43683 40001
rect 24578 39924 24584 39976
rect 24636 39924 24642 39976
rect 32306 39924 32312 39976
rect 32364 39964 32370 39976
rect 32401 39967 32459 39973
rect 32401 39964 32413 39967
rect 32364 39936 32413 39964
rect 32364 39924 32370 39936
rect 32401 39933 32413 39936
rect 32447 39933 32459 39967
rect 32401 39927 32459 39933
rect 34241 39967 34299 39973
rect 34241 39933 34253 39967
rect 34287 39933 34299 39967
rect 34241 39927 34299 39933
rect 24210 39896 24216 39908
rect 24044 39868 24216 39896
rect 24210 39856 24216 39868
rect 24268 39896 24274 39908
rect 24268 39868 26740 39896
rect 24268 39856 24274 39868
rect 26712 39840 26740 39868
rect 22428 39800 22508 39828
rect 22428 39788 22434 39800
rect 25222 39788 25228 39840
rect 25280 39788 25286 39840
rect 25314 39788 25320 39840
rect 25372 39788 25378 39840
rect 26694 39788 26700 39840
rect 26752 39788 26758 39840
rect 26786 39788 26792 39840
rect 26844 39828 26850 39840
rect 26973 39831 27031 39837
rect 26973 39828 26985 39831
rect 26844 39800 26985 39828
rect 26844 39788 26850 39800
rect 26973 39797 26985 39800
rect 27019 39797 27031 39831
rect 26973 39791 27031 39797
rect 32766 39788 32772 39840
rect 32824 39828 32830 39840
rect 33045 39831 33103 39837
rect 33045 39828 33057 39831
rect 32824 39800 33057 39828
rect 32824 39788 32830 39800
rect 33045 39797 33057 39800
rect 33091 39797 33103 39831
rect 34256 39828 34284 39927
rect 34514 39924 34520 39976
rect 34572 39924 34578 39976
rect 38470 39924 38476 39976
rect 38528 39924 38534 39976
rect 38746 39924 38752 39976
rect 38804 39924 38810 39976
rect 40221 39967 40279 39973
rect 40221 39933 40233 39967
rect 40267 39964 40279 39967
rect 40604 39964 40632 39992
rect 40267 39936 40632 39964
rect 42705 39967 42763 39973
rect 40267 39933 40279 39936
rect 40221 39927 40279 39933
rect 42705 39933 42717 39967
rect 42751 39964 42763 39967
rect 42794 39964 42800 39976
rect 42751 39936 42800 39964
rect 42751 39933 42763 39936
rect 42705 39927 42763 39933
rect 42794 39924 42800 39936
rect 42852 39924 42858 39976
rect 34698 39828 34704 39840
rect 34256 39800 34704 39828
rect 33045 39791 33103 39797
rect 34698 39788 34704 39800
rect 34756 39788 34762 39840
rect 41138 39788 41144 39840
rect 41196 39788 41202 39840
rect 41230 39788 41236 39840
rect 41288 39788 41294 39840
rect 42886 39788 42892 39840
rect 42944 39828 42950 39840
rect 43625 39831 43683 39837
rect 43625 39828 43637 39831
rect 42944 39800 43637 39828
rect 42944 39788 42950 39800
rect 43625 39797 43637 39800
rect 43671 39797 43683 39831
rect 43625 39791 43683 39797
rect 1104 39738 44620 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 44620 39738
rect 1104 39664 44620 39686
rect 7098 39584 7104 39636
rect 7156 39624 7162 39636
rect 7377 39627 7435 39633
rect 7377 39624 7389 39627
rect 7156 39596 7389 39624
rect 7156 39584 7162 39596
rect 7377 39593 7389 39596
rect 7423 39593 7435 39627
rect 7377 39587 7435 39593
rect 13265 39627 13323 39633
rect 13265 39593 13277 39627
rect 13311 39624 13323 39627
rect 13538 39624 13544 39636
rect 13311 39596 13544 39624
rect 13311 39593 13323 39596
rect 13265 39587 13323 39593
rect 13538 39584 13544 39596
rect 13596 39584 13602 39636
rect 15746 39624 15752 39636
rect 13740 39596 15752 39624
rect 8478 39448 8484 39500
rect 8536 39488 8542 39500
rect 9398 39488 9404 39500
rect 8536 39460 9404 39488
rect 8536 39448 8542 39460
rect 9398 39448 9404 39460
rect 9456 39488 9462 39500
rect 9585 39491 9643 39497
rect 9585 39488 9597 39491
rect 9456 39460 9597 39488
rect 9456 39448 9462 39460
rect 9585 39457 9597 39460
rect 9631 39488 9643 39491
rect 11517 39491 11575 39497
rect 11517 39488 11529 39491
rect 9631 39460 11529 39488
rect 9631 39457 9643 39460
rect 9585 39451 9643 39457
rect 11517 39457 11529 39460
rect 11563 39457 11575 39491
rect 11517 39451 11575 39457
rect 11793 39491 11851 39497
rect 11793 39457 11805 39491
rect 11839 39488 11851 39491
rect 11882 39488 11888 39500
rect 11839 39460 11888 39488
rect 11839 39457 11851 39460
rect 11793 39451 11851 39457
rect 11882 39448 11888 39460
rect 11940 39448 11946 39500
rect 7561 39423 7619 39429
rect 7561 39389 7573 39423
rect 7607 39420 7619 39423
rect 8662 39420 8668 39432
rect 7607 39392 8668 39420
rect 7607 39389 7619 39392
rect 7561 39383 7619 39389
rect 8662 39380 8668 39392
rect 8720 39380 8726 39432
rect 13740 39429 13768 39596
rect 15746 39584 15752 39596
rect 15804 39584 15810 39636
rect 17037 39627 17095 39633
rect 17037 39593 17049 39627
rect 17083 39624 17095 39627
rect 17954 39624 17960 39636
rect 17083 39596 17960 39624
rect 17083 39593 17095 39596
rect 17037 39587 17095 39593
rect 17954 39584 17960 39596
rect 18012 39584 18018 39636
rect 20714 39624 20720 39636
rect 19352 39596 20720 39624
rect 16025 39559 16083 39565
rect 16025 39525 16037 39559
rect 16071 39556 16083 39559
rect 17497 39559 17555 39565
rect 16071 39528 17172 39556
rect 16071 39525 16083 39528
rect 16025 39519 16083 39525
rect 16114 39448 16120 39500
rect 16172 39488 16178 39500
rect 17144 39497 17172 39528
rect 17497 39525 17509 39559
rect 17543 39556 17555 39559
rect 19352 39556 19380 39596
rect 20714 39584 20720 39596
rect 20772 39584 20778 39636
rect 25866 39584 25872 39636
rect 25924 39624 25930 39636
rect 26145 39627 26203 39633
rect 26145 39624 26157 39627
rect 25924 39596 26157 39624
rect 25924 39584 25930 39596
rect 26145 39593 26157 39596
rect 26191 39593 26203 39627
rect 26145 39587 26203 39593
rect 34514 39584 34520 39636
rect 34572 39624 34578 39636
rect 35069 39627 35127 39633
rect 35069 39624 35081 39627
rect 34572 39596 35081 39624
rect 34572 39584 34578 39596
rect 35069 39593 35081 39596
rect 35115 39593 35127 39627
rect 35069 39587 35127 39593
rect 38746 39584 38752 39636
rect 38804 39624 38810 39636
rect 39393 39627 39451 39633
rect 39393 39624 39405 39627
rect 38804 39596 39405 39624
rect 38804 39584 38810 39596
rect 39393 39593 39405 39596
rect 39439 39593 39451 39627
rect 39393 39587 39451 39593
rect 39942 39584 39948 39636
rect 40000 39624 40006 39636
rect 40037 39627 40095 39633
rect 40037 39624 40049 39627
rect 40000 39596 40049 39624
rect 40000 39584 40006 39596
rect 40037 39593 40049 39596
rect 40083 39593 40095 39627
rect 40037 39587 40095 39593
rect 40126 39584 40132 39636
rect 40184 39624 40190 39636
rect 40221 39627 40279 39633
rect 40221 39624 40233 39627
rect 40184 39596 40233 39624
rect 40184 39584 40190 39596
rect 40221 39593 40233 39596
rect 40267 39593 40279 39627
rect 40221 39587 40279 39593
rect 42429 39627 42487 39633
rect 42429 39593 42441 39627
rect 42475 39624 42487 39627
rect 42794 39624 42800 39636
rect 42475 39596 42800 39624
rect 42475 39593 42487 39596
rect 42429 39587 42487 39593
rect 42794 39584 42800 39596
rect 42852 39584 42858 39636
rect 42886 39584 42892 39636
rect 42944 39584 42950 39636
rect 39960 39556 39988 39584
rect 42904 39556 42932 39584
rect 17543 39528 19380 39556
rect 39224 39528 39988 39556
rect 42352 39528 42932 39556
rect 17543 39525 17555 39528
rect 17497 39519 17555 39525
rect 16393 39491 16451 39497
rect 16393 39488 16405 39491
rect 16172 39460 16405 39488
rect 16172 39448 16178 39460
rect 16393 39457 16405 39460
rect 16439 39457 16451 39491
rect 16393 39451 16451 39457
rect 17129 39491 17187 39497
rect 17129 39457 17141 39491
rect 17175 39488 17187 39491
rect 17678 39488 17684 39500
rect 17175 39460 17684 39488
rect 17175 39457 17187 39460
rect 17129 39451 17187 39457
rect 17678 39448 17684 39460
rect 17736 39448 17742 39500
rect 18233 39491 18291 39497
rect 18233 39457 18245 39491
rect 18279 39488 18291 39491
rect 18414 39488 18420 39500
rect 18279 39460 18420 39488
rect 18279 39457 18291 39460
rect 18233 39451 18291 39457
rect 18414 39448 18420 39460
rect 18472 39448 18478 39500
rect 18506 39448 18512 39500
rect 18564 39488 18570 39500
rect 19245 39491 19303 39497
rect 19245 39488 19257 39491
rect 18564 39460 19257 39488
rect 18564 39448 18570 39460
rect 19245 39457 19257 39460
rect 19291 39457 19303 39491
rect 19245 39451 19303 39457
rect 24394 39448 24400 39500
rect 24452 39488 24458 39500
rect 26142 39488 26148 39500
rect 24452 39460 26148 39488
rect 24452 39448 24458 39460
rect 26142 39448 26148 39460
rect 26200 39488 26206 39500
rect 26421 39491 26479 39497
rect 26421 39488 26433 39491
rect 26200 39460 26433 39488
rect 26200 39448 26206 39460
rect 26421 39457 26433 39460
rect 26467 39457 26479 39491
rect 26421 39451 26479 39457
rect 26697 39491 26755 39497
rect 26697 39457 26709 39491
rect 26743 39488 26755 39491
rect 26786 39488 26792 39500
rect 26743 39460 26792 39488
rect 26743 39457 26755 39460
rect 26697 39451 26755 39457
rect 26786 39448 26792 39460
rect 26844 39448 26850 39500
rect 27430 39448 27436 39500
rect 27488 39488 27494 39500
rect 27488 39460 27844 39488
rect 27488 39448 27494 39460
rect 13725 39423 13783 39429
rect 13725 39389 13737 39423
rect 13771 39389 13783 39423
rect 13725 39383 13783 39389
rect 13998 39380 14004 39432
rect 14056 39420 14062 39432
rect 14277 39423 14335 39429
rect 14277 39420 14289 39423
rect 14056 39392 14289 39420
rect 14056 39380 14062 39392
rect 14277 39389 14289 39392
rect 14323 39389 14335 39423
rect 14277 39383 14335 39389
rect 17313 39423 17371 39429
rect 17313 39389 17325 39423
rect 17359 39420 17371 39423
rect 17359 39392 18184 39420
rect 17359 39389 17371 39392
rect 17313 39383 17371 39389
rect 9858 39312 9864 39364
rect 9916 39312 9922 39364
rect 10870 39312 10876 39364
rect 10928 39312 10934 39364
rect 14553 39355 14611 39361
rect 14553 39352 14565 39355
rect 11256 39324 12291 39352
rect 9582 39244 9588 39296
rect 9640 39284 9646 39296
rect 11256 39284 11284 39324
rect 9640 39256 11284 39284
rect 11333 39287 11391 39293
rect 9640 39244 9646 39256
rect 11333 39253 11345 39287
rect 11379 39284 11391 39287
rect 11514 39284 11520 39296
rect 11379 39256 11520 39284
rect 11379 39253 11391 39256
rect 11333 39247 11391 39253
rect 11514 39244 11520 39256
rect 11572 39244 11578 39296
rect 12263 39284 12291 39324
rect 13924 39324 14565 39352
rect 12618 39284 12624 39296
rect 12263 39256 12624 39284
rect 12618 39244 12624 39256
rect 12676 39244 12682 39296
rect 13924 39293 13952 39324
rect 14553 39321 14565 39324
rect 14599 39321 14611 39355
rect 16022 39352 16028 39364
rect 15778 39324 16028 39352
rect 14553 39315 14611 39321
rect 16022 39312 16028 39324
rect 16080 39312 16086 39364
rect 16669 39355 16727 39361
rect 16669 39321 16681 39355
rect 16715 39352 16727 39355
rect 17589 39355 17647 39361
rect 17589 39352 17601 39355
rect 16715 39324 17601 39352
rect 16715 39321 16727 39324
rect 16669 39315 16727 39321
rect 17589 39321 17601 39324
rect 17635 39321 17647 39355
rect 17589 39315 17647 39321
rect 18156 39296 18184 39392
rect 18874 39380 18880 39432
rect 18932 39380 18938 39432
rect 20622 39380 20628 39432
rect 20680 39380 20686 39432
rect 20806 39380 20812 39432
rect 20864 39420 20870 39432
rect 22281 39423 22339 39429
rect 22281 39420 22293 39423
rect 20864 39392 22293 39420
rect 20864 39380 20870 39392
rect 22281 39389 22293 39392
rect 22327 39389 22339 39423
rect 22281 39383 22339 39389
rect 19521 39355 19579 39361
rect 19521 39352 19533 39355
rect 19076 39324 19533 39352
rect 13909 39287 13967 39293
rect 13909 39253 13921 39287
rect 13955 39253 13967 39287
rect 13909 39247 13967 39253
rect 16574 39244 16580 39296
rect 16632 39244 16638 39296
rect 18138 39244 18144 39296
rect 18196 39244 18202 39296
rect 19076 39293 19104 39324
rect 19521 39321 19533 39324
rect 19567 39321 19579 39355
rect 22296 39352 22324 39383
rect 22554 39380 22560 39432
rect 22612 39420 22618 39432
rect 22922 39420 22928 39432
rect 22612 39392 22928 39420
rect 22612 39380 22618 39392
rect 22922 39380 22928 39392
rect 22980 39380 22986 39432
rect 24673 39355 24731 39361
rect 22296 39324 23796 39352
rect 19521 39315 19579 39321
rect 23768 39296 23796 39324
rect 24673 39321 24685 39355
rect 24719 39352 24731 39355
rect 24946 39352 24952 39364
rect 24719 39324 24952 39352
rect 24719 39321 24731 39324
rect 24673 39315 24731 39321
rect 24946 39312 24952 39324
rect 25004 39312 25010 39364
rect 25898 39324 26556 39352
rect 19061 39287 19119 39293
rect 19061 39253 19073 39287
rect 19107 39253 19119 39287
rect 19061 39247 19119 39253
rect 20346 39244 20352 39296
rect 20404 39284 20410 39296
rect 20993 39287 21051 39293
rect 20993 39284 21005 39287
rect 20404 39256 21005 39284
rect 20404 39244 20410 39256
rect 20993 39253 21005 39256
rect 21039 39284 21051 39287
rect 21266 39284 21272 39296
rect 21039 39256 21272 39284
rect 21039 39253 21051 39256
rect 20993 39247 21051 39253
rect 21266 39244 21272 39256
rect 21324 39244 21330 39296
rect 22094 39244 22100 39296
rect 22152 39244 22158 39296
rect 22278 39244 22284 39296
rect 22336 39284 22342 39296
rect 22465 39287 22523 39293
rect 22465 39284 22477 39287
rect 22336 39256 22477 39284
rect 22336 39244 22342 39256
rect 22465 39253 22477 39256
rect 22511 39253 22523 39287
rect 22465 39247 22523 39253
rect 23750 39244 23756 39296
rect 23808 39244 23814 39296
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 26326 39284 26332 39296
rect 24360 39256 26332 39284
rect 24360 39244 24366 39256
rect 26326 39244 26332 39256
rect 26384 39244 26390 39296
rect 26528 39284 26556 39324
rect 27816 39284 27844 39460
rect 27890 39448 27896 39500
rect 27948 39488 27954 39500
rect 28169 39491 28227 39497
rect 28169 39488 28181 39491
rect 27948 39460 28181 39488
rect 27948 39448 27954 39460
rect 28169 39457 28181 39460
rect 28215 39488 28227 39491
rect 28902 39488 28908 39500
rect 28215 39460 28908 39488
rect 28215 39457 28227 39460
rect 28169 39451 28227 39457
rect 28902 39448 28908 39460
rect 28960 39488 28966 39500
rect 31662 39488 31668 39500
rect 28960 39460 29040 39488
rect 28960 39448 28966 39460
rect 29012 39429 29040 39460
rect 30576 39460 31668 39488
rect 28997 39423 29055 39429
rect 28997 39389 29009 39423
rect 29043 39389 29055 39423
rect 28997 39383 29055 39389
rect 28813 39355 28871 39361
rect 28813 39321 28825 39355
rect 28859 39352 28871 39355
rect 29454 39352 29460 39364
rect 28859 39324 29460 39352
rect 28859 39321 28871 39324
rect 28813 39315 28871 39321
rect 29454 39312 29460 39324
rect 29512 39312 29518 39364
rect 30374 39352 30380 39364
rect 30208 39324 30380 39352
rect 26528 39256 27844 39284
rect 28534 39244 28540 39296
rect 28592 39284 28598 39296
rect 28629 39287 28687 39293
rect 28629 39284 28641 39287
rect 28592 39256 28641 39284
rect 28592 39244 28598 39256
rect 28629 39253 28641 39256
rect 28675 39253 28687 39287
rect 28629 39247 28687 39253
rect 28718 39244 28724 39296
rect 28776 39284 28782 39296
rect 30208 39284 30236 39324
rect 30374 39312 30380 39324
rect 30432 39352 30438 39364
rect 30576 39352 30604 39460
rect 31662 39448 31668 39460
rect 31720 39448 31726 39500
rect 31754 39448 31760 39500
rect 31812 39448 31818 39500
rect 32030 39448 32036 39500
rect 32088 39488 32094 39500
rect 32125 39491 32183 39497
rect 32125 39488 32137 39491
rect 32088 39460 32137 39488
rect 32088 39448 32094 39460
rect 32125 39457 32137 39460
rect 32171 39457 32183 39491
rect 32125 39451 32183 39457
rect 32401 39491 32459 39497
rect 32401 39457 32413 39491
rect 32447 39488 32459 39491
rect 32490 39488 32496 39500
rect 32447 39460 32496 39488
rect 32447 39457 32459 39460
rect 32401 39451 32459 39457
rect 32490 39448 32496 39460
rect 32548 39448 32554 39500
rect 34606 39380 34612 39432
rect 34664 39420 34670 39432
rect 35069 39423 35127 39429
rect 35069 39420 35081 39423
rect 34664 39392 35081 39420
rect 34664 39380 34670 39392
rect 35069 39389 35081 39392
rect 35115 39389 35127 39423
rect 35069 39383 35127 39389
rect 35253 39423 35311 39429
rect 35253 39389 35265 39423
rect 35299 39420 35311 39423
rect 35526 39420 35532 39432
rect 35299 39392 35532 39420
rect 35299 39389 35311 39392
rect 35253 39383 35311 39389
rect 35526 39380 35532 39392
rect 35584 39380 35590 39432
rect 38013 39423 38071 39429
rect 38013 39389 38025 39423
rect 38059 39389 38071 39423
rect 38013 39383 38071 39389
rect 38197 39423 38255 39429
rect 38197 39389 38209 39423
rect 38243 39420 38255 39423
rect 38746 39420 38752 39432
rect 38243 39392 38752 39420
rect 38243 39389 38255 39392
rect 38197 39383 38255 39389
rect 30432 39338 30604 39352
rect 30432 39324 30590 39338
rect 30432 39312 30438 39324
rect 31662 39312 31668 39364
rect 31720 39352 31726 39364
rect 38028 39352 38056 39383
rect 38746 39380 38752 39392
rect 38804 39380 38810 39432
rect 39224 39429 39252 39528
rect 40589 39491 40647 39497
rect 40589 39488 40601 39491
rect 39408 39460 40601 39488
rect 39408 39429 39436 39460
rect 40589 39457 40601 39460
rect 40635 39457 40647 39491
rect 40589 39451 40647 39457
rect 39209 39423 39267 39429
rect 39209 39389 39221 39423
rect 39255 39389 39267 39423
rect 39209 39383 39267 39389
rect 39393 39423 39451 39429
rect 39393 39389 39405 39423
rect 39439 39389 39451 39423
rect 39393 39383 39451 39389
rect 40218 39380 40224 39432
rect 40276 39420 40282 39432
rect 40497 39423 40555 39429
rect 40497 39420 40509 39423
rect 40276 39392 40509 39420
rect 40276 39380 40282 39392
rect 40497 39389 40509 39392
rect 40543 39389 40555 39423
rect 40497 39383 40555 39389
rect 40681 39423 40739 39429
rect 40681 39389 40693 39423
rect 40727 39420 40739 39423
rect 41138 39420 41144 39432
rect 40727 39392 41144 39420
rect 40727 39389 40739 39392
rect 40681 39383 40739 39389
rect 41138 39380 41144 39392
rect 41196 39380 41202 39432
rect 42150 39380 42156 39432
rect 42208 39380 42214 39432
rect 42352 39429 42380 39528
rect 42426 39448 42432 39500
rect 42484 39488 42490 39500
rect 44174 39488 44180 39500
rect 42484 39460 44180 39488
rect 42484 39448 42490 39460
rect 44174 39448 44180 39460
rect 44232 39448 44238 39500
rect 42337 39423 42395 39429
rect 42337 39389 42349 39423
rect 42383 39389 42395 39423
rect 42337 39383 42395 39389
rect 42518 39380 42524 39432
rect 42576 39420 42582 39432
rect 42576 39392 42826 39420
rect 42576 39380 42582 39392
rect 40405 39355 40463 39361
rect 31720 39324 32352 39352
rect 31720 39312 31726 39324
rect 28776 39256 30236 39284
rect 30285 39287 30343 39293
rect 28776 39244 28782 39256
rect 30285 39253 30297 39287
rect 30331 39284 30343 39287
rect 32214 39284 32220 39296
rect 30331 39256 32220 39284
rect 30331 39253 30343 39256
rect 30285 39247 30343 39253
rect 32214 39244 32220 39256
rect 32272 39244 32278 39296
rect 32324 39284 32352 39324
rect 32508 39324 32890 39352
rect 38028 39324 40172 39352
rect 32508 39284 32536 39324
rect 38212 39296 38240 39324
rect 32324 39256 32536 39284
rect 33870 39244 33876 39296
rect 33928 39244 33934 39296
rect 38102 39244 38108 39296
rect 38160 39244 38166 39296
rect 38194 39244 38200 39296
rect 38252 39244 38258 39296
rect 40144 39284 40172 39324
rect 40405 39321 40417 39355
rect 40451 39352 40463 39355
rect 40586 39352 40592 39364
rect 40451 39324 40592 39352
rect 40451 39321 40463 39324
rect 40405 39315 40463 39321
rect 40586 39312 40592 39324
rect 40644 39312 40650 39364
rect 42245 39355 42303 39361
rect 42245 39321 42257 39355
rect 42291 39352 42303 39355
rect 43901 39355 43959 39361
rect 42291 39324 42656 39352
rect 42291 39321 42303 39324
rect 42245 39315 42303 39321
rect 40200 39287 40258 39293
rect 40200 39284 40212 39287
rect 40144 39256 40212 39284
rect 40200 39253 40212 39256
rect 40246 39284 40258 39287
rect 40310 39284 40316 39296
rect 40246 39256 40316 39284
rect 40246 39253 40258 39256
rect 40200 39247 40258 39253
rect 40310 39244 40316 39256
rect 40368 39244 40374 39296
rect 42628 39284 42656 39324
rect 43901 39321 43913 39355
rect 43947 39321 43959 39355
rect 43901 39315 43959 39321
rect 43916 39284 43944 39315
rect 42628 39256 43944 39284
rect 1104 39194 44620 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 44620 39194
rect 1104 39120 44620 39142
rect 7653 39083 7711 39089
rect 7653 39049 7665 39083
rect 7699 39049 7711 39083
rect 7653 39043 7711 39049
rect 7285 38947 7343 38953
rect 7285 38913 7297 38947
rect 7331 38944 7343 38947
rect 7668 38944 7696 39043
rect 9582 39040 9588 39092
rect 9640 39040 9646 39092
rect 9858 39040 9864 39092
rect 9916 39080 9922 39092
rect 10045 39083 10103 39089
rect 10045 39080 10057 39083
rect 9916 39052 10057 39080
rect 9916 39040 9922 39052
rect 10045 39049 10057 39052
rect 10091 39049 10103 39083
rect 10045 39043 10103 39049
rect 10505 39083 10563 39089
rect 10505 39049 10517 39083
rect 10551 39049 10563 39083
rect 10505 39043 10563 39049
rect 7331 38916 7696 38944
rect 8021 38947 8079 38953
rect 7331 38913 7343 38916
rect 7285 38907 7343 38913
rect 8021 38913 8033 38947
rect 8067 38944 8079 38947
rect 8481 38947 8539 38953
rect 8481 38944 8493 38947
rect 8067 38916 8493 38944
rect 8067 38913 8079 38916
rect 8021 38907 8079 38913
rect 8481 38913 8493 38916
rect 8527 38913 8539 38947
rect 8481 38907 8539 38913
rect 9214 38904 9220 38956
rect 9272 38944 9278 38956
rect 9309 38947 9367 38953
rect 9309 38944 9321 38947
rect 9272 38916 9321 38944
rect 9272 38904 9278 38916
rect 9309 38913 9321 38916
rect 9355 38944 9367 38947
rect 10229 38947 10287 38953
rect 9355 38916 10180 38944
rect 9355 38913 9367 38916
rect 9309 38907 9367 38913
rect 7834 38836 7840 38888
rect 7892 38876 7898 38888
rect 8113 38879 8171 38885
rect 8113 38876 8125 38879
rect 7892 38848 8125 38876
rect 7892 38836 7898 38848
rect 8113 38845 8125 38848
rect 8159 38845 8171 38879
rect 8113 38839 8171 38845
rect 8297 38879 8355 38885
rect 8297 38845 8309 38879
rect 8343 38845 8355 38879
rect 8297 38839 8355 38845
rect 8202 38768 8208 38820
rect 8260 38808 8266 38820
rect 8312 38808 8340 38839
rect 9030 38836 9036 38888
rect 9088 38836 9094 38888
rect 9490 38836 9496 38888
rect 9548 38836 9554 38888
rect 10152 38876 10180 38916
rect 10229 38913 10241 38947
rect 10275 38944 10287 38947
rect 10520 38944 10548 39043
rect 10962 39040 10968 39092
rect 11020 39040 11026 39092
rect 12066 39040 12072 39092
rect 12124 39040 12130 39092
rect 12802 39040 12808 39092
rect 12860 39040 12866 39092
rect 13354 39080 13360 39092
rect 12912 39052 13360 39080
rect 12437 39015 12495 39021
rect 12437 38981 12449 39015
rect 12483 39012 12495 39015
rect 12526 39012 12532 39024
rect 12483 38984 12532 39012
rect 12483 38981 12495 38984
rect 12437 38975 12495 38981
rect 12526 38972 12532 38984
rect 12584 38972 12590 39024
rect 12912 39012 12940 39052
rect 13354 39040 13360 39052
rect 13412 39040 13418 39092
rect 15286 39080 15292 39092
rect 13924 39052 15292 39080
rect 13924 39012 13952 39052
rect 15286 39040 15292 39052
rect 15344 39080 15350 39092
rect 15473 39083 15531 39089
rect 15473 39080 15485 39083
rect 15344 39052 15485 39080
rect 15344 39040 15350 39052
rect 15473 39049 15485 39052
rect 15519 39049 15531 39083
rect 15473 39043 15531 39049
rect 18874 39040 18880 39092
rect 18932 39080 18938 39092
rect 19521 39083 19579 39089
rect 19521 39080 19533 39083
rect 18932 39052 19533 39080
rect 18932 39040 18938 39052
rect 19521 39049 19533 39052
rect 19567 39049 19579 39083
rect 19521 39043 19579 39049
rect 19981 39083 20039 39089
rect 19981 39049 19993 39083
rect 20027 39080 20039 39083
rect 20070 39080 20076 39092
rect 20027 39052 20076 39080
rect 20027 39049 20039 39052
rect 19981 39043 20039 39049
rect 20070 39040 20076 39052
rect 20128 39040 20134 39092
rect 20806 39040 20812 39092
rect 20864 39040 20870 39092
rect 24302 39040 24308 39092
rect 24360 39040 24366 39092
rect 24397 39083 24455 39089
rect 24397 39049 24409 39083
rect 24443 39080 24455 39083
rect 24578 39080 24584 39092
rect 24443 39052 24584 39080
rect 24443 39049 24455 39052
rect 24397 39043 24455 39049
rect 24578 39040 24584 39052
rect 24636 39040 24642 39092
rect 31754 39040 31760 39092
rect 31812 39080 31818 39092
rect 32125 39083 32183 39089
rect 32125 39080 32137 39083
rect 31812 39052 32137 39080
rect 31812 39040 31818 39052
rect 32125 39049 32137 39052
rect 32171 39049 32183 39083
rect 32950 39080 32956 39092
rect 32125 39043 32183 39049
rect 32784 39052 32956 39080
rect 12636 38984 12940 39012
rect 13846 38984 13952 39012
rect 10275 38916 10548 38944
rect 10873 38947 10931 38953
rect 10275 38913 10287 38916
rect 10229 38907 10287 38913
rect 10873 38913 10885 38947
rect 10919 38944 10931 38947
rect 11514 38944 11520 38956
rect 10919 38916 11520 38944
rect 10919 38913 10931 38916
rect 10873 38907 10931 38913
rect 11514 38904 11520 38916
rect 11572 38904 11578 38956
rect 12636 38953 12664 38984
rect 13998 38972 14004 39024
rect 14056 39012 14062 39024
rect 18141 39015 18199 39021
rect 14056 38984 14596 39012
rect 14056 38972 14062 38984
rect 12248 38947 12306 38953
rect 12248 38913 12260 38947
rect 12294 38913 12306 38947
rect 12248 38907 12306 38913
rect 12345 38947 12403 38953
rect 12345 38913 12357 38947
rect 12391 38913 12403 38947
rect 12345 38907 12403 38913
rect 12620 38947 12678 38953
rect 12620 38913 12632 38947
rect 12666 38913 12678 38947
rect 12620 38907 12678 38913
rect 10962 38876 10968 38888
rect 10152 38848 10968 38876
rect 10962 38836 10968 38848
rect 11020 38836 11026 38888
rect 11149 38879 11207 38885
rect 11149 38845 11161 38879
rect 11195 38876 11207 38879
rect 11330 38876 11336 38888
rect 11195 38848 11336 38876
rect 11195 38845 11207 38848
rect 11149 38839 11207 38845
rect 11330 38836 11336 38848
rect 11388 38876 11394 38888
rect 11974 38876 11980 38888
rect 11388 38848 11980 38876
rect 11388 38836 11394 38848
rect 11974 38836 11980 38848
rect 12032 38836 12038 38888
rect 9508 38808 9536 38836
rect 8260 38780 9536 38808
rect 12268 38808 12296 38907
rect 12360 38876 12388 38907
rect 12710 38904 12716 38956
rect 12768 38904 12774 38956
rect 14568 38953 14596 38984
rect 18141 38981 18153 39015
rect 18187 39012 18199 39015
rect 20824 39012 20852 39040
rect 18187 38984 20852 39012
rect 24121 39015 24179 39021
rect 18187 38981 18199 38984
rect 18141 38975 18199 38981
rect 24121 38981 24133 39015
rect 24167 39012 24179 39015
rect 24320 39012 24348 39040
rect 25038 39012 25044 39024
rect 24167 38984 24348 39012
rect 24504 38984 25044 39012
rect 24167 38981 24179 38984
rect 24121 38975 24179 38981
rect 14553 38947 14611 38953
rect 14553 38913 14565 38947
rect 14599 38913 14611 38947
rect 14553 38907 14611 38913
rect 15749 38947 15807 38953
rect 15749 38913 15761 38947
rect 15795 38944 15807 38947
rect 17957 38947 18015 38953
rect 15795 38916 15884 38944
rect 15795 38913 15807 38916
rect 15749 38907 15807 38913
rect 13538 38876 13544 38888
rect 12360 38848 13544 38876
rect 13538 38836 13544 38848
rect 13596 38836 13602 38888
rect 14277 38879 14335 38885
rect 14277 38845 14289 38879
rect 14323 38876 14335 38879
rect 14645 38879 14703 38885
rect 14645 38876 14657 38879
rect 14323 38848 14657 38876
rect 14323 38845 14335 38848
rect 14277 38839 14335 38845
rect 14645 38845 14657 38848
rect 14691 38845 14703 38879
rect 14645 38839 14703 38845
rect 14734 38836 14740 38888
rect 14792 38876 14798 38888
rect 15197 38879 15255 38885
rect 15197 38876 15209 38879
rect 14792 38848 15209 38876
rect 14792 38836 14798 38848
rect 15197 38845 15209 38848
rect 15243 38845 15255 38879
rect 15197 38839 15255 38845
rect 12268 38780 12434 38808
rect 8260 38768 8266 38780
rect 7006 38700 7012 38752
rect 7064 38740 7070 38752
rect 7101 38743 7159 38749
rect 7101 38740 7113 38743
rect 7064 38712 7113 38740
rect 7064 38700 7070 38712
rect 7101 38709 7113 38712
rect 7147 38709 7159 38743
rect 12406 38740 12434 38780
rect 12894 38740 12900 38752
rect 12406 38712 12900 38740
rect 7101 38703 7159 38709
rect 12894 38700 12900 38712
rect 12952 38740 12958 38752
rect 13722 38740 13728 38752
rect 12952 38712 13728 38740
rect 12952 38700 12958 38712
rect 13722 38700 13728 38712
rect 13780 38700 13786 38752
rect 15856 38740 15884 38916
rect 17957 38913 17969 38947
rect 18003 38944 18015 38947
rect 19889 38947 19947 38953
rect 18003 38916 18184 38944
rect 18003 38913 18015 38916
rect 17957 38907 18015 38913
rect 17494 38836 17500 38888
rect 17552 38876 17558 38888
rect 17773 38879 17831 38885
rect 17773 38876 17785 38879
rect 17552 38848 17785 38876
rect 17552 38836 17558 38848
rect 17773 38845 17785 38848
rect 17819 38845 17831 38879
rect 17773 38839 17831 38845
rect 18156 38820 18184 38916
rect 19889 38913 19901 38947
rect 19935 38944 19947 38947
rect 20346 38944 20352 38956
rect 19935 38916 20352 38944
rect 19935 38913 19947 38916
rect 19889 38907 19947 38913
rect 20346 38904 20352 38916
rect 20404 38904 20410 38956
rect 20441 38947 20499 38953
rect 20441 38913 20453 38947
rect 20487 38913 20499 38947
rect 20441 38907 20499 38913
rect 20165 38879 20223 38885
rect 20165 38845 20177 38879
rect 20211 38876 20223 38879
rect 20254 38876 20260 38888
rect 20211 38848 20260 38876
rect 20211 38845 20223 38848
rect 20165 38839 20223 38845
rect 20254 38836 20260 38848
rect 20312 38836 20318 38888
rect 18138 38768 18144 38820
rect 18196 38768 18202 38820
rect 18966 38740 18972 38752
rect 15856 38712 18972 38740
rect 18966 38700 18972 38712
rect 19024 38740 19030 38752
rect 20456 38740 20484 38907
rect 23750 38904 23756 38956
rect 23808 38904 23814 38956
rect 23901 38947 23959 38953
rect 23901 38913 23913 38947
rect 23947 38944 23959 38947
rect 23947 38913 23980 38944
rect 23901 38907 23980 38913
rect 21634 38836 21640 38888
rect 21692 38876 21698 38888
rect 22005 38879 22063 38885
rect 22005 38876 22017 38879
rect 21692 38848 22017 38876
rect 21692 38836 21698 38848
rect 22005 38845 22017 38848
rect 22051 38845 22063 38879
rect 22005 38839 22063 38845
rect 22278 38836 22284 38888
rect 22336 38876 22342 38888
rect 23017 38879 23075 38885
rect 23017 38876 23029 38879
rect 22336 38848 23029 38876
rect 22336 38836 22342 38848
rect 23017 38845 23029 38848
rect 23063 38845 23075 38879
rect 23017 38839 23075 38845
rect 23566 38836 23572 38888
rect 23624 38836 23630 38888
rect 19024 38712 20484 38740
rect 20533 38743 20591 38749
rect 19024 38700 19030 38712
rect 20533 38709 20545 38743
rect 20579 38740 20591 38743
rect 20622 38740 20628 38752
rect 20579 38712 20628 38740
rect 20579 38709 20591 38712
rect 20533 38703 20591 38709
rect 20622 38700 20628 38712
rect 20680 38700 20686 38752
rect 22646 38700 22652 38752
rect 22704 38700 22710 38752
rect 23952 38740 23980 38907
rect 24026 38904 24032 38956
rect 24084 38904 24090 38956
rect 24210 38904 24216 38956
rect 24268 38953 24274 38956
rect 24268 38944 24276 38953
rect 24268 38916 24313 38944
rect 24268 38907 24276 38916
rect 24268 38904 24274 38907
rect 24394 38904 24400 38956
rect 24452 38944 24458 38956
rect 24504 38953 24532 38984
rect 25038 38972 25044 38984
rect 25096 38972 25102 39024
rect 26697 39015 26755 39021
rect 26697 38981 26709 39015
rect 26743 39012 26755 39015
rect 26878 39012 26884 39024
rect 26743 38984 26884 39012
rect 26743 38981 26755 38984
rect 26697 38975 26755 38981
rect 26878 38972 26884 38984
rect 26936 38972 26942 39024
rect 28718 39012 28724 39024
rect 27264 38984 28724 39012
rect 24489 38947 24547 38953
rect 24489 38944 24501 38947
rect 24452 38916 24501 38944
rect 24452 38904 24458 38916
rect 24489 38913 24501 38916
rect 24535 38913 24547 38947
rect 26329 38947 26387 38953
rect 26329 38944 26341 38947
rect 25898 38916 26341 38944
rect 24489 38907 24547 38913
rect 26329 38913 26341 38916
rect 26375 38944 26387 38947
rect 26786 38944 26792 38956
rect 26375 38916 26792 38944
rect 26375 38913 26387 38916
rect 26329 38907 26387 38913
rect 26786 38904 26792 38916
rect 26844 38944 26850 38956
rect 27264 38944 27292 38984
rect 28718 38972 28724 38984
rect 28776 38972 28782 39024
rect 32631 39015 32689 39021
rect 32631 38981 32643 39015
rect 32677 39012 32689 39015
rect 32784 39012 32812 39052
rect 32950 39040 32956 39052
rect 33008 39080 33014 39092
rect 33008 39052 33364 39080
rect 33008 39040 33014 39052
rect 32677 38984 32812 39012
rect 32677 38981 32689 38984
rect 32631 38975 32689 38981
rect 32858 38972 32864 39024
rect 32916 38972 32922 39024
rect 33137 39015 33195 39021
rect 33137 38981 33149 39015
rect 33183 38981 33195 39015
rect 33137 38975 33195 38981
rect 26844 38916 27292 38944
rect 27341 38947 27399 38953
rect 26844 38904 26850 38916
rect 27341 38913 27353 38947
rect 27387 38944 27399 38947
rect 27522 38944 27528 38956
rect 27387 38916 27528 38944
rect 27387 38913 27399 38916
rect 27341 38907 27399 38913
rect 27522 38904 27528 38916
rect 27580 38904 27586 38956
rect 27985 38947 28043 38953
rect 27985 38913 27997 38947
rect 28031 38913 28043 38947
rect 27985 38907 28043 38913
rect 32309 38947 32367 38953
rect 32309 38913 32321 38947
rect 32355 38913 32367 38947
rect 32309 38907 32367 38913
rect 24044 38876 24072 38904
rect 24765 38879 24823 38885
rect 24044 38848 24532 38876
rect 24504 38820 24532 38848
rect 24765 38845 24777 38879
rect 24811 38876 24823 38879
rect 25222 38876 25228 38888
rect 24811 38848 25228 38876
rect 24811 38845 24823 38848
rect 24765 38839 24823 38845
rect 25222 38836 25228 38848
rect 25280 38836 25286 38888
rect 26142 38836 26148 38888
rect 26200 38836 26206 38888
rect 26694 38836 26700 38888
rect 26752 38876 26758 38888
rect 27433 38879 27491 38885
rect 27433 38876 27445 38879
rect 26752 38848 27445 38876
rect 26752 38836 26758 38848
rect 27433 38845 27445 38848
rect 27479 38845 27491 38879
rect 27433 38839 27491 38845
rect 27617 38879 27675 38885
rect 27617 38845 27629 38879
rect 27663 38876 27675 38879
rect 27890 38876 27896 38888
rect 27663 38848 27896 38876
rect 27663 38845 27675 38848
rect 27617 38839 27675 38845
rect 27890 38836 27896 38848
rect 27948 38836 27954 38888
rect 24486 38768 24492 38820
rect 24544 38768 24550 38820
rect 26160 38808 26188 38836
rect 28000 38808 28028 38907
rect 28258 38836 28264 38888
rect 28316 38836 28322 38888
rect 29454 38836 29460 38888
rect 29512 38876 29518 38888
rect 29733 38879 29791 38885
rect 29733 38876 29745 38879
rect 29512 38848 29745 38876
rect 29512 38836 29518 38848
rect 29733 38845 29745 38848
rect 29779 38876 29791 38879
rect 30377 38879 30435 38885
rect 30377 38876 30389 38879
rect 29779 38848 30389 38876
rect 29779 38845 29791 38848
rect 29733 38839 29791 38845
rect 30377 38845 30389 38848
rect 30423 38845 30435 38879
rect 30377 38839 30435 38845
rect 26160 38780 28028 38808
rect 25314 38740 25320 38752
rect 23952 38712 25320 38740
rect 25314 38700 25320 38712
rect 25372 38700 25378 38752
rect 26237 38743 26295 38749
rect 26237 38709 26249 38743
rect 26283 38740 26295 38743
rect 26326 38740 26332 38752
rect 26283 38712 26332 38740
rect 26283 38709 26295 38712
rect 26237 38703 26295 38709
rect 26326 38700 26332 38712
rect 26384 38700 26390 38752
rect 26970 38700 26976 38752
rect 27028 38700 27034 38752
rect 28000 38740 28028 38780
rect 29362 38768 29368 38820
rect 29420 38808 29426 38820
rect 29825 38811 29883 38817
rect 29825 38808 29837 38811
rect 29420 38780 29837 38808
rect 29420 38768 29426 38780
rect 29825 38777 29837 38780
rect 29871 38777 29883 38811
rect 29825 38771 29883 38777
rect 29546 38740 29552 38752
rect 28000 38712 29552 38740
rect 29546 38700 29552 38712
rect 29604 38700 29610 38752
rect 32324 38740 32352 38907
rect 32398 38904 32404 38956
rect 32456 38904 32462 38956
rect 32493 38947 32551 38953
rect 32493 38913 32505 38947
rect 32539 38944 32551 38947
rect 32876 38944 32904 38972
rect 32539 38916 32904 38944
rect 33045 38947 33103 38953
rect 32539 38913 32551 38916
rect 32493 38907 32551 38913
rect 33045 38913 33057 38947
rect 33091 38913 33103 38947
rect 33045 38907 33103 38913
rect 32766 38836 32772 38888
rect 32824 38836 32830 38888
rect 32490 38768 32496 38820
rect 32548 38808 32554 38820
rect 32861 38811 32919 38817
rect 32861 38808 32873 38811
rect 32548 38780 32873 38808
rect 32548 38768 32554 38780
rect 32861 38777 32873 38780
rect 32907 38777 32919 38811
rect 33060 38808 33088 38907
rect 33152 38888 33180 38975
rect 33226 38972 33232 39024
rect 33284 39021 33290 39024
rect 33284 39015 33300 39021
rect 33288 38981 33300 39015
rect 33284 38975 33300 38981
rect 33284 38972 33290 38975
rect 33336 38953 33364 39052
rect 38378 39040 38384 39092
rect 38436 39040 38442 39092
rect 43993 39083 44051 39089
rect 43993 39049 44005 39083
rect 44039 39080 44051 39083
rect 44174 39080 44180 39092
rect 44039 39052 44180 39080
rect 44039 39049 44051 39052
rect 43993 39043 44051 39049
rect 44174 39040 44180 39052
rect 44232 39040 44238 39092
rect 35894 38972 35900 39024
rect 35952 39012 35958 39024
rect 36725 39015 36783 39021
rect 36725 39012 36737 39015
rect 35952 38984 36737 39012
rect 35952 38972 35958 38984
rect 36725 38981 36737 38984
rect 36771 38981 36783 39015
rect 36725 38975 36783 38981
rect 38286 38972 38292 39024
rect 38344 38972 38350 39024
rect 38396 39012 38424 39040
rect 42521 39015 42579 39021
rect 42521 39012 42533 39015
rect 38396 38984 42533 39012
rect 42521 38981 42533 38984
rect 42567 38981 42579 39015
rect 42521 38975 42579 38981
rect 33336 38947 33405 38953
rect 33336 38916 33359 38947
rect 33347 38913 33359 38916
rect 33393 38913 33405 38947
rect 33347 38907 33405 38913
rect 33870 38904 33876 38956
rect 33928 38944 33934 38956
rect 34146 38944 34152 38956
rect 33928 38916 34152 38944
rect 33928 38904 33934 38916
rect 34146 38904 34152 38916
rect 34204 38944 34210 38956
rect 34241 38947 34299 38953
rect 34241 38944 34253 38947
rect 34204 38916 34253 38944
rect 34204 38904 34210 38916
rect 34241 38913 34253 38916
rect 34287 38913 34299 38947
rect 34241 38907 34299 38913
rect 40310 38904 40316 38956
rect 40368 38944 40374 38956
rect 40589 38947 40647 38953
rect 40589 38944 40601 38947
rect 40368 38916 40601 38944
rect 40368 38904 40374 38916
rect 40589 38913 40601 38916
rect 40635 38913 40647 38947
rect 40589 38907 40647 38913
rect 40773 38947 40831 38953
rect 40773 38913 40785 38947
rect 40819 38944 40831 38947
rect 40862 38944 40868 38956
rect 40819 38916 40868 38944
rect 40819 38913 40831 38916
rect 40773 38907 40831 38913
rect 33134 38836 33140 38888
rect 33192 38836 33198 38888
rect 33505 38879 33563 38885
rect 33505 38845 33517 38879
rect 33551 38876 33563 38879
rect 33689 38879 33747 38885
rect 33689 38876 33701 38879
rect 33551 38848 33701 38876
rect 33551 38845 33563 38848
rect 33505 38839 33563 38845
rect 33689 38845 33701 38848
rect 33735 38845 33747 38879
rect 33689 38839 33747 38845
rect 36541 38879 36599 38885
rect 36541 38845 36553 38879
rect 36587 38876 36599 38879
rect 36722 38876 36728 38888
rect 36587 38848 36728 38876
rect 36587 38845 36599 38848
rect 36541 38839 36599 38845
rect 36722 38836 36728 38848
rect 36780 38836 36786 38888
rect 38102 38836 38108 38888
rect 38160 38876 38166 38888
rect 38749 38879 38807 38885
rect 38749 38876 38761 38879
rect 38160 38848 38761 38876
rect 38160 38836 38166 38848
rect 38749 38845 38761 38848
rect 38795 38845 38807 38879
rect 38749 38839 38807 38845
rect 39025 38879 39083 38885
rect 39025 38845 39037 38879
rect 39071 38876 39083 38879
rect 39850 38876 39856 38888
rect 39071 38848 39856 38876
rect 39071 38845 39083 38848
rect 39025 38839 39083 38845
rect 39850 38836 39856 38848
rect 39908 38836 39914 38888
rect 40126 38836 40132 38888
rect 40184 38876 40190 38888
rect 40788 38876 40816 38907
rect 40862 38904 40868 38916
rect 40920 38904 40926 38956
rect 40184 38848 40816 38876
rect 40184 38836 40190 38848
rect 33594 38808 33600 38820
rect 33060 38780 33600 38808
rect 32861 38771 32919 38777
rect 33594 38768 33600 38780
rect 33652 38768 33658 38820
rect 36906 38768 36912 38820
rect 36964 38808 36970 38820
rect 37001 38811 37059 38817
rect 37001 38808 37013 38811
rect 36964 38780 37013 38808
rect 36964 38768 36970 38780
rect 37001 38777 37013 38780
rect 37047 38808 37059 38811
rect 37047 38780 37780 38808
rect 37047 38777 37059 38780
rect 37001 38771 37059 38777
rect 33226 38740 33232 38752
rect 32324 38712 33232 38740
rect 33226 38700 33232 38712
rect 33284 38700 33290 38752
rect 35894 38700 35900 38752
rect 35952 38700 35958 38752
rect 37274 38700 37280 38752
rect 37332 38700 37338 38752
rect 37752 38740 37780 38780
rect 40310 38768 40316 38820
rect 40368 38808 40374 38820
rect 40589 38811 40647 38817
rect 40589 38808 40601 38811
rect 40368 38780 40601 38808
rect 40368 38768 40374 38780
rect 40589 38777 40601 38780
rect 40635 38777 40647 38811
rect 40589 38771 40647 38777
rect 38286 38740 38292 38752
rect 37752 38712 38292 38740
rect 38286 38700 38292 38712
rect 38344 38700 38350 38752
rect 40218 38700 40224 38752
rect 40276 38740 40282 38752
rect 40497 38743 40555 38749
rect 40497 38740 40509 38743
rect 40276 38712 40509 38740
rect 40276 38700 40282 38712
rect 40497 38709 40509 38712
rect 40543 38709 40555 38743
rect 40497 38703 40555 38709
rect 1104 38650 44620 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 44620 38650
rect 1104 38576 44620 38598
rect 8386 38536 8392 38548
rect 7852 38508 8392 38536
rect 6457 38403 6515 38409
rect 6457 38369 6469 38403
rect 6503 38400 6515 38403
rect 6730 38400 6736 38412
rect 6503 38372 6736 38400
rect 6503 38369 6515 38372
rect 6457 38363 6515 38369
rect 6730 38360 6736 38372
rect 6788 38360 6794 38412
rect 7852 38318 7880 38508
rect 8386 38496 8392 38508
rect 8444 38536 8450 38548
rect 9582 38536 9588 38548
rect 8444 38508 9588 38536
rect 8444 38496 8450 38508
rect 9582 38496 9588 38508
rect 9640 38496 9646 38548
rect 13633 38539 13691 38545
rect 13633 38505 13645 38539
rect 13679 38536 13691 38539
rect 14734 38536 14740 38548
rect 13679 38508 14740 38536
rect 13679 38505 13691 38508
rect 13633 38499 13691 38505
rect 14734 38496 14740 38508
rect 14792 38496 14798 38548
rect 23566 38496 23572 38548
rect 23624 38496 23630 38548
rect 28258 38496 28264 38548
rect 28316 38536 28322 38548
rect 28353 38539 28411 38545
rect 28353 38536 28365 38539
rect 28316 38508 28365 38536
rect 28316 38496 28322 38508
rect 28353 38505 28365 38508
rect 28399 38505 28411 38539
rect 28353 38499 28411 38505
rect 29362 38496 29368 38548
rect 29420 38496 29426 38548
rect 32398 38496 32404 38548
rect 32456 38536 32462 38548
rect 32677 38539 32735 38545
rect 32677 38536 32689 38539
rect 32456 38508 32689 38536
rect 32456 38496 32462 38508
rect 32677 38505 32689 38508
rect 32723 38505 32735 38539
rect 32677 38499 32735 38505
rect 33226 38496 33232 38548
rect 33284 38496 33290 38548
rect 33594 38496 33600 38548
rect 33652 38536 33658 38548
rect 33689 38539 33747 38545
rect 33689 38536 33701 38539
rect 33652 38508 33701 38536
rect 33652 38496 33658 38508
rect 33689 38505 33701 38508
rect 33735 38505 33747 38539
rect 33689 38499 33747 38505
rect 40862 38496 40868 38548
rect 40920 38536 40926 38548
rect 41601 38539 41659 38545
rect 41601 38536 41613 38539
rect 40920 38508 41613 38536
rect 40920 38496 40926 38508
rect 41601 38505 41613 38508
rect 41647 38505 41659 38539
rect 41601 38499 41659 38505
rect 42518 38496 42524 38548
rect 42576 38496 42582 38548
rect 9309 38471 9367 38477
rect 9309 38437 9321 38471
rect 9355 38468 9367 38471
rect 12710 38468 12716 38480
rect 9355 38440 12716 38468
rect 9355 38437 9367 38440
rect 9309 38431 9367 38437
rect 8205 38403 8263 38409
rect 8205 38369 8217 38403
rect 8251 38400 8263 38403
rect 8941 38403 8999 38409
rect 8941 38400 8953 38403
rect 8251 38372 8953 38400
rect 8251 38369 8263 38372
rect 8205 38363 8263 38369
rect 8941 38369 8953 38372
rect 8987 38400 8999 38403
rect 9030 38400 9036 38412
rect 8987 38372 9036 38400
rect 8987 38369 8999 38372
rect 8941 38363 8999 38369
rect 9030 38360 9036 38372
rect 9088 38360 9094 38412
rect 9125 38335 9183 38341
rect 9125 38301 9137 38335
rect 9171 38332 9183 38335
rect 9324 38332 9352 38431
rect 12710 38428 12716 38440
rect 12768 38428 12774 38480
rect 25038 38428 25044 38480
rect 25096 38428 25102 38480
rect 29380 38468 29408 38496
rect 33134 38468 33140 38480
rect 29012 38440 29408 38468
rect 33060 38440 33140 38468
rect 9401 38403 9459 38409
rect 9401 38369 9413 38403
rect 9447 38400 9459 38403
rect 10505 38403 10563 38409
rect 10505 38400 10517 38403
rect 9447 38372 10517 38400
rect 9447 38369 9459 38372
rect 9401 38363 9459 38369
rect 10505 38369 10517 38372
rect 10551 38369 10563 38403
rect 15473 38403 15531 38409
rect 10505 38363 10563 38369
rect 12544 38372 13308 38400
rect 12544 38344 12572 38372
rect 9585 38335 9643 38341
rect 9585 38332 9597 38335
rect 9171 38304 9260 38332
rect 9324 38304 9597 38332
rect 9171 38301 9183 38304
rect 9125 38295 9183 38301
rect 9232 38276 9260 38304
rect 9585 38301 9597 38304
rect 9631 38301 9643 38335
rect 9585 38295 9643 38301
rect 9674 38292 9680 38344
rect 9732 38332 9738 38344
rect 9861 38335 9919 38341
rect 9861 38332 9873 38335
rect 9732 38304 9873 38332
rect 9732 38292 9738 38304
rect 9861 38301 9873 38304
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 11422 38292 11428 38344
rect 11480 38292 11486 38344
rect 12526 38292 12532 38344
rect 12584 38292 12590 38344
rect 12894 38292 12900 38344
rect 12952 38332 12958 38344
rect 13280 38341 13308 38372
rect 15473 38369 15485 38403
rect 15519 38400 15531 38403
rect 16485 38403 16543 38409
rect 16485 38400 16497 38403
rect 15519 38372 16497 38400
rect 15519 38369 15531 38372
rect 15473 38363 15531 38369
rect 16485 38369 16497 38372
rect 16531 38369 16543 38403
rect 18233 38403 18291 38409
rect 18233 38400 18245 38403
rect 16485 38363 16543 38369
rect 16960 38372 18245 38400
rect 16960 38344 16988 38372
rect 18233 38369 18245 38372
rect 18279 38400 18291 38403
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 18279 38372 19993 38400
rect 18279 38369 18291 38372
rect 18233 38363 18291 38369
rect 19981 38369 19993 38372
rect 20027 38400 20039 38403
rect 20714 38400 20720 38412
rect 20027 38372 20720 38400
rect 20027 38369 20039 38372
rect 19981 38363 20039 38369
rect 20714 38360 20720 38372
rect 20772 38400 20778 38412
rect 21821 38403 21879 38409
rect 21821 38400 21833 38403
rect 20772 38372 21833 38400
rect 20772 38360 20778 38372
rect 21821 38369 21833 38372
rect 21867 38369 21879 38403
rect 21821 38363 21879 38369
rect 22094 38360 22100 38412
rect 22152 38360 22158 38412
rect 25056 38400 25084 38428
rect 25406 38400 25412 38412
rect 25056 38372 25412 38400
rect 25406 38360 25412 38372
rect 25464 38360 25470 38412
rect 28902 38360 28908 38412
rect 28960 38360 28966 38412
rect 29012 38409 29040 38440
rect 28997 38403 29055 38409
rect 28997 38369 29009 38403
rect 29043 38369 29055 38403
rect 28997 38363 29055 38369
rect 29546 38360 29552 38412
rect 29604 38400 29610 38412
rect 29641 38403 29699 38409
rect 29641 38400 29653 38403
rect 29604 38372 29653 38400
rect 29604 38360 29610 38372
rect 29641 38369 29653 38372
rect 29687 38369 29699 38403
rect 29641 38363 29699 38369
rect 31389 38403 31447 38409
rect 31389 38369 31401 38403
rect 31435 38400 31447 38403
rect 31570 38400 31576 38412
rect 31435 38372 31576 38400
rect 31435 38369 31447 38372
rect 31389 38363 31447 38369
rect 31570 38360 31576 38372
rect 31628 38400 31634 38412
rect 32033 38403 32091 38409
rect 32033 38400 32045 38403
rect 31628 38372 32045 38400
rect 31628 38360 31634 38372
rect 32033 38369 32045 38372
rect 32079 38369 32091 38403
rect 32033 38363 32091 38369
rect 12989 38335 13047 38341
rect 12989 38332 13001 38335
rect 12952 38304 13001 38332
rect 12952 38292 12958 38304
rect 12989 38301 13001 38304
rect 13035 38301 13047 38335
rect 12989 38295 13047 38301
rect 13137 38335 13195 38341
rect 13137 38301 13149 38335
rect 13183 38332 13195 38335
rect 13265 38335 13323 38341
rect 13183 38301 13216 38332
rect 13137 38295 13216 38301
rect 13265 38301 13277 38335
rect 13311 38301 13323 38335
rect 13265 38295 13323 38301
rect 6733 38267 6791 38273
rect 6733 38233 6745 38267
rect 6779 38264 6791 38267
rect 7006 38264 7012 38276
rect 6779 38236 7012 38264
rect 6779 38233 6791 38236
rect 6733 38227 6791 38233
rect 7006 38224 7012 38236
rect 7064 38224 7070 38276
rect 9214 38224 9220 38276
rect 9272 38224 9278 38276
rect 9769 38267 9827 38273
rect 9769 38233 9781 38267
rect 9815 38264 9827 38267
rect 10870 38264 10876 38276
rect 9815 38236 10876 38264
rect 9815 38233 9827 38236
rect 9769 38227 9827 38233
rect 10870 38224 10876 38236
rect 10928 38224 10934 38276
rect 9950 38156 9956 38208
rect 10008 38156 10014 38208
rect 13188 38196 13216 38295
rect 13354 38292 13360 38344
rect 13412 38292 13418 38344
rect 13495 38335 13553 38341
rect 13495 38301 13507 38335
rect 13541 38332 13553 38335
rect 13722 38332 13728 38344
rect 13541 38304 13728 38332
rect 13541 38301 13553 38304
rect 13495 38295 13553 38301
rect 13722 38292 13728 38304
rect 13780 38292 13786 38344
rect 16942 38292 16948 38344
rect 17000 38292 17006 38344
rect 18874 38292 18880 38344
rect 18932 38292 18938 38344
rect 28534 38292 28540 38344
rect 28592 38292 28598 38344
rect 28920 38332 28948 38360
rect 29089 38335 29147 38341
rect 29089 38332 29101 38335
rect 28920 38304 29101 38332
rect 29089 38301 29101 38304
rect 29135 38301 29147 38335
rect 29089 38295 29147 38301
rect 29273 38335 29331 38341
rect 29273 38301 29285 38335
rect 29319 38332 29331 38335
rect 29454 38332 29460 38344
rect 29319 38304 29460 38332
rect 29319 38301 29331 38304
rect 29273 38295 29331 38301
rect 29454 38292 29460 38304
rect 29512 38292 29518 38344
rect 32861 38335 32919 38341
rect 32861 38301 32873 38335
rect 32907 38301 32919 38335
rect 33060 38332 33088 38440
rect 33134 38428 33140 38440
rect 33192 38468 33198 38480
rect 42536 38468 42564 38496
rect 33192 38440 33364 38468
rect 33192 38428 33198 38440
rect 33137 38335 33195 38341
rect 33137 38332 33149 38335
rect 33060 38304 33149 38332
rect 32861 38295 32919 38301
rect 33137 38301 33149 38304
rect 33183 38301 33195 38335
rect 33137 38295 33195 38301
rect 15286 38224 15292 38276
rect 15344 38264 15350 38276
rect 16482 38264 16488 38276
rect 15344 38236 16488 38264
rect 15344 38224 15350 38236
rect 16482 38224 16488 38236
rect 16540 38264 16546 38276
rect 16540 38236 16790 38264
rect 16540 38224 16546 38236
rect 17954 38224 17960 38276
rect 18012 38224 18018 38276
rect 20254 38224 20260 38276
rect 20312 38224 20318 38276
rect 20640 38236 20746 38264
rect 20640 38208 20668 38236
rect 22554 38224 22560 38276
rect 22612 38224 22618 38276
rect 27154 38224 27160 38276
rect 27212 38224 27218 38276
rect 28626 38224 28632 38276
rect 28684 38224 28690 38276
rect 28721 38267 28779 38273
rect 28721 38233 28733 38267
rect 28767 38233 28779 38267
rect 28721 38227 28779 38233
rect 28859 38267 28917 38273
rect 28859 38233 28871 38267
rect 28905 38264 28917 38267
rect 28905 38236 29868 38264
rect 28905 38233 28917 38236
rect 28859 38227 28917 38233
rect 14829 38199 14887 38205
rect 14829 38196 14841 38199
rect 13188 38168 14841 38196
rect 14829 38165 14841 38168
rect 14875 38196 14887 38199
rect 17310 38196 17316 38208
rect 14875 38168 17316 38196
rect 14875 38165 14887 38168
rect 14829 38159 14887 38165
rect 17310 38156 17316 38168
rect 17368 38156 17374 38208
rect 17770 38156 17776 38208
rect 17828 38196 17834 38208
rect 18325 38199 18383 38205
rect 18325 38196 18337 38199
rect 17828 38168 18337 38196
rect 17828 38156 17834 38168
rect 18325 38165 18337 38168
rect 18371 38165 18383 38199
rect 18325 38159 18383 38165
rect 20622 38156 20628 38208
rect 20680 38156 20686 38208
rect 21634 38156 21640 38208
rect 21692 38196 21698 38208
rect 21729 38199 21787 38205
rect 21729 38196 21741 38199
rect 21692 38168 21741 38196
rect 21692 38156 21698 38168
rect 21729 38165 21741 38168
rect 21775 38165 21787 38199
rect 28736 38196 28764 38227
rect 29181 38199 29239 38205
rect 29181 38196 29193 38199
rect 28736 38168 29193 38196
rect 21729 38159 21787 38165
rect 29181 38165 29193 38168
rect 29227 38165 29239 38199
rect 29840 38196 29868 38236
rect 29914 38224 29920 38276
rect 29972 38224 29978 38276
rect 30374 38224 30380 38276
rect 30432 38224 30438 38276
rect 32876 38264 32904 38295
rect 33226 38292 33232 38344
rect 33284 38292 33290 38344
rect 33336 38341 33364 38440
rect 41386 38440 42564 38468
rect 33502 38360 33508 38412
rect 33560 38400 33566 38412
rect 38013 38403 38071 38409
rect 38013 38400 38025 38403
rect 33560 38372 33824 38400
rect 33560 38360 33566 38372
rect 33321 38335 33379 38341
rect 33321 38301 33333 38335
rect 33367 38301 33379 38335
rect 33321 38295 33379 38301
rect 33410 38292 33416 38344
rect 33468 38332 33474 38344
rect 33796 38341 33824 38372
rect 37292 38372 38025 38400
rect 37292 38344 37320 38372
rect 38013 38369 38025 38372
rect 38059 38369 38071 38403
rect 38013 38363 38071 38369
rect 38286 38360 38292 38412
rect 38344 38400 38350 38412
rect 38344 38372 41276 38400
rect 38344 38360 38350 38372
rect 33597 38335 33655 38341
rect 33597 38332 33609 38335
rect 33468 38304 33609 38332
rect 33468 38292 33474 38304
rect 33597 38301 33609 38304
rect 33643 38301 33655 38335
rect 33597 38295 33655 38301
rect 33781 38335 33839 38341
rect 33781 38301 33793 38335
rect 33827 38301 33839 38335
rect 33781 38295 33839 38301
rect 34790 38292 34796 38344
rect 34848 38332 34854 38344
rect 34977 38335 35035 38341
rect 34977 38332 34989 38335
rect 34848 38304 34989 38332
rect 34848 38292 34854 38304
rect 34977 38301 34989 38304
rect 35023 38301 35035 38335
rect 36906 38332 36912 38344
rect 36386 38304 36912 38332
rect 34977 38295 35035 38301
rect 36906 38292 36912 38304
rect 36964 38292 36970 38344
rect 37274 38292 37280 38344
rect 37332 38292 37338 38344
rect 37366 38292 37372 38344
rect 37424 38332 37430 38344
rect 37737 38335 37795 38341
rect 37737 38332 37749 38335
rect 37424 38304 37749 38332
rect 37424 38292 37430 38304
rect 37737 38301 37749 38304
rect 37783 38301 37795 38335
rect 37737 38295 37795 38301
rect 37918 38292 37924 38344
rect 37976 38292 37982 38344
rect 39850 38292 39856 38344
rect 39908 38292 39914 38344
rect 41248 38332 41276 38372
rect 41386 38332 41414 38440
rect 42702 38360 42708 38412
rect 42760 38360 42766 38412
rect 42794 38360 42800 38412
rect 42852 38400 42858 38412
rect 43441 38403 43499 38409
rect 43441 38400 43453 38403
rect 42852 38372 43453 38400
rect 42852 38360 42858 38372
rect 43441 38369 43453 38372
rect 43487 38369 43499 38403
rect 43441 38363 43499 38369
rect 41248 38318 41414 38332
rect 41262 38304 41414 38318
rect 42610 38292 42616 38344
rect 42668 38292 42674 38344
rect 43254 38292 43260 38344
rect 43312 38292 43318 38344
rect 33505 38267 33563 38273
rect 33505 38264 33517 38267
rect 32876 38236 33517 38264
rect 33505 38233 33517 38236
rect 33551 38264 33563 38267
rect 33870 38264 33876 38276
rect 33551 38236 33876 38264
rect 33551 38233 33563 38236
rect 33505 38227 33563 38233
rect 33870 38224 33876 38236
rect 33928 38224 33934 38276
rect 35250 38224 35256 38276
rect 35308 38224 35314 38276
rect 37829 38267 37887 38273
rect 37829 38233 37841 38267
rect 37875 38264 37887 38267
rect 40034 38264 40040 38276
rect 37875 38236 40040 38264
rect 37875 38233 37887 38236
rect 37829 38227 37887 38233
rect 40034 38224 40040 38236
rect 40092 38224 40098 38276
rect 40126 38224 40132 38276
rect 40184 38224 40190 38276
rect 43073 38267 43131 38273
rect 43073 38264 43085 38267
rect 42168 38236 43085 38264
rect 42168 38208 42196 38236
rect 43073 38233 43085 38236
rect 43119 38233 43131 38267
rect 43073 38227 43131 38233
rect 30098 38196 30104 38208
rect 29840 38168 30104 38196
rect 29181 38159 29239 38165
rect 30098 38156 30104 38168
rect 30156 38156 30162 38208
rect 31478 38156 31484 38208
rect 31536 38156 31542 38208
rect 33045 38199 33103 38205
rect 33045 38165 33057 38199
rect 33091 38196 33103 38199
rect 33226 38196 33232 38208
rect 33091 38168 33232 38196
rect 33091 38165 33103 38168
rect 33045 38159 33103 38165
rect 33226 38156 33232 38168
rect 33284 38156 33290 38208
rect 36722 38156 36728 38208
rect 36780 38156 36786 38208
rect 38654 38156 38660 38208
rect 38712 38156 38718 38208
rect 42150 38156 42156 38208
rect 42208 38156 42214 38208
rect 42978 38156 42984 38208
rect 43036 38156 43042 38208
rect 1104 38106 44620 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 44620 38106
rect 1104 38032 44620 38054
rect 9950 37992 9956 38004
rect 9692 37964 9956 37992
rect 6730 37924 6736 37936
rect 6564 37896 6736 37924
rect 6564 37865 6592 37896
rect 6730 37884 6736 37896
rect 6788 37884 6794 37936
rect 8386 37924 8392 37936
rect 8050 37896 8392 37924
rect 8386 37884 8392 37896
rect 8444 37884 8450 37936
rect 9692 37933 9720 37964
rect 9950 37952 9956 37964
rect 10008 37952 10014 38004
rect 11149 37995 11207 38001
rect 11149 37961 11161 37995
rect 11195 37992 11207 37995
rect 11422 37992 11428 38004
rect 11195 37964 11428 37992
rect 11195 37961 11207 37964
rect 11149 37955 11207 37961
rect 11422 37952 11428 37964
rect 11480 37952 11486 38004
rect 13722 37952 13728 38004
rect 13780 37992 13786 38004
rect 13780 37964 16712 37992
rect 13780 37952 13786 37964
rect 9677 37927 9735 37933
rect 9677 37893 9689 37927
rect 9723 37893 9735 37927
rect 9677 37887 9735 37893
rect 15286 37884 15292 37936
rect 15344 37884 15350 37936
rect 6549 37859 6607 37865
rect 6549 37825 6561 37859
rect 6595 37825 6607 37859
rect 6549 37819 6607 37825
rect 9398 37816 9404 37868
rect 9456 37816 9462 37868
rect 10962 37856 10968 37868
rect 10810 37828 10968 37856
rect 10962 37816 10968 37828
rect 11020 37816 11026 37868
rect 12894 37816 12900 37868
rect 12952 37856 12958 37868
rect 13173 37859 13231 37865
rect 13173 37856 13185 37859
rect 12952 37828 13185 37856
rect 12952 37816 12958 37828
rect 13173 37825 13185 37828
rect 13219 37825 13231 37859
rect 13173 37819 13231 37825
rect 13354 37816 13360 37868
rect 13412 37816 13418 37868
rect 13449 37859 13507 37865
rect 13449 37825 13461 37859
rect 13495 37825 13507 37859
rect 13449 37819 13507 37825
rect 6825 37791 6883 37797
rect 6825 37757 6837 37791
rect 6871 37788 6883 37791
rect 6914 37788 6920 37800
rect 6871 37760 6920 37788
rect 6871 37757 6883 37760
rect 6825 37751 6883 37757
rect 6914 37748 6920 37760
rect 6972 37748 6978 37800
rect 8297 37791 8355 37797
rect 8297 37757 8309 37791
rect 8343 37788 8355 37791
rect 8938 37788 8944 37800
rect 8343 37760 8944 37788
rect 8343 37757 8355 37760
rect 8297 37751 8355 37757
rect 8938 37748 8944 37760
rect 8996 37748 9002 37800
rect 8386 37612 8392 37664
rect 8444 37612 8450 37664
rect 12986 37612 12992 37664
rect 13044 37612 13050 37664
rect 13464 37652 13492 37819
rect 13998 37748 14004 37800
rect 14056 37788 14062 37800
rect 14277 37791 14335 37797
rect 14277 37788 14289 37791
rect 14056 37760 14289 37788
rect 14056 37748 14062 37760
rect 14277 37757 14289 37760
rect 14323 37757 14335 37791
rect 14277 37751 14335 37757
rect 14553 37791 14611 37797
rect 14553 37757 14565 37791
rect 14599 37788 14611 37791
rect 15286 37788 15292 37800
rect 14599 37760 15292 37788
rect 14599 37757 14611 37760
rect 14553 37751 14611 37757
rect 15286 37748 15292 37760
rect 15344 37748 15350 37800
rect 16684 37788 16712 37964
rect 17770 37952 17776 38004
rect 17828 37952 17834 38004
rect 17954 37952 17960 38004
rect 18012 37992 18018 38004
rect 18509 37995 18567 38001
rect 18509 37992 18521 37995
rect 18012 37964 18521 37992
rect 18012 37952 18018 37964
rect 18509 37961 18521 37964
rect 18555 37961 18567 37995
rect 19242 37992 19248 38004
rect 18509 37955 18567 37961
rect 18800 37964 19248 37992
rect 17788 37924 17816 37952
rect 18800 37924 18828 37964
rect 19242 37952 19248 37964
rect 19300 37952 19306 38004
rect 20254 37952 20260 38004
rect 20312 37992 20318 38004
rect 21177 37995 21235 38001
rect 21177 37992 21189 37995
rect 20312 37964 21189 37992
rect 20312 37952 20318 37964
rect 21177 37961 21189 37964
rect 21223 37961 21235 37995
rect 21177 37955 21235 37961
rect 21821 37995 21879 38001
rect 21821 37961 21833 37995
rect 21867 37961 21879 37995
rect 21821 37955 21879 37961
rect 22189 37995 22247 38001
rect 22189 37961 22201 37995
rect 22235 37992 22247 37995
rect 22646 37992 22652 38004
rect 22235 37964 22652 37992
rect 22235 37961 22247 37964
rect 22189 37955 22247 37961
rect 17236 37896 17816 37924
rect 17880 37896 18828 37924
rect 17034 37816 17040 37868
rect 17092 37816 17098 37868
rect 17236 37865 17264 37896
rect 17185 37859 17264 37865
rect 17185 37825 17197 37859
rect 17231 37828 17264 37859
rect 17231 37825 17243 37828
rect 17185 37819 17243 37825
rect 17310 37816 17316 37868
rect 17368 37816 17374 37868
rect 17402 37816 17408 37868
rect 17460 37816 17466 37868
rect 17541 37859 17599 37865
rect 17541 37825 17553 37859
rect 17587 37856 17599 37859
rect 17880 37856 17908 37896
rect 17587 37828 17908 37856
rect 17587 37825 17599 37828
rect 17541 37819 17599 37825
rect 17558 37788 17586 37819
rect 18506 37816 18512 37868
rect 18564 37856 18570 37868
rect 20349 37859 20407 37865
rect 18564 37842 18998 37856
rect 18564 37828 19012 37842
rect 18564 37816 18570 37828
rect 16684 37760 17586 37788
rect 17865 37791 17923 37797
rect 17865 37757 17877 37791
rect 17911 37757 17923 37791
rect 17865 37751 17923 37757
rect 16666 37720 16672 37732
rect 15948 37692 16672 37720
rect 15948 37652 15976 37692
rect 16666 37680 16672 37692
rect 16724 37680 16730 37732
rect 17681 37723 17739 37729
rect 17681 37689 17693 37723
rect 17727 37720 17739 37723
rect 17880 37720 17908 37751
rect 17727 37692 17908 37720
rect 17727 37689 17739 37692
rect 17681 37683 17739 37689
rect 13464 37624 15976 37652
rect 16022 37612 16028 37664
rect 16080 37612 16086 37664
rect 18601 37655 18659 37661
rect 18601 37621 18613 37655
rect 18647 37652 18659 37655
rect 18874 37652 18880 37664
rect 18647 37624 18880 37652
rect 18647 37621 18659 37624
rect 18601 37615 18659 37621
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 18984 37652 19012 37828
rect 20349 37825 20361 37859
rect 20395 37856 20407 37859
rect 20714 37856 20720 37868
rect 20395 37828 20720 37856
rect 20395 37825 20407 37828
rect 20349 37819 20407 37825
rect 20714 37816 20720 37828
rect 20772 37816 20778 37868
rect 21361 37859 21419 37865
rect 21361 37825 21373 37859
rect 21407 37856 21419 37859
rect 21836 37856 21864 37955
rect 22646 37952 22652 37964
rect 22704 37952 22710 38004
rect 24854 37952 24860 38004
rect 24912 37992 24918 38004
rect 25225 37995 25283 38001
rect 25225 37992 25237 37995
rect 24912 37964 25237 37992
rect 24912 37952 24918 37964
rect 25225 37961 25237 37964
rect 25271 37992 25283 37995
rect 27522 37992 27528 38004
rect 25271 37964 27528 37992
rect 25271 37961 25283 37964
rect 25225 37955 25283 37961
rect 27522 37952 27528 37964
rect 27580 37952 27586 38004
rect 28644 37964 29408 37992
rect 22278 37884 22284 37936
rect 22336 37884 22342 37936
rect 27706 37924 27712 37936
rect 27172 37896 27712 37924
rect 21407 37828 21864 37856
rect 24765 37859 24823 37865
rect 21407 37825 21419 37828
rect 21361 37819 21419 37825
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25314 37856 25320 37868
rect 24811 37828 25320 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25314 37816 25320 37828
rect 25372 37816 25378 37868
rect 27172 37865 27200 37896
rect 27706 37884 27712 37896
rect 27764 37884 27770 37936
rect 27157 37859 27215 37865
rect 27157 37825 27169 37859
rect 27203 37825 27215 37859
rect 27157 37819 27215 37825
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 27341 37859 27399 37865
rect 27341 37825 27353 37859
rect 27387 37825 27399 37859
rect 27341 37819 27399 37825
rect 20073 37791 20131 37797
rect 20073 37757 20085 37791
rect 20119 37788 20131 37791
rect 20441 37791 20499 37797
rect 20441 37788 20453 37791
rect 20119 37760 20453 37788
rect 20119 37757 20131 37760
rect 20073 37751 20131 37757
rect 20441 37757 20453 37760
rect 20487 37757 20499 37791
rect 20441 37751 20499 37757
rect 20990 37748 20996 37800
rect 21048 37748 21054 37800
rect 22370 37748 22376 37800
rect 22428 37748 22434 37800
rect 24581 37723 24639 37729
rect 24581 37689 24593 37723
rect 24627 37720 24639 37723
rect 24762 37720 24768 37732
rect 24627 37692 24768 37720
rect 24627 37689 24639 37692
rect 24581 37683 24639 37689
rect 24762 37680 24768 37692
rect 24820 37720 24826 37732
rect 27264 37720 27292 37819
rect 27356 37788 27384 37819
rect 27430 37816 27436 37868
rect 27488 37865 27494 37868
rect 28644 37865 28672 37964
rect 28718 37884 28724 37936
rect 28776 37924 28782 37936
rect 29380 37933 29408 37964
rect 29914 37952 29920 38004
rect 29972 37992 29978 38004
rect 30561 37995 30619 38001
rect 30561 37992 30573 37995
rect 29972 37964 30573 37992
rect 29972 37952 29978 37964
rect 30561 37961 30573 37964
rect 30607 37961 30619 37995
rect 30561 37955 30619 37961
rect 33134 37952 33140 38004
rect 33192 37952 33198 38004
rect 35526 37952 35532 38004
rect 35584 37952 35590 38004
rect 35621 37995 35679 38001
rect 35621 37961 35633 37995
rect 35667 37992 35679 37995
rect 35667 37964 36308 37992
rect 35667 37961 35679 37964
rect 35621 37955 35679 37961
rect 29149 37927 29207 37933
rect 29149 37924 29161 37927
rect 28776 37896 29161 37924
rect 28776 37884 28782 37896
rect 27488 37859 27517 37865
rect 27505 37825 27517 37859
rect 28629 37859 28687 37865
rect 28629 37856 28641 37859
rect 27488 37819 27517 37825
rect 28276 37828 28641 37856
rect 27488 37816 27494 37819
rect 27617 37791 27675 37797
rect 27356 37760 27476 37788
rect 24820 37692 27292 37720
rect 27448 37720 27476 37760
rect 27617 37757 27629 37791
rect 27663 37788 27675 37791
rect 27709 37791 27767 37797
rect 27709 37788 27721 37791
rect 27663 37760 27721 37788
rect 27663 37757 27675 37760
rect 27617 37751 27675 37757
rect 27709 37757 27721 37760
rect 27755 37757 27767 37791
rect 27709 37751 27767 37757
rect 27798 37748 27804 37800
rect 27856 37788 27862 37800
rect 28276 37797 28304 37828
rect 28629 37825 28641 37828
rect 28675 37825 28687 37859
rect 28629 37819 28687 37825
rect 28813 37859 28871 37865
rect 28813 37825 28825 37859
rect 28859 37825 28871 37859
rect 28813 37819 28871 37825
rect 28905 37859 28963 37865
rect 28905 37825 28917 37859
rect 28951 37856 28963 37859
rect 29012 37856 29040 37896
rect 29149 37893 29161 37896
rect 29195 37893 29207 37927
rect 29149 37887 29207 37893
rect 29365 37927 29423 37933
rect 29365 37893 29377 37927
rect 29411 37893 29423 37927
rect 31047 37927 31105 37933
rect 31047 37924 31059 37927
rect 29365 37887 29423 37893
rect 30116 37896 31059 37924
rect 30116 37868 30144 37896
rect 31047 37893 31059 37896
rect 31093 37924 31105 37927
rect 32950 37924 32956 37936
rect 31093 37896 32956 37924
rect 31093 37893 31105 37896
rect 31047 37887 31105 37893
rect 32950 37884 32956 37896
rect 33008 37884 33014 37936
rect 35544 37924 35572 37952
rect 36280 37933 36308 37964
rect 37918 37952 37924 38004
rect 37976 37992 37982 38004
rect 38013 37995 38071 38001
rect 38013 37992 38025 37995
rect 37976 37964 38025 37992
rect 37976 37952 37982 37964
rect 38013 37961 38025 37964
rect 38059 37961 38071 37995
rect 38013 37955 38071 37961
rect 38654 37952 38660 38004
rect 38712 37952 38718 38004
rect 38746 37952 38752 38004
rect 38804 37992 38810 38004
rect 38841 37995 38899 38001
rect 38841 37992 38853 37995
rect 38804 37964 38853 37992
rect 38804 37952 38810 37964
rect 38841 37961 38853 37964
rect 38887 37961 38899 37995
rect 38841 37955 38899 37961
rect 40126 37952 40132 38004
rect 40184 37992 40190 38004
rect 40221 37995 40279 38001
rect 40221 37992 40233 37995
rect 40184 37964 40233 37992
rect 40184 37952 40190 37964
rect 40221 37961 40233 37964
rect 40267 37961 40279 37995
rect 40221 37955 40279 37961
rect 42610 37952 42616 38004
rect 42668 37952 42674 38004
rect 42978 37952 42984 38004
rect 43036 37952 43042 38004
rect 36049 37927 36107 37933
rect 36049 37924 36061 37927
rect 35544 37896 36061 37924
rect 28951 37828 29040 37856
rect 28951 37825 28963 37828
rect 28905 37819 28963 37825
rect 28261 37791 28319 37797
rect 28261 37788 28273 37791
rect 27856 37760 28273 37788
rect 27856 37748 27862 37760
rect 28261 37757 28273 37760
rect 28307 37757 28319 37791
rect 28828 37788 28856 37819
rect 30098 37816 30104 37868
rect 30156 37816 30162 37868
rect 30745 37859 30803 37865
rect 30745 37825 30757 37859
rect 30791 37825 30803 37859
rect 30745 37819 30803 37825
rect 30837 37859 30895 37865
rect 30837 37825 30849 37859
rect 30883 37825 30895 37859
rect 30837 37819 30895 37825
rect 30929 37859 30987 37865
rect 30929 37825 30941 37859
rect 30975 37825 30987 37859
rect 30929 37819 30987 37825
rect 31205 37859 31263 37865
rect 31205 37825 31217 37859
rect 31251 37856 31263 37859
rect 31478 37856 31484 37868
rect 31251 37828 31484 37856
rect 31251 37825 31263 37828
rect 31205 37819 31263 37825
rect 28828 37760 29224 37788
rect 28261 37751 28319 37757
rect 27890 37720 27896 37732
rect 27448 37692 27896 37720
rect 24820 37680 24826 37692
rect 22554 37652 22560 37664
rect 18984 37624 22560 37652
rect 22554 37612 22560 37624
rect 22612 37612 22618 37664
rect 26970 37612 26976 37664
rect 27028 37612 27034 37664
rect 27264 37652 27292 37692
rect 27890 37680 27896 37692
rect 27948 37720 27954 37732
rect 28445 37723 28503 37729
rect 28445 37720 28457 37723
rect 27948 37692 28457 37720
rect 27948 37680 27954 37692
rect 28445 37689 28457 37692
rect 28491 37689 28503 37723
rect 28445 37683 28503 37689
rect 28626 37680 28632 37732
rect 28684 37680 28690 37732
rect 28644 37652 28672 37680
rect 27264 37624 28672 37652
rect 28994 37612 29000 37664
rect 29052 37612 29058 37664
rect 29196 37661 29224 37760
rect 29181 37655 29239 37661
rect 29181 37621 29193 37655
rect 29227 37652 29239 37655
rect 29454 37652 29460 37664
rect 29227 37624 29460 37652
rect 29227 37621 29239 37624
rect 29181 37615 29239 37621
rect 29454 37612 29460 37624
rect 29512 37612 29518 37664
rect 30760 37652 30788 37819
rect 30852 37720 30880 37819
rect 30944 37788 30972 37819
rect 31478 37816 31484 37828
rect 31536 37816 31542 37868
rect 33321 37859 33379 37865
rect 33321 37825 33333 37859
rect 33367 37856 33379 37859
rect 33410 37856 33416 37868
rect 33367 37828 33416 37856
rect 33367 37825 33379 37828
rect 33321 37819 33379 37825
rect 33410 37816 33416 37828
rect 33468 37816 33474 37868
rect 33502 37816 33508 37868
rect 33560 37816 33566 37868
rect 35544 37865 35572 37896
rect 36049 37893 36061 37896
rect 36095 37893 36107 37927
rect 36049 37887 36107 37893
rect 36265 37927 36323 37933
rect 36265 37893 36277 37927
rect 36311 37924 36323 37927
rect 36722 37924 36728 37936
rect 36311 37896 36728 37924
rect 36311 37893 36323 37896
rect 36265 37887 36323 37893
rect 36722 37884 36728 37896
rect 36780 37924 36786 37936
rect 38257 37927 38315 37933
rect 38257 37924 38269 37927
rect 36780 37896 37872 37924
rect 36780 37884 36786 37896
rect 34977 37859 35035 37865
rect 34977 37825 34989 37859
rect 35023 37825 35035 37859
rect 35529 37859 35587 37865
rect 35529 37856 35541 37859
rect 34977 37819 35035 37825
rect 35084 37828 35541 37856
rect 32858 37788 32864 37800
rect 30944 37760 32864 37788
rect 32858 37748 32864 37760
rect 32916 37748 32922 37800
rect 31202 37720 31208 37732
rect 30852 37692 31208 37720
rect 31202 37680 31208 37692
rect 31260 37680 31266 37732
rect 34992 37720 35020 37819
rect 35084 37797 35112 37828
rect 35529 37825 35541 37828
rect 35575 37825 35587 37859
rect 35529 37819 35587 37825
rect 35805 37859 35863 37865
rect 35805 37825 35817 37859
rect 35851 37856 35863 37859
rect 36357 37859 36415 37865
rect 36357 37856 36369 37859
rect 35851 37828 36369 37856
rect 35851 37825 35863 37828
rect 35805 37819 35863 37825
rect 36357 37825 36369 37828
rect 36403 37825 36415 37859
rect 36357 37819 36415 37825
rect 36814 37816 36820 37868
rect 36872 37856 36878 37868
rect 37844 37865 37872 37896
rect 38028 37896 38269 37924
rect 37001 37859 37059 37865
rect 37001 37856 37013 37859
rect 36872 37828 37013 37856
rect 36872 37816 36878 37828
rect 37001 37825 37013 37828
rect 37047 37856 37059 37859
rect 37461 37859 37519 37865
rect 37461 37856 37473 37859
rect 37047 37828 37473 37856
rect 37047 37825 37059 37828
rect 37001 37819 37059 37825
rect 37461 37825 37473 37828
rect 37507 37825 37519 37859
rect 37461 37819 37519 37825
rect 37829 37859 37887 37865
rect 37829 37825 37841 37859
rect 37875 37825 37887 37859
rect 37829 37819 37887 37825
rect 35069 37791 35127 37797
rect 35069 37757 35081 37791
rect 35115 37757 35127 37791
rect 35069 37751 35127 37757
rect 35250 37748 35256 37800
rect 35308 37788 35314 37800
rect 35345 37791 35403 37797
rect 35345 37788 35357 37791
rect 35308 37760 35357 37788
rect 35308 37748 35314 37760
rect 35345 37757 35357 37760
rect 35391 37757 35403 37791
rect 35894 37788 35900 37800
rect 35345 37751 35403 37757
rect 35866 37748 35900 37788
rect 35952 37748 35958 37800
rect 35866 37720 35894 37748
rect 34992 37692 35894 37720
rect 32950 37652 32956 37664
rect 30760 37624 32956 37652
rect 32950 37612 32956 37624
rect 33008 37612 33014 37664
rect 35802 37612 35808 37664
rect 35860 37612 35866 37664
rect 35897 37655 35955 37661
rect 35897 37621 35909 37655
rect 35943 37652 35955 37655
rect 35986 37652 35992 37664
rect 35943 37624 35992 37652
rect 35943 37621 35955 37624
rect 35897 37615 35955 37621
rect 35986 37612 35992 37624
rect 36044 37612 36050 37664
rect 36081 37655 36139 37661
rect 36081 37621 36093 37655
rect 36127 37652 36139 37655
rect 36832 37652 36860 37816
rect 38028 37800 38056 37896
rect 38257 37893 38269 37896
rect 38303 37893 38315 37927
rect 38257 37887 38315 37893
rect 38473 37927 38531 37933
rect 38473 37893 38485 37927
rect 38519 37893 38531 37927
rect 38473 37887 38531 37893
rect 37274 37748 37280 37800
rect 37332 37788 37338 37800
rect 37369 37791 37427 37797
rect 37369 37788 37381 37791
rect 37332 37760 37381 37788
rect 37332 37748 37338 37760
rect 37369 37757 37381 37760
rect 37415 37757 37427 37791
rect 37369 37751 37427 37757
rect 37384 37720 37412 37751
rect 38010 37748 38016 37800
rect 38068 37748 38074 37800
rect 38488 37720 38516 37887
rect 38565 37859 38623 37865
rect 38565 37825 38577 37859
rect 38611 37856 38623 37859
rect 38672 37856 38700 37952
rect 38611 37828 38700 37856
rect 38611 37825 38623 37828
rect 38565 37819 38623 37825
rect 40218 37816 40224 37868
rect 40276 37816 40282 37868
rect 40310 37816 40316 37868
rect 40368 37816 40374 37868
rect 42996 37856 43024 37952
rect 43533 37859 43591 37865
rect 43533 37856 43545 37859
rect 42996 37828 43545 37856
rect 43533 37825 43545 37828
rect 43579 37825 43591 37859
rect 43533 37819 43591 37825
rect 38841 37791 38899 37797
rect 38841 37757 38853 37791
rect 38887 37788 38899 37791
rect 39482 37788 39488 37800
rect 38887 37760 39488 37788
rect 38887 37757 38899 37760
rect 38841 37751 38899 37757
rect 39482 37748 39488 37760
rect 39540 37748 39546 37800
rect 39942 37748 39948 37800
rect 40000 37748 40006 37800
rect 40129 37791 40187 37797
rect 40129 37757 40141 37791
rect 40175 37788 40187 37791
rect 40328 37788 40356 37816
rect 40175 37760 40356 37788
rect 40175 37757 40187 37760
rect 40129 37751 40187 37757
rect 43162 37748 43168 37800
rect 43220 37748 43226 37800
rect 37384 37692 38332 37720
rect 38488 37692 38884 37720
rect 36127 37624 36860 37652
rect 36127 37621 36139 37624
rect 36081 37615 36139 37621
rect 37826 37612 37832 37664
rect 37884 37612 37890 37664
rect 38105 37655 38163 37661
rect 38105 37621 38117 37655
rect 38151 37652 38163 37655
rect 38194 37652 38200 37664
rect 38151 37624 38200 37652
rect 38151 37621 38163 37624
rect 38105 37615 38163 37621
rect 38194 37612 38200 37624
rect 38252 37612 38258 37664
rect 38304 37661 38332 37692
rect 38856 37664 38884 37692
rect 38289 37655 38347 37661
rect 38289 37621 38301 37655
rect 38335 37621 38347 37655
rect 38289 37615 38347 37621
rect 38654 37612 38660 37664
rect 38712 37612 38718 37664
rect 38838 37612 38844 37664
rect 38896 37612 38902 37664
rect 44177 37655 44235 37661
rect 44177 37621 44189 37655
rect 44223 37652 44235 37655
rect 44223 37624 44680 37652
rect 44223 37621 44235 37624
rect 44177 37615 44235 37621
rect 1104 37562 44620 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 44620 37562
rect 1104 37488 44620 37510
rect 6914 37408 6920 37460
rect 6972 37448 6978 37460
rect 7101 37451 7159 37457
rect 7101 37448 7113 37451
rect 6972 37420 7113 37448
rect 6972 37408 6978 37420
rect 7101 37417 7113 37420
rect 7147 37417 7159 37451
rect 7101 37411 7159 37417
rect 8938 37408 8944 37460
rect 8996 37408 9002 37460
rect 16669 37451 16727 37457
rect 16669 37417 16681 37451
rect 16715 37448 16727 37451
rect 17034 37448 17040 37460
rect 16715 37420 17040 37448
rect 16715 37417 16727 37420
rect 16669 37411 16727 37417
rect 17034 37408 17040 37420
rect 17092 37408 17098 37460
rect 20714 37408 20720 37460
rect 20772 37408 20778 37460
rect 22462 37448 22468 37460
rect 22066 37420 22468 37448
rect 8202 37272 8208 37324
rect 8260 37272 8266 37324
rect 8956 37321 8984 37408
rect 9214 37380 9220 37392
rect 9140 37352 9220 37380
rect 8941 37315 8999 37321
rect 8941 37281 8953 37315
rect 8987 37281 8999 37315
rect 8941 37275 8999 37281
rect 934 37204 940 37256
rect 992 37244 998 37256
rect 1397 37247 1455 37253
rect 1397 37244 1409 37247
rect 992 37216 1409 37244
rect 992 37204 998 37216
rect 1397 37213 1409 37216
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 5534 37244 5540 37256
rect 1820 37216 5540 37244
rect 1820 37204 1826 37216
rect 5534 37204 5540 37216
rect 5592 37204 5598 37256
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37244 7343 37247
rect 8021 37247 8079 37253
rect 7331 37216 7696 37244
rect 7331 37213 7343 37216
rect 7285 37207 7343 37213
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37108 1639 37111
rect 2130 37108 2136 37120
rect 1627 37080 2136 37108
rect 1627 37077 1639 37080
rect 1581 37071 1639 37077
rect 2130 37068 2136 37080
rect 2188 37068 2194 37120
rect 7668 37117 7696 37216
rect 8021 37213 8033 37247
rect 8067 37244 8079 37247
rect 8386 37244 8392 37256
rect 8067 37216 8392 37244
rect 8067 37213 8079 37216
rect 8021 37207 8079 37213
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 9140 37253 9168 37352
rect 9214 37340 9220 37352
rect 9272 37380 9278 37392
rect 11054 37380 11060 37392
rect 9272 37352 11060 37380
rect 9272 37340 9278 37352
rect 11054 37340 11060 37352
rect 11112 37380 11118 37392
rect 11112 37352 16436 37380
rect 11112 37340 11118 37352
rect 10870 37272 10876 37324
rect 10928 37312 10934 37324
rect 11149 37315 11207 37321
rect 11149 37312 11161 37315
rect 10928 37284 11161 37312
rect 10928 37272 10934 37284
rect 11149 37281 11161 37284
rect 11195 37281 11207 37315
rect 11149 37275 11207 37281
rect 11333 37315 11391 37321
rect 11333 37281 11345 37315
rect 11379 37312 11391 37315
rect 11422 37312 11428 37324
rect 11379 37284 11428 37312
rect 11379 37281 11391 37284
rect 11333 37275 11391 37281
rect 11422 37272 11428 37284
rect 11480 37272 11486 37324
rect 12621 37315 12679 37321
rect 12621 37281 12633 37315
rect 12667 37312 12679 37315
rect 12986 37312 12992 37324
rect 12667 37284 12992 37312
rect 12667 37281 12679 37284
rect 12621 37275 12679 37281
rect 12986 37272 12992 37284
rect 13044 37272 13050 37324
rect 14645 37315 14703 37321
rect 14645 37281 14657 37315
rect 14691 37312 14703 37315
rect 14691 37284 15700 37312
rect 14691 37281 14703 37284
rect 14645 37275 14703 37281
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 12250 37204 12256 37256
rect 12308 37244 12314 37256
rect 13265 37247 13323 37253
rect 13265 37244 13277 37247
rect 12308 37216 13277 37244
rect 12308 37204 12314 37216
rect 13265 37213 13277 37216
rect 13311 37213 13323 37247
rect 13265 37207 13323 37213
rect 13354 37204 13360 37256
rect 13412 37244 13418 37256
rect 13909 37247 13967 37253
rect 13909 37244 13921 37247
rect 13412 37216 13921 37244
rect 13412 37204 13418 37216
rect 13909 37213 13921 37216
rect 13955 37213 13967 37247
rect 15672 37244 15700 37284
rect 16022 37272 16028 37324
rect 16080 37312 16086 37324
rect 16301 37315 16359 37321
rect 16301 37312 16313 37315
rect 16080 37284 16313 37312
rect 16080 37272 16086 37284
rect 16301 37281 16313 37284
rect 16347 37281 16359 37315
rect 16301 37275 16359 37281
rect 16408 37244 16436 37352
rect 16482 37340 16488 37392
rect 16540 37340 16546 37392
rect 16500 37312 16528 37340
rect 18506 37312 18512 37324
rect 16500 37284 18512 37312
rect 16485 37247 16543 37253
rect 16485 37244 16497 37247
rect 15672 37216 16068 37244
rect 16408 37216 16497 37244
rect 13909 37207 13967 37213
rect 16040 37188 16068 37216
rect 16485 37213 16497 37216
rect 16531 37244 16543 37247
rect 16850 37244 16856 37256
rect 16531 37216 16856 37244
rect 16531 37213 16543 37216
rect 16485 37207 16543 37213
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 16942 37204 16948 37256
rect 17000 37244 17006 37256
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 17000 37216 17049 37244
rect 17000 37204 17006 37216
rect 17037 37213 17049 37216
rect 17083 37213 17095 37247
rect 18432 37230 18460 37284
rect 18506 37272 18512 37284
rect 18564 37272 18570 37324
rect 22066 37312 22094 37420
rect 22462 37408 22468 37420
rect 22520 37448 22526 37460
rect 25225 37451 25283 37457
rect 25225 37448 25237 37451
rect 22520 37420 25237 37448
rect 22520 37408 22526 37420
rect 25225 37417 25237 37420
rect 25271 37417 25283 37451
rect 25225 37411 25283 37417
rect 27798 37408 27804 37460
rect 27856 37408 27862 37460
rect 36814 37408 36820 37460
rect 36872 37408 36878 37460
rect 39482 37408 39488 37460
rect 39540 37448 39546 37460
rect 40497 37451 40555 37457
rect 40497 37448 40509 37451
rect 39540 37420 40509 37448
rect 39540 37408 39546 37420
rect 40497 37417 40509 37420
rect 40543 37448 40555 37451
rect 40543 37420 42104 37448
rect 40543 37417 40555 37420
rect 40497 37411 40555 37417
rect 28626 37340 28632 37392
rect 28684 37380 28690 37392
rect 30006 37380 30012 37392
rect 28684 37352 30012 37380
rect 28684 37340 28690 37352
rect 30006 37340 30012 37352
rect 30064 37340 30070 37392
rect 41049 37383 41107 37389
rect 41049 37380 41061 37383
rect 40144 37352 41061 37380
rect 21652 37284 22094 37312
rect 17037 37207 17095 37213
rect 19150 37204 19156 37256
rect 19208 37244 19214 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 19208 37216 19257 37244
rect 19208 37204 19214 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 9309 37179 9367 37185
rect 9309 37145 9321 37179
rect 9355 37176 9367 37179
rect 12894 37176 12900 37188
rect 9355 37148 12900 37176
rect 9355 37145 9367 37148
rect 9309 37139 9367 37145
rect 12894 37136 12900 37148
rect 12952 37136 12958 37188
rect 14829 37179 14887 37185
rect 14829 37145 14841 37179
rect 14875 37176 14887 37179
rect 15473 37179 15531 37185
rect 15473 37176 15485 37179
rect 14875 37148 15485 37176
rect 14875 37145 14887 37148
rect 14829 37139 14887 37145
rect 15473 37145 15485 37148
rect 15519 37145 15531 37179
rect 15473 37139 15531 37145
rect 16022 37136 16028 37188
rect 16080 37136 16086 37188
rect 17310 37136 17316 37188
rect 17368 37136 17374 37188
rect 19058 37136 19064 37188
rect 19116 37176 19122 37188
rect 21652 37176 21680 37284
rect 25406 37272 25412 37324
rect 25464 37312 25470 37324
rect 26053 37315 26111 37321
rect 26053 37312 26065 37315
rect 25464 37284 26065 37312
rect 25464 37272 25470 37284
rect 26053 37281 26065 37284
rect 26099 37281 26111 37315
rect 26053 37275 26111 37281
rect 26329 37315 26387 37321
rect 26329 37281 26341 37315
rect 26375 37312 26387 37315
rect 26970 37312 26976 37324
rect 26375 37284 26976 37312
rect 26375 37281 26387 37284
rect 26329 37275 26387 37281
rect 26970 37272 26976 37284
rect 27028 37272 27034 37324
rect 27522 37272 27528 37324
rect 27580 37312 27586 37324
rect 32766 37312 32772 37324
rect 27580 37284 32772 37312
rect 27580 37272 27586 37284
rect 32766 37272 32772 37284
rect 32824 37272 32830 37324
rect 34790 37272 34796 37324
rect 34848 37312 34854 37324
rect 35069 37315 35127 37321
rect 35069 37312 35081 37315
rect 34848 37284 35081 37312
rect 34848 37272 34854 37284
rect 35069 37281 35081 37284
rect 35115 37281 35127 37315
rect 35069 37275 35127 37281
rect 35986 37272 35992 37324
rect 36044 37312 36050 37324
rect 36044 37284 37228 37312
rect 36044 37272 36050 37284
rect 21726 37204 21732 37256
rect 21784 37244 21790 37256
rect 22465 37247 22523 37253
rect 22465 37244 22477 37247
rect 21784 37216 22477 37244
rect 21784 37204 21790 37216
rect 22465 37213 22477 37216
rect 22511 37213 22523 37247
rect 22465 37207 22523 37213
rect 23842 37204 23848 37256
rect 23900 37204 23906 37256
rect 24394 37204 24400 37256
rect 24452 37204 24458 37256
rect 25314 37204 25320 37256
rect 25372 37244 25378 37256
rect 25501 37247 25559 37253
rect 25501 37244 25513 37247
rect 25372 37216 25513 37244
rect 25372 37204 25378 37216
rect 25501 37213 25513 37216
rect 25547 37213 25559 37247
rect 25501 37207 25559 37213
rect 19116 37148 21680 37176
rect 23109 37179 23167 37185
rect 19116 37136 19122 37148
rect 23109 37145 23121 37179
rect 23155 37176 23167 37179
rect 25516 37176 25544 37207
rect 25682 37204 25688 37256
rect 25740 37204 25746 37256
rect 25869 37247 25927 37253
rect 25869 37213 25881 37247
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 33229 37247 33287 37253
rect 33229 37213 33241 37247
rect 33275 37244 33287 37247
rect 33502 37244 33508 37256
rect 33275 37216 33508 37244
rect 33275 37213 33287 37216
rect 33229 37207 33287 37213
rect 25777 37179 25835 37185
rect 25777 37176 25789 37179
rect 23155 37148 23980 37176
rect 25516 37148 25789 37176
rect 23155 37145 23167 37148
rect 23109 37139 23167 37145
rect 23952 37120 23980 37148
rect 25777 37145 25789 37148
rect 25823 37145 25835 37179
rect 25777 37139 25835 37145
rect 7653 37111 7711 37117
rect 7653 37077 7665 37111
rect 7699 37077 7711 37111
rect 7653 37071 7711 37077
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8113 37111 8171 37117
rect 8113 37108 8125 37111
rect 7800 37080 8125 37108
rect 7800 37068 7806 37080
rect 8113 37077 8125 37080
rect 8159 37077 8171 37111
rect 8113 37071 8171 37077
rect 10686 37068 10692 37120
rect 10744 37068 10750 37120
rect 11054 37068 11060 37120
rect 11112 37068 11118 37120
rect 13173 37111 13231 37117
rect 13173 37077 13185 37111
rect 13219 37108 13231 37111
rect 13446 37108 13452 37120
rect 13219 37080 13452 37108
rect 13219 37077 13231 37080
rect 13173 37071 13231 37077
rect 13446 37068 13452 37080
rect 13504 37068 13510 37120
rect 13630 37068 13636 37120
rect 13688 37108 13694 37120
rect 14737 37111 14795 37117
rect 14737 37108 14749 37111
rect 13688 37080 14749 37108
rect 13688 37068 13694 37080
rect 14737 37077 14749 37080
rect 14783 37077 14795 37111
rect 14737 37071 14795 37077
rect 15194 37068 15200 37120
rect 15252 37068 15258 37120
rect 18782 37068 18788 37120
rect 18840 37068 18846 37120
rect 18966 37068 18972 37120
rect 19024 37108 19030 37120
rect 23201 37111 23259 37117
rect 23201 37108 23213 37111
rect 19024 37080 23213 37108
rect 19024 37068 19030 37080
rect 23201 37077 23213 37080
rect 23247 37108 23259 37111
rect 23750 37108 23756 37120
rect 23247 37080 23756 37108
rect 23247 37077 23259 37080
rect 23201 37071 23259 37077
rect 23750 37068 23756 37080
rect 23808 37068 23814 37120
rect 23934 37068 23940 37120
rect 23992 37068 23998 37120
rect 25038 37068 25044 37120
rect 25096 37068 25102 37120
rect 25884 37108 25912 37207
rect 33502 37204 33508 37216
rect 33560 37244 33566 37256
rect 36906 37244 36912 37256
rect 33560 37216 34100 37244
rect 36478 37216 36912 37244
rect 33560 37204 33566 37216
rect 34072 37188 34100 37216
rect 36906 37204 36912 37216
rect 36964 37204 36970 37256
rect 37200 37244 37228 37284
rect 37826 37272 37832 37324
rect 37884 37312 37890 37324
rect 37884 37284 38884 37312
rect 37884 37272 37890 37284
rect 38856 37256 38884 37284
rect 38010 37244 38016 37256
rect 37200 37216 38016 37244
rect 38010 37204 38016 37216
rect 38068 37204 38074 37256
rect 38197 37247 38255 37253
rect 38197 37213 38209 37247
rect 38243 37244 38255 37247
rect 38654 37244 38660 37256
rect 38243 37216 38660 37244
rect 38243 37213 38255 37216
rect 38197 37207 38255 37213
rect 38654 37204 38660 37216
rect 38712 37204 38718 37256
rect 38838 37204 38844 37256
rect 38896 37204 38902 37256
rect 40034 37204 40040 37256
rect 40092 37244 40098 37256
rect 40144 37253 40172 37352
rect 41049 37349 41061 37352
rect 41095 37349 41107 37383
rect 41049 37343 41107 37349
rect 41230 37312 41236 37324
rect 40696 37284 41236 37312
rect 40129 37247 40187 37253
rect 40129 37244 40141 37247
rect 40092 37216 40141 37244
rect 40092 37204 40098 37216
rect 40129 37213 40141 37216
rect 40175 37213 40187 37247
rect 40129 37207 40187 37213
rect 40497 37247 40555 37253
rect 40497 37213 40509 37247
rect 40543 37244 40555 37247
rect 40696 37244 40724 37284
rect 41230 37272 41236 37284
rect 41288 37272 41294 37324
rect 40543 37216 40724 37244
rect 40773 37247 40831 37253
rect 40543 37213 40555 37216
rect 40497 37207 40555 37213
rect 40773 37213 40785 37247
rect 40819 37213 40831 37247
rect 40773 37207 40831 37213
rect 40957 37247 41015 37253
rect 40957 37213 40969 37247
rect 41003 37244 41015 37247
rect 41003 37216 41460 37244
rect 41003 37213 41015 37216
rect 40957 37207 41015 37213
rect 26786 37136 26792 37188
rect 26844 37136 26850 37188
rect 33413 37179 33471 37185
rect 33413 37145 33425 37179
rect 33459 37176 33471 37179
rect 33870 37176 33876 37188
rect 33459 37148 33876 37176
rect 33459 37145 33471 37148
rect 33413 37139 33471 37145
rect 33870 37136 33876 37148
rect 33928 37136 33934 37188
rect 34054 37136 34060 37188
rect 34112 37136 34118 37188
rect 35342 37136 35348 37188
rect 35400 37136 35406 37188
rect 40788 37176 40816 37207
rect 41325 37179 41383 37185
rect 41325 37176 41337 37179
rect 40788 37148 40908 37176
rect 27614 37108 27620 37120
rect 25884 37080 27620 37108
rect 27614 37068 27620 37080
rect 27672 37068 27678 37120
rect 33045 37111 33103 37117
rect 33045 37077 33057 37111
rect 33091 37108 33103 37111
rect 33318 37108 33324 37120
rect 33091 37080 33324 37108
rect 33091 37077 33103 37080
rect 33045 37071 33103 37077
rect 33318 37068 33324 37080
rect 33376 37068 33382 37120
rect 40880 37108 40908 37148
rect 41156 37148 41337 37176
rect 41156 37120 41184 37148
rect 41325 37145 41337 37148
rect 41371 37145 41383 37179
rect 41325 37139 41383 37145
rect 41432 37120 41460 37216
rect 42076 37185 42104 37420
rect 42242 37408 42248 37460
rect 42300 37408 42306 37460
rect 43993 37315 44051 37321
rect 43993 37281 44005 37315
rect 44039 37312 44051 37315
rect 44652 37312 44680 37624
rect 44039 37284 44680 37312
rect 44039 37281 44051 37284
rect 43993 37275 44051 37281
rect 42978 37244 42984 37256
rect 42918 37216 42984 37244
rect 42978 37204 42984 37216
rect 43036 37204 43042 37256
rect 44266 37204 44272 37256
rect 44324 37204 44330 37256
rect 42061 37179 42119 37185
rect 42061 37145 42073 37179
rect 42107 37145 42119 37179
rect 42061 37139 42119 37145
rect 42277 37179 42335 37185
rect 42277 37145 42289 37179
rect 42323 37176 42335 37179
rect 42610 37176 42616 37188
rect 42323 37148 42616 37176
rect 42323 37145 42335 37148
rect 42277 37139 42335 37145
rect 42610 37136 42616 37148
rect 42668 37136 42674 37188
rect 41138 37108 41144 37120
rect 40880 37080 41144 37108
rect 41138 37068 41144 37080
rect 41196 37068 41202 37120
rect 41230 37068 41236 37120
rect 41288 37068 41294 37120
rect 41414 37068 41420 37120
rect 41472 37068 41478 37120
rect 41598 37068 41604 37120
rect 41656 37068 41662 37120
rect 41782 37068 41788 37120
rect 41840 37108 41846 37120
rect 42429 37111 42487 37117
rect 42429 37108 42441 37111
rect 41840 37080 42441 37108
rect 41840 37068 41846 37080
rect 42429 37077 42441 37080
rect 42475 37077 42487 37111
rect 42429 37071 42487 37077
rect 42521 37111 42579 37117
rect 42521 37077 42533 37111
rect 42567 37108 42579 37111
rect 43162 37108 43168 37120
rect 42567 37080 43168 37108
rect 42567 37077 42579 37080
rect 42521 37071 42579 37077
rect 43162 37068 43168 37080
rect 43220 37068 43226 37120
rect 1104 37018 44620 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 44620 37018
rect 1104 36944 44620 36966
rect 4448 36876 6776 36904
rect 4448 36836 4476 36876
rect 6748 36848 6776 36876
rect 12250 36864 12256 36916
rect 12308 36864 12314 36916
rect 13446 36864 13452 36916
rect 13504 36904 13510 36916
rect 13504 36876 13768 36904
rect 13504 36864 13510 36876
rect 4356 36808 4476 36836
rect 4356 36777 4384 36808
rect 6730 36796 6736 36848
rect 6788 36796 6794 36848
rect 13740 36845 13768 36876
rect 15194 36864 15200 36916
rect 15252 36864 15258 36916
rect 15286 36864 15292 36916
rect 15344 36864 15350 36916
rect 16666 36864 16672 36916
rect 16724 36864 16730 36916
rect 17310 36864 17316 36916
rect 17368 36864 17374 36916
rect 18782 36864 18788 36916
rect 18840 36864 18846 36916
rect 18874 36864 18880 36916
rect 18932 36904 18938 36916
rect 19429 36907 19487 36913
rect 18932 36876 19196 36904
rect 18932 36864 18938 36876
rect 13725 36839 13783 36845
rect 13725 36805 13737 36839
rect 13771 36805 13783 36839
rect 13725 36799 13783 36805
rect 4341 36771 4399 36777
rect 4341 36737 4353 36771
rect 4387 36737 4399 36771
rect 6917 36771 6975 36777
rect 5750 36740 5856 36768
rect 4341 36731 4399 36737
rect 1762 36660 1768 36712
rect 1820 36660 1826 36712
rect 4614 36660 4620 36712
rect 4672 36660 4678 36712
rect 2130 36592 2136 36644
rect 2188 36592 2194 36644
rect 5828 36576 5856 36740
rect 6917 36737 6929 36771
rect 6963 36768 6975 36771
rect 8202 36768 8208 36780
rect 6963 36740 8208 36768
rect 6963 36737 6975 36740
rect 6917 36731 6975 36737
rect 8202 36728 8208 36740
rect 8260 36728 8266 36780
rect 10962 36728 10968 36780
rect 11020 36768 11026 36780
rect 11020 36740 12204 36768
rect 11020 36728 11026 36740
rect 12176 36712 12204 36740
rect 12618 36728 12624 36780
rect 12676 36728 12682 36780
rect 13998 36728 14004 36780
rect 14056 36728 14062 36780
rect 15212 36768 15240 36864
rect 16022 36796 16028 36848
rect 16080 36796 16086 36848
rect 16684 36836 16712 36864
rect 17126 36836 17132 36848
rect 16684 36808 17132 36836
rect 15473 36771 15531 36777
rect 15473 36768 15485 36771
rect 15212 36740 15485 36768
rect 15473 36737 15485 36740
rect 15519 36737 15531 36771
rect 15473 36731 15531 36737
rect 16393 36771 16451 36777
rect 16393 36737 16405 36771
rect 16439 36768 16451 36771
rect 16666 36768 16672 36780
rect 16439 36740 16672 36768
rect 16439 36737 16451 36740
rect 16393 36731 16451 36737
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 16776 36777 16804 36808
rect 17126 36796 17132 36808
rect 17184 36796 17190 36848
rect 17218 36796 17224 36848
rect 17276 36836 17282 36848
rect 18800 36836 18828 36864
rect 19168 36845 19196 36876
rect 19429 36873 19441 36907
rect 19475 36904 19487 36907
rect 20990 36904 20996 36916
rect 19475 36876 20996 36904
rect 19475 36873 19487 36876
rect 19429 36867 19487 36873
rect 20990 36864 20996 36876
rect 21048 36864 21054 36916
rect 23842 36864 23848 36916
rect 23900 36864 23906 36916
rect 25038 36864 25044 36916
rect 25096 36864 25102 36916
rect 25406 36864 25412 36916
rect 25464 36864 25470 36916
rect 27706 36864 27712 36916
rect 27764 36904 27770 36916
rect 28353 36907 28411 36913
rect 28353 36904 28365 36907
rect 27764 36876 28365 36904
rect 27764 36864 27770 36876
rect 28353 36873 28365 36876
rect 28399 36873 28411 36907
rect 28353 36867 28411 36873
rect 31202 36864 31208 36916
rect 31260 36904 31266 36916
rect 31662 36904 31668 36916
rect 31260 36876 31668 36904
rect 31260 36864 31266 36876
rect 31662 36864 31668 36876
rect 31720 36904 31726 36916
rect 32217 36907 32275 36913
rect 32217 36904 32229 36907
rect 31720 36876 32229 36904
rect 31720 36864 31726 36876
rect 32217 36873 32229 36876
rect 32263 36873 32275 36907
rect 33045 36907 33103 36913
rect 33045 36904 33057 36907
rect 32217 36867 32275 36873
rect 32324 36876 33057 36904
rect 17276 36808 18644 36836
rect 17276 36796 17282 36808
rect 16761 36771 16819 36777
rect 16761 36737 16773 36771
rect 16807 36737 16819 36771
rect 16761 36731 16819 36737
rect 16853 36771 16911 36777
rect 16853 36737 16865 36771
rect 16899 36768 16911 36771
rect 16899 36740 16988 36768
rect 16899 36737 16911 36740
rect 16853 36731 16911 36737
rect 6089 36703 6147 36709
rect 6089 36669 6101 36703
rect 6135 36700 6147 36703
rect 6362 36700 6368 36712
rect 6135 36672 6368 36700
rect 6135 36669 6147 36672
rect 6089 36663 6147 36669
rect 6362 36660 6368 36672
rect 6420 36700 6426 36712
rect 8294 36700 8300 36712
rect 6420 36672 8300 36700
rect 6420 36660 6426 36672
rect 8294 36660 8300 36672
rect 8352 36660 8358 36712
rect 8665 36703 8723 36709
rect 8665 36669 8677 36703
rect 8711 36700 8723 36703
rect 9398 36700 9404 36712
rect 8711 36672 9404 36700
rect 8711 36669 8723 36672
rect 8665 36663 8723 36669
rect 9398 36660 9404 36672
rect 9456 36700 9462 36712
rect 9585 36703 9643 36709
rect 9585 36700 9597 36703
rect 9456 36672 9597 36700
rect 9456 36660 9462 36672
rect 9585 36669 9597 36672
rect 9631 36669 9643 36703
rect 9585 36663 9643 36669
rect 9858 36660 9864 36712
rect 9916 36660 9922 36712
rect 12158 36660 12164 36712
rect 12216 36660 12222 36712
rect 16960 36632 16988 36740
rect 17034 36728 17040 36780
rect 17092 36728 17098 36780
rect 17221 36703 17279 36709
rect 17221 36669 17233 36703
rect 17267 36700 17279 36703
rect 17865 36703 17923 36709
rect 17865 36700 17877 36703
rect 17267 36672 17877 36700
rect 17267 36669 17279 36672
rect 17221 36663 17279 36669
rect 17865 36669 17877 36672
rect 17911 36669 17923 36703
rect 18616 36700 18644 36808
rect 18708 36808 18828 36836
rect 19153 36839 19211 36845
rect 18708 36777 18736 36808
rect 19153 36805 19165 36839
rect 19199 36805 19211 36839
rect 22649 36839 22707 36845
rect 19153 36799 19211 36805
rect 19352 36808 22094 36836
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36737 18751 36771
rect 18693 36731 18751 36737
rect 18782 36728 18788 36780
rect 18840 36728 18846 36780
rect 18966 36777 18972 36780
rect 18933 36771 18972 36777
rect 18933 36737 18945 36771
rect 18933 36731 18972 36737
rect 18966 36728 18972 36731
rect 19024 36728 19030 36780
rect 19058 36728 19064 36780
rect 19116 36728 19122 36780
rect 19242 36768 19248 36780
rect 19300 36777 19306 36780
rect 19208 36740 19248 36768
rect 19242 36728 19248 36740
rect 19300 36768 19308 36777
rect 19352 36768 19380 36808
rect 19300 36740 19380 36768
rect 19889 36771 19947 36777
rect 19300 36731 19308 36740
rect 19889 36737 19901 36771
rect 19935 36768 19947 36771
rect 20441 36771 20499 36777
rect 20441 36768 20453 36771
rect 19935 36740 20453 36768
rect 19935 36737 19947 36740
rect 19889 36731 19947 36737
rect 20441 36737 20453 36740
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 21361 36771 21419 36777
rect 21361 36737 21373 36771
rect 21407 36737 21419 36771
rect 21361 36731 21419 36737
rect 19300 36728 19306 36731
rect 19076 36700 19104 36728
rect 18616 36672 19104 36700
rect 17865 36663 17923 36669
rect 19334 36660 19340 36712
rect 19392 36700 19398 36712
rect 19613 36703 19671 36709
rect 19613 36700 19625 36703
rect 19392 36672 19625 36700
rect 19392 36660 19398 36672
rect 19613 36669 19625 36672
rect 19659 36669 19671 36703
rect 19613 36663 19671 36669
rect 19797 36703 19855 36709
rect 19797 36669 19809 36703
rect 19843 36669 19855 36703
rect 19797 36663 19855 36669
rect 18049 36635 18107 36641
rect 18049 36632 18061 36635
rect 10980 36604 12204 36632
rect 16960 36604 18061 36632
rect 2222 36524 2228 36576
rect 2280 36524 2286 36576
rect 5810 36524 5816 36576
rect 5868 36524 5874 36576
rect 8662 36524 8668 36576
rect 8720 36564 8726 36576
rect 10980 36564 11008 36604
rect 8720 36536 11008 36564
rect 8720 36524 8726 36536
rect 11054 36524 11060 36576
rect 11112 36564 11118 36576
rect 11333 36567 11391 36573
rect 11333 36564 11345 36567
rect 11112 36536 11345 36564
rect 11112 36524 11118 36536
rect 11333 36533 11345 36536
rect 11379 36564 11391 36567
rect 12066 36564 12072 36576
rect 11379 36536 12072 36564
rect 11379 36533 11391 36536
rect 11333 36527 11391 36533
rect 12066 36524 12072 36536
rect 12124 36524 12130 36576
rect 12176 36564 12204 36604
rect 18049 36601 18061 36604
rect 18095 36632 18107 36635
rect 19812 36632 19840 36663
rect 20530 36660 20536 36712
rect 20588 36700 20594 36712
rect 20993 36703 21051 36709
rect 20993 36700 21005 36703
rect 20588 36672 21005 36700
rect 20588 36660 20594 36672
rect 20993 36669 21005 36672
rect 21039 36669 21051 36703
rect 20993 36663 21051 36669
rect 18095 36604 19840 36632
rect 20257 36635 20315 36641
rect 18095 36601 18107 36604
rect 18049 36595 18107 36601
rect 20257 36601 20269 36635
rect 20303 36632 20315 36635
rect 21376 36632 21404 36731
rect 20303 36604 21404 36632
rect 22066 36632 22094 36808
rect 22649 36805 22661 36839
rect 22695 36836 22707 36839
rect 23934 36836 23940 36848
rect 22695 36808 23940 36836
rect 22695 36805 22707 36808
rect 22649 36799 22707 36805
rect 23934 36796 23940 36808
rect 23992 36796 23998 36848
rect 25056 36836 25084 36864
rect 25317 36839 25375 36845
rect 25317 36836 25329 36839
rect 25056 36808 25329 36836
rect 25317 36805 25329 36808
rect 25363 36805 25375 36839
rect 25424 36836 25452 36864
rect 25424 36808 25636 36836
rect 25317 36799 25375 36805
rect 22554 36728 22560 36780
rect 22612 36728 22618 36780
rect 25608 36777 25636 36808
rect 25593 36771 25651 36777
rect 22738 36660 22744 36712
rect 22796 36660 22802 36712
rect 23658 36660 23664 36712
rect 23716 36660 23722 36712
rect 24228 36700 24256 36754
rect 25593 36737 25605 36771
rect 25639 36737 25651 36771
rect 25593 36731 25651 36737
rect 25958 36728 25964 36780
rect 26016 36728 26022 36780
rect 27062 36728 27068 36780
rect 27120 36768 27126 36780
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 27120 36740 27169 36768
rect 27120 36728 27126 36740
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27724 36768 27752 36864
rect 28994 36836 29000 36848
rect 28460 36808 29000 36836
rect 27893 36771 27951 36777
rect 27893 36768 27905 36771
rect 27724 36740 27905 36768
rect 27157 36731 27215 36737
rect 27893 36737 27905 36740
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 28166 36728 28172 36780
rect 28224 36728 28230 36780
rect 28460 36777 28488 36808
rect 28994 36796 29000 36808
rect 29052 36796 29058 36848
rect 28445 36771 28503 36777
rect 28445 36737 28457 36771
rect 28491 36737 28503 36771
rect 28445 36731 28503 36737
rect 30190 36728 30196 36780
rect 30248 36768 30254 36780
rect 30285 36771 30343 36777
rect 30285 36768 30297 36771
rect 30248 36740 30297 36768
rect 30248 36728 30254 36740
rect 30285 36737 30297 36740
rect 30331 36737 30343 36771
rect 30285 36731 30343 36737
rect 25222 36700 25228 36712
rect 24228 36672 25228 36700
rect 25222 36660 25228 36672
rect 25280 36660 25286 36712
rect 27801 36703 27859 36709
rect 27801 36669 27813 36703
rect 27847 36700 27859 36703
rect 28077 36703 28135 36709
rect 28077 36700 28089 36703
rect 27847 36672 28089 36700
rect 27847 36669 27859 36672
rect 27801 36663 27859 36669
rect 28077 36669 28089 36672
rect 28123 36669 28135 36703
rect 32324 36700 32352 36876
rect 33045 36873 33057 36876
rect 33091 36904 33103 36907
rect 33134 36904 33140 36916
rect 33091 36876 33140 36904
rect 33091 36873 33103 36876
rect 33045 36867 33103 36873
rect 33134 36864 33140 36876
rect 33192 36904 33198 36916
rect 33192 36876 33824 36904
rect 33192 36864 33198 36876
rect 33689 36839 33747 36845
rect 33689 36836 33701 36839
rect 32876 36808 33701 36836
rect 32876 36777 32904 36808
rect 33689 36805 33701 36808
rect 33735 36805 33747 36839
rect 33689 36799 33747 36805
rect 32401 36771 32459 36777
rect 32401 36737 32413 36771
rect 32447 36768 32459 36771
rect 32861 36771 32919 36777
rect 32861 36768 32873 36771
rect 32447 36740 32873 36768
rect 32447 36737 32459 36740
rect 32401 36731 32459 36737
rect 32861 36737 32873 36740
rect 32907 36737 32919 36771
rect 32861 36731 32919 36737
rect 32953 36771 33011 36777
rect 32953 36737 32965 36771
rect 32999 36737 33011 36771
rect 32953 36731 33011 36737
rect 33321 36771 33379 36777
rect 33321 36737 33333 36771
rect 33367 36737 33379 36771
rect 33321 36731 33379 36737
rect 32493 36703 32551 36709
rect 32493 36700 32505 36703
rect 32324 36672 32505 36700
rect 28077 36663 28135 36669
rect 32493 36669 32505 36672
rect 32539 36669 32551 36703
rect 32493 36663 32551 36669
rect 32585 36703 32643 36709
rect 32585 36669 32597 36703
rect 32631 36669 32643 36703
rect 32585 36663 32643 36669
rect 26237 36635 26295 36641
rect 22066 36604 24348 36632
rect 20303 36601 20315 36604
rect 20257 36595 20315 36601
rect 16390 36564 16396 36576
rect 12176 36536 16396 36564
rect 16390 36524 16396 36536
rect 16448 36524 16454 36576
rect 21174 36524 21180 36576
rect 21232 36524 21238 36576
rect 22186 36524 22192 36576
rect 22244 36524 22250 36576
rect 23106 36524 23112 36576
rect 23164 36524 23170 36576
rect 24320 36564 24348 36604
rect 26237 36601 26249 36635
rect 26283 36632 26295 36635
rect 26283 36604 27476 36632
rect 26283 36601 26295 36604
rect 26237 36595 26295 36601
rect 27448 36576 27476 36604
rect 24854 36564 24860 36576
rect 24320 36536 24860 36564
rect 24854 36524 24860 36536
rect 24912 36524 24918 36576
rect 26970 36524 26976 36576
rect 27028 36524 27034 36576
rect 27430 36524 27436 36576
rect 27488 36524 27494 36576
rect 27522 36524 27528 36576
rect 27580 36524 27586 36576
rect 27614 36524 27620 36576
rect 27672 36564 27678 36576
rect 27709 36567 27767 36573
rect 27709 36564 27721 36567
rect 27672 36536 27721 36564
rect 27672 36524 27678 36536
rect 27709 36533 27721 36536
rect 27755 36533 27767 36567
rect 27709 36527 27767 36533
rect 30101 36567 30159 36573
rect 30101 36533 30113 36567
rect 30147 36564 30159 36567
rect 31110 36564 31116 36576
rect 30147 36536 31116 36564
rect 30147 36533 30159 36536
rect 30101 36527 30159 36533
rect 31110 36524 31116 36536
rect 31168 36524 31174 36576
rect 32600 36564 32628 36663
rect 32674 36660 32680 36712
rect 32732 36700 32738 36712
rect 32968 36700 32996 36731
rect 32732 36672 32996 36700
rect 32732 36660 32738 36672
rect 33226 36660 33232 36712
rect 33284 36660 33290 36712
rect 33336 36644 33364 36731
rect 33410 36728 33416 36780
rect 33468 36768 33474 36780
rect 33796 36777 33824 36876
rect 33870 36864 33876 36916
rect 33928 36864 33934 36916
rect 34054 36864 34060 36916
rect 34112 36864 34118 36916
rect 35342 36864 35348 36916
rect 35400 36904 35406 36916
rect 35897 36907 35955 36913
rect 35897 36904 35909 36907
rect 35400 36876 35909 36904
rect 35400 36864 35406 36876
rect 35897 36873 35909 36876
rect 35943 36873 35955 36907
rect 41598 36904 41604 36916
rect 35897 36867 35955 36873
rect 40696 36876 41604 36904
rect 35621 36839 35679 36845
rect 35621 36805 35633 36839
rect 35667 36836 35679 36839
rect 35802 36836 35808 36848
rect 35667 36808 35808 36836
rect 35667 36805 35679 36808
rect 35621 36799 35679 36805
rect 35802 36796 35808 36808
rect 35860 36796 35866 36848
rect 40696 36845 40724 36876
rect 41598 36864 41604 36876
rect 41656 36864 41662 36916
rect 41782 36864 41788 36916
rect 41840 36864 41846 36916
rect 41877 36907 41935 36913
rect 41877 36873 41889 36907
rect 41923 36904 41935 36907
rect 42242 36904 42248 36916
rect 41923 36876 42248 36904
rect 41923 36873 41935 36876
rect 41877 36867 41935 36873
rect 42242 36864 42248 36876
rect 42300 36864 42306 36916
rect 44266 36904 44272 36916
rect 42444 36876 44272 36904
rect 38105 36839 38163 36845
rect 38105 36836 38117 36839
rect 37752 36808 38117 36836
rect 33505 36771 33563 36777
rect 33505 36768 33517 36771
rect 33468 36740 33517 36768
rect 33468 36728 33474 36740
rect 33505 36737 33517 36740
rect 33551 36737 33563 36771
rect 33505 36731 33563 36737
rect 33781 36771 33839 36777
rect 33781 36737 33793 36771
rect 33827 36737 33839 36771
rect 33781 36731 33839 36737
rect 33520 36700 33548 36731
rect 33870 36728 33876 36780
rect 33928 36728 33934 36780
rect 33962 36728 33968 36780
rect 34020 36728 34026 36780
rect 34057 36771 34115 36777
rect 34057 36737 34069 36771
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 33888 36700 33916 36728
rect 34072 36700 34100 36731
rect 34238 36728 34244 36780
rect 34296 36728 34302 36780
rect 37752 36777 37780 36808
rect 38105 36805 38117 36808
rect 38151 36805 38163 36839
rect 38105 36799 38163 36805
rect 40681 36839 40739 36845
rect 40681 36805 40693 36839
rect 40727 36805 40739 36839
rect 41800 36836 41828 36864
rect 40681 36799 40739 36805
rect 41616 36808 41828 36836
rect 35897 36771 35955 36777
rect 35897 36737 35909 36771
rect 35943 36737 35955 36771
rect 35897 36731 35955 36737
rect 37737 36771 37795 36777
rect 37737 36737 37749 36771
rect 37783 36737 37795 36771
rect 37737 36731 37795 36737
rect 37921 36771 37979 36777
rect 37921 36737 37933 36771
rect 37967 36737 37979 36771
rect 37921 36731 37979 36737
rect 33520 36672 33916 36700
rect 33980 36672 34100 36700
rect 32950 36592 32956 36644
rect 33008 36632 33014 36644
rect 33137 36635 33195 36641
rect 33137 36632 33149 36635
rect 33008 36604 33149 36632
rect 33008 36592 33014 36604
rect 33137 36601 33149 36604
rect 33183 36601 33195 36635
rect 33137 36595 33195 36601
rect 33318 36592 33324 36644
rect 33376 36592 33382 36644
rect 33226 36564 33232 36576
rect 32600 36536 33232 36564
rect 33226 36524 33232 36536
rect 33284 36564 33290 36576
rect 33980 36564 34008 36672
rect 35805 36635 35863 36641
rect 35805 36601 35817 36635
rect 35851 36601 35863 36635
rect 35912 36632 35940 36731
rect 37936 36700 37964 36731
rect 38010 36728 38016 36780
rect 38068 36728 38074 36780
rect 38197 36771 38255 36777
rect 38197 36737 38209 36771
rect 38243 36768 38255 36771
rect 38565 36771 38623 36777
rect 38565 36768 38577 36771
rect 38243 36740 38577 36768
rect 38243 36737 38255 36740
rect 38197 36731 38255 36737
rect 38565 36737 38577 36740
rect 38611 36737 38623 36771
rect 38565 36731 38623 36737
rect 38654 36728 38660 36780
rect 38712 36728 38718 36780
rect 41616 36777 41644 36808
rect 41601 36771 41659 36777
rect 41601 36737 41613 36771
rect 41647 36737 41659 36771
rect 42061 36771 42119 36777
rect 42061 36768 42073 36771
rect 41601 36731 41659 36737
rect 41708 36740 42073 36768
rect 38672 36700 38700 36728
rect 37936 36672 38700 36700
rect 38838 36660 38844 36712
rect 38896 36700 38902 36712
rect 39117 36703 39175 36709
rect 39117 36700 39129 36703
rect 38896 36672 39129 36700
rect 38896 36660 38902 36672
rect 39117 36669 39129 36672
rect 39163 36669 39175 36703
rect 39117 36663 39175 36669
rect 39942 36632 39948 36644
rect 35912 36604 39948 36632
rect 35805 36595 35863 36601
rect 33284 36536 34008 36564
rect 35820 36564 35848 36595
rect 39942 36592 39948 36604
rect 40000 36632 40006 36644
rect 40126 36632 40132 36644
rect 40000 36604 40132 36632
rect 40000 36592 40006 36604
rect 40126 36592 40132 36604
rect 40184 36632 40190 36644
rect 40405 36635 40463 36641
rect 40405 36632 40417 36635
rect 40184 36604 40417 36632
rect 40184 36592 40190 36604
rect 40405 36601 40417 36604
rect 40451 36601 40463 36635
rect 40405 36595 40463 36601
rect 35986 36564 35992 36576
rect 35820 36536 35992 36564
rect 33284 36524 33290 36536
rect 35986 36524 35992 36536
rect 36044 36524 36050 36576
rect 37734 36524 37740 36576
rect 37792 36524 37798 36576
rect 41708 36564 41736 36740
rect 42061 36737 42073 36740
rect 42107 36737 42119 36771
rect 42061 36731 42119 36737
rect 42242 36728 42248 36780
rect 42300 36728 42306 36780
rect 42444 36777 42472 36876
rect 44266 36864 44272 36876
rect 44324 36864 44330 36916
rect 42978 36796 42984 36848
rect 43036 36836 43042 36848
rect 43036 36808 43194 36836
rect 43036 36796 43042 36808
rect 42429 36771 42487 36777
rect 42429 36737 42441 36771
rect 42475 36737 42487 36771
rect 42429 36731 42487 36737
rect 42705 36703 42763 36709
rect 42705 36700 42717 36703
rect 41800 36672 42717 36700
rect 41800 36641 41828 36672
rect 42705 36669 42717 36672
rect 42751 36669 42763 36703
rect 42705 36663 42763 36669
rect 41785 36635 41843 36641
rect 41785 36601 41797 36635
rect 41831 36601 41843 36635
rect 41785 36595 41843 36601
rect 43070 36564 43076 36576
rect 41708 36536 43076 36564
rect 43070 36524 43076 36536
rect 43128 36564 43134 36576
rect 44177 36567 44235 36573
rect 44177 36564 44189 36567
rect 43128 36536 44189 36564
rect 43128 36524 43134 36536
rect 44177 36533 44189 36536
rect 44223 36533 44235 36567
rect 44177 36527 44235 36533
rect 1104 36474 44620 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 44620 36474
rect 1104 36400 44620 36422
rect 4614 36320 4620 36372
rect 4672 36360 4678 36372
rect 5905 36363 5963 36369
rect 5905 36360 5917 36363
rect 4672 36332 5917 36360
rect 4672 36320 4678 36332
rect 5905 36329 5917 36332
rect 5951 36329 5963 36363
rect 5905 36323 5963 36329
rect 8202 36320 8208 36372
rect 8260 36360 8266 36372
rect 13262 36360 13268 36372
rect 8260 36332 13268 36360
rect 8260 36320 8266 36332
rect 13262 36320 13268 36332
rect 13320 36320 13326 36372
rect 20735 36363 20793 36369
rect 20735 36329 20747 36363
rect 20781 36360 20793 36363
rect 21174 36360 21180 36372
rect 20781 36332 21180 36360
rect 20781 36329 20793 36332
rect 20735 36323 20793 36329
rect 21174 36320 21180 36332
rect 21232 36320 21238 36372
rect 21726 36320 21732 36372
rect 21784 36320 21790 36372
rect 22186 36320 22192 36372
rect 22244 36320 22250 36372
rect 23569 36363 23627 36369
rect 23569 36329 23581 36363
rect 23615 36360 23627 36363
rect 23658 36360 23664 36372
rect 23615 36332 23664 36360
rect 23615 36329 23627 36332
rect 23569 36323 23627 36329
rect 23658 36320 23664 36332
rect 23716 36320 23722 36372
rect 24394 36320 24400 36372
rect 24452 36320 24458 36372
rect 27985 36363 28043 36369
rect 27985 36329 27997 36363
rect 28031 36360 28043 36363
rect 28166 36360 28172 36372
rect 28031 36332 28172 36360
rect 28031 36329 28043 36332
rect 27985 36323 28043 36329
rect 28166 36320 28172 36332
rect 28224 36320 28230 36372
rect 31662 36320 31668 36372
rect 31720 36360 31726 36372
rect 31720 36332 32260 36360
rect 31720 36320 31726 36332
rect 8662 36252 8668 36304
rect 8720 36292 8726 36304
rect 8846 36292 8852 36304
rect 8720 36264 8852 36292
rect 8720 36252 8726 36264
rect 8846 36252 8852 36264
rect 8904 36252 8910 36304
rect 9858 36252 9864 36304
rect 9916 36292 9922 36304
rect 10321 36295 10379 36301
rect 10321 36292 10333 36295
rect 9916 36264 10333 36292
rect 9916 36252 9922 36264
rect 10321 36261 10333 36264
rect 10367 36261 10379 36295
rect 10321 36255 10379 36261
rect 10686 36252 10692 36304
rect 10744 36252 10750 36304
rect 16669 36295 16727 36301
rect 16669 36261 16681 36295
rect 16715 36292 16727 36295
rect 21637 36295 21695 36301
rect 16715 36264 17448 36292
rect 16715 36261 16727 36264
rect 16669 36255 16727 36261
rect 3789 36227 3847 36233
rect 3789 36193 3801 36227
rect 3835 36224 3847 36227
rect 6730 36224 6736 36236
rect 3835 36196 6736 36224
rect 3835 36193 3847 36196
rect 3789 36187 3847 36193
rect 6730 36184 6736 36196
rect 6788 36224 6794 36236
rect 6917 36227 6975 36233
rect 6917 36224 6929 36227
rect 6788 36196 6929 36224
rect 6788 36184 6794 36196
rect 6917 36193 6929 36196
rect 6963 36224 6975 36227
rect 9398 36224 9404 36236
rect 6963 36196 9404 36224
rect 6963 36193 6975 36196
rect 6917 36187 6975 36193
rect 9398 36184 9404 36196
rect 9456 36184 9462 36236
rect 6086 36116 6092 36168
rect 6144 36116 6150 36168
rect 8478 36156 8484 36168
rect 8326 36142 8484 36156
rect 8312 36128 8484 36142
rect 4062 36048 4068 36100
rect 4120 36048 4126 36100
rect 5810 36088 5816 36100
rect 5290 36060 5816 36088
rect 5810 36048 5816 36060
rect 5868 36088 5874 36100
rect 5868 36060 5948 36088
rect 5868 36048 5874 36060
rect 5537 36023 5595 36029
rect 5537 35989 5549 36023
rect 5583 36020 5595 36023
rect 5718 36020 5724 36032
rect 5583 35992 5724 36020
rect 5583 35989 5595 35992
rect 5537 35983 5595 35989
rect 5718 35980 5724 35992
rect 5776 35980 5782 36032
rect 5920 36020 5948 36060
rect 7190 36048 7196 36100
rect 7248 36048 7254 36100
rect 7374 36020 7380 36032
rect 5920 35992 7380 36020
rect 7374 35980 7380 35992
rect 7432 36020 7438 36032
rect 8312 36020 8340 36128
rect 8478 36116 8484 36128
rect 8536 36116 8542 36168
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36156 10563 36159
rect 10704 36156 10732 36252
rect 11793 36227 11851 36233
rect 11793 36193 11805 36227
rect 11839 36224 11851 36227
rect 13998 36224 14004 36236
rect 11839 36196 14004 36224
rect 11839 36193 11851 36196
rect 11793 36187 11851 36193
rect 13998 36184 14004 36196
rect 14056 36184 14062 36236
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 16942 36224 16948 36236
rect 14967 36196 16948 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 16942 36184 16948 36196
rect 17000 36184 17006 36236
rect 17420 36233 17448 36264
rect 21637 36261 21649 36295
rect 21683 36292 21695 36295
rect 22094 36292 22100 36304
rect 21683 36264 22100 36292
rect 21683 36261 21695 36264
rect 21637 36255 21695 36261
rect 22094 36252 22100 36264
rect 22152 36252 22158 36304
rect 17405 36227 17463 36233
rect 17405 36193 17417 36227
rect 17451 36224 17463 36227
rect 17494 36224 17500 36236
rect 17451 36196 17500 36224
rect 17451 36193 17463 36196
rect 17405 36187 17463 36193
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 20714 36184 20720 36236
rect 20772 36224 20778 36236
rect 20993 36227 21051 36233
rect 20993 36224 21005 36227
rect 20772 36196 21005 36224
rect 20772 36184 20778 36196
rect 20993 36193 21005 36196
rect 21039 36193 21051 36227
rect 22204 36224 22232 36320
rect 24854 36252 24860 36304
rect 24912 36292 24918 36304
rect 25317 36295 25375 36301
rect 25317 36292 25329 36295
rect 24912 36264 25329 36292
rect 24912 36252 24918 36264
rect 25317 36261 25329 36264
rect 25363 36261 25375 36295
rect 25317 36255 25375 36261
rect 20993 36187 21051 36193
rect 21468 36196 22232 36224
rect 10551 36128 10732 36156
rect 14645 36159 14703 36165
rect 10551 36125 10563 36128
rect 10505 36119 10563 36125
rect 14645 36125 14657 36159
rect 14691 36125 14703 36159
rect 16482 36156 16488 36168
rect 16330 36128 16488 36156
rect 14645 36119 14703 36125
rect 12069 36091 12127 36097
rect 12069 36057 12081 36091
rect 12115 36057 12127 36091
rect 12069 36051 12127 36057
rect 7432 35992 8340 36020
rect 12084 36020 12112 36051
rect 12158 36048 12164 36100
rect 12216 36088 12222 36100
rect 14660 36088 14688 36119
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 21468 36165 21496 36196
rect 23106 36184 23112 36236
rect 23164 36224 23170 36236
rect 23201 36227 23259 36233
rect 23201 36224 23213 36227
rect 23164 36196 23213 36224
rect 23164 36184 23170 36196
rect 23201 36193 23213 36196
rect 23247 36193 23259 36227
rect 23201 36187 23259 36193
rect 23477 36227 23535 36233
rect 23477 36193 23489 36227
rect 23523 36224 23535 36227
rect 23566 36224 23572 36236
rect 23523 36196 23572 36224
rect 23523 36193 23535 36196
rect 23477 36187 23535 36193
rect 23566 36184 23572 36196
rect 23624 36224 23630 36236
rect 25406 36224 25412 36236
rect 23624 36196 25412 36224
rect 23624 36184 23630 36196
rect 25406 36184 25412 36196
rect 25464 36224 25470 36236
rect 26237 36227 26295 36233
rect 26237 36224 26249 36227
rect 25464 36196 26249 36224
rect 25464 36184 25470 36196
rect 26237 36193 26249 36196
rect 26283 36193 26295 36227
rect 26237 36187 26295 36193
rect 26513 36227 26571 36233
rect 26513 36193 26525 36227
rect 26559 36224 26571 36227
rect 26970 36224 26976 36236
rect 26559 36196 26976 36224
rect 26559 36193 26571 36196
rect 26513 36187 26571 36193
rect 26970 36184 26976 36196
rect 27028 36184 27034 36236
rect 21453 36159 21511 36165
rect 21453 36125 21465 36159
rect 21499 36125 21511 36159
rect 21453 36119 21511 36125
rect 23750 36116 23756 36168
rect 23808 36116 23814 36168
rect 23934 36116 23940 36168
rect 23992 36116 23998 36168
rect 24026 36116 24032 36168
rect 24084 36116 24090 36168
rect 24576 36159 24634 36165
rect 24576 36125 24588 36159
rect 24622 36156 24634 36159
rect 24854 36156 24860 36168
rect 24622 36128 24860 36156
rect 24622 36125 24634 36128
rect 24576 36119 24634 36125
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 24946 36116 24952 36168
rect 25004 36116 25010 36168
rect 25041 36159 25099 36165
rect 25041 36125 25053 36159
rect 25087 36125 25099 36159
rect 25041 36119 25099 36125
rect 12216 36060 12558 36088
rect 13556 36060 14688 36088
rect 12216 36048 12222 36060
rect 12434 36020 12440 36032
rect 12084 35992 12440 36020
rect 7432 35980 7438 35992
rect 12434 35980 12440 35992
rect 12492 35980 12498 36032
rect 13446 35980 13452 36032
rect 13504 36020 13510 36032
rect 13556 36029 13584 36060
rect 15194 36048 15200 36100
rect 15252 36048 15258 36100
rect 20622 36088 20628 36100
rect 20286 36060 20628 36088
rect 20622 36048 20628 36060
rect 20680 36048 20686 36100
rect 22462 36048 22468 36100
rect 22520 36048 22526 36100
rect 13541 36023 13599 36029
rect 13541 36020 13553 36023
rect 13504 35992 13553 36020
rect 13504 35980 13510 35992
rect 13541 35989 13553 35992
rect 13587 35989 13599 36023
rect 13541 35983 13599 35989
rect 14090 35980 14096 36032
rect 14148 35980 14154 36032
rect 16758 35980 16764 36032
rect 16816 35980 16822 36032
rect 19245 36023 19303 36029
rect 19245 35989 19257 36023
rect 19291 36020 19303 36023
rect 20530 36020 20536 36032
rect 19291 35992 20536 36020
rect 19291 35989 19303 35992
rect 19245 35983 19303 35989
rect 20530 35980 20536 35992
rect 20588 35980 20594 36032
rect 23768 36020 23796 36116
rect 23842 36048 23848 36100
rect 23900 36088 23906 36100
rect 24673 36091 24731 36097
rect 24673 36088 24685 36091
rect 23900 36060 24685 36088
rect 23900 36048 23906 36060
rect 24673 36057 24685 36060
rect 24719 36057 24731 36091
rect 24673 36051 24731 36057
rect 24762 36048 24768 36100
rect 24820 36048 24826 36100
rect 25056 36088 25084 36119
rect 25222 36116 25228 36168
rect 25280 36116 25286 36168
rect 25593 36159 25651 36165
rect 25593 36125 25605 36159
rect 25639 36156 25651 36159
rect 25958 36156 25964 36168
rect 25639 36128 25964 36156
rect 25639 36125 25651 36128
rect 25593 36119 25651 36125
rect 25958 36116 25964 36128
rect 26016 36116 26022 36168
rect 28184 36156 28212 36320
rect 31757 36295 31815 36301
rect 31757 36292 31769 36295
rect 29932 36264 31769 36292
rect 28261 36159 28319 36165
rect 28261 36156 28273 36159
rect 28184 36128 28273 36156
rect 28261 36125 28273 36128
rect 28307 36125 28319 36159
rect 28261 36119 28319 36125
rect 28537 36159 28595 36165
rect 28537 36125 28549 36159
rect 28583 36156 28595 36159
rect 28994 36156 29000 36168
rect 28583 36128 29000 36156
rect 28583 36125 28595 36128
rect 28537 36119 28595 36125
rect 28994 36116 29000 36128
rect 29052 36116 29058 36168
rect 29932 36165 29960 36264
rect 31757 36261 31769 36264
rect 31803 36261 31815 36295
rect 31757 36255 31815 36261
rect 31110 36184 31116 36236
rect 31168 36224 31174 36236
rect 31386 36224 31392 36236
rect 31168 36196 31392 36224
rect 31168 36184 31174 36196
rect 31386 36184 31392 36196
rect 31444 36184 31450 36236
rect 29825 36159 29883 36165
rect 29825 36125 29837 36159
rect 29871 36125 29883 36159
rect 29825 36119 29883 36125
rect 29917 36159 29975 36165
rect 29917 36125 29929 36159
rect 29963 36125 29975 36159
rect 29917 36119 29975 36125
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36156 30343 36159
rect 30377 36159 30435 36165
rect 30377 36156 30389 36159
rect 30331 36128 30389 36156
rect 30331 36125 30343 36128
rect 30285 36119 30343 36125
rect 30377 36125 30389 36128
rect 30423 36125 30435 36159
rect 30377 36119 30435 36125
rect 24964 36060 25084 36088
rect 25240 36088 25268 36116
rect 26786 36088 26792 36100
rect 25240 36060 26792 36088
rect 24964 36020 24992 36060
rect 26786 36048 26792 36060
rect 26844 36088 26850 36100
rect 29362 36088 29368 36100
rect 26844 36060 27002 36088
rect 28000 36060 29368 36088
rect 26844 36048 26850 36060
rect 23768 35992 24992 36020
rect 26896 36020 26924 36060
rect 28000 36020 28028 36060
rect 29362 36048 29368 36060
rect 29420 36048 29426 36100
rect 26896 35992 28028 36020
rect 28074 35980 28080 36032
rect 28132 35980 28138 36032
rect 28445 36023 28503 36029
rect 28445 35989 28457 36023
rect 28491 36020 28503 36023
rect 28534 36020 28540 36032
rect 28491 35992 28540 36020
rect 28491 35989 28503 35992
rect 28445 35983 28503 35989
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 29638 35980 29644 36032
rect 29696 35980 29702 36032
rect 29840 36020 29868 36119
rect 30558 36116 30564 36168
rect 30616 36156 30622 36168
rect 30929 36159 30987 36165
rect 30929 36156 30941 36159
rect 30616 36128 30941 36156
rect 30616 36116 30622 36128
rect 30929 36125 30941 36128
rect 30975 36125 30987 36159
rect 30929 36119 30987 36125
rect 31481 36159 31539 36165
rect 31481 36125 31493 36159
rect 31527 36156 31539 36159
rect 31570 36156 31576 36168
rect 31527 36128 31576 36156
rect 31527 36125 31539 36128
rect 31481 36119 31539 36125
rect 31570 36116 31576 36128
rect 31628 36116 31634 36168
rect 32232 36165 32260 36332
rect 32398 36320 32404 36372
rect 32456 36360 32462 36372
rect 32674 36360 32680 36372
rect 32456 36332 32680 36360
rect 32456 36320 32462 36332
rect 32674 36320 32680 36332
rect 32732 36320 32738 36372
rect 33134 36320 33140 36372
rect 33192 36360 33198 36372
rect 33229 36363 33287 36369
rect 33229 36360 33241 36363
rect 33192 36332 33241 36360
rect 33192 36320 33198 36332
rect 33229 36329 33241 36332
rect 33275 36329 33287 36363
rect 33229 36323 33287 36329
rect 33873 36363 33931 36369
rect 33873 36329 33885 36363
rect 33919 36360 33931 36363
rect 33962 36360 33968 36372
rect 33919 36332 33968 36360
rect 33919 36329 33931 36332
rect 33873 36323 33931 36329
rect 33962 36320 33968 36332
rect 34020 36320 34026 36372
rect 34238 36320 34244 36372
rect 34296 36320 34302 36372
rect 38838 36320 38844 36372
rect 38896 36320 38902 36372
rect 41414 36320 41420 36372
rect 41472 36360 41478 36372
rect 42429 36363 42487 36369
rect 42429 36360 42441 36363
rect 41472 36332 42441 36360
rect 41472 36320 41478 36332
rect 42429 36329 42441 36332
rect 42475 36329 42487 36363
rect 42429 36323 42487 36329
rect 42610 36320 42616 36372
rect 42668 36360 42674 36372
rect 43073 36363 43131 36369
rect 43073 36360 43085 36363
rect 42668 36332 43085 36360
rect 42668 36320 42674 36332
rect 43073 36329 43085 36332
rect 43119 36329 43131 36363
rect 43073 36323 43131 36329
rect 43162 36320 43168 36372
rect 43220 36320 43226 36372
rect 33318 36292 33324 36304
rect 32508 36264 33324 36292
rect 32508 36233 32536 36264
rect 33318 36252 33324 36264
rect 33376 36252 33382 36304
rect 33781 36295 33839 36301
rect 33781 36261 33793 36295
rect 33827 36292 33839 36295
rect 34256 36292 34284 36320
rect 33827 36264 34284 36292
rect 33827 36261 33839 36264
rect 33781 36255 33839 36261
rect 32493 36227 32551 36233
rect 32493 36193 32505 36227
rect 32539 36193 32551 36227
rect 33870 36224 33876 36236
rect 32493 36187 32551 36193
rect 32600 36196 33876 36224
rect 32600 36165 32628 36196
rect 33870 36184 33876 36196
rect 33928 36184 33934 36236
rect 37369 36227 37427 36233
rect 37369 36193 37381 36227
rect 37415 36224 37427 36227
rect 37734 36224 37740 36236
rect 37415 36196 37740 36224
rect 37415 36193 37427 36196
rect 37369 36187 37427 36193
rect 37734 36184 37740 36196
rect 37792 36184 37798 36236
rect 40126 36184 40132 36236
rect 40184 36184 40190 36236
rect 42613 36227 42671 36233
rect 42613 36193 42625 36227
rect 42659 36224 42671 36227
rect 43180 36224 43208 36320
rect 42659 36196 43208 36224
rect 42659 36193 42671 36196
rect 42613 36187 42671 36193
rect 31941 36159 31999 36165
rect 31941 36125 31953 36159
rect 31987 36125 31999 36159
rect 31941 36119 31999 36125
rect 32217 36159 32275 36165
rect 32217 36125 32229 36159
rect 32263 36125 32275 36159
rect 32217 36119 32275 36125
rect 32585 36159 32643 36165
rect 32585 36125 32597 36159
rect 32631 36125 32643 36159
rect 32585 36119 32643 36125
rect 33137 36159 33195 36165
rect 33137 36125 33149 36159
rect 33183 36125 33195 36159
rect 33137 36119 33195 36125
rect 30006 36048 30012 36100
rect 30064 36048 30070 36100
rect 30098 36048 30104 36100
rect 30156 36097 30162 36100
rect 30156 36091 30185 36097
rect 30173 36057 30185 36091
rect 31956 36088 31984 36119
rect 32309 36091 32367 36097
rect 32309 36088 32321 36091
rect 30156 36051 30185 36057
rect 31726 36060 32321 36088
rect 30156 36048 30162 36051
rect 30650 36020 30656 36032
rect 29840 35992 30656 36020
rect 30650 35980 30656 35992
rect 30708 35980 30714 36032
rect 31110 35980 31116 36032
rect 31168 36020 31174 36032
rect 31726 36020 31754 36060
rect 32309 36057 32321 36060
rect 32355 36057 32367 36091
rect 32309 36051 32367 36057
rect 33152 36032 33180 36119
rect 33318 36116 33324 36168
rect 33376 36116 33382 36168
rect 33413 36159 33471 36165
rect 33413 36125 33425 36159
rect 33459 36156 33471 36159
rect 33502 36156 33508 36168
rect 33459 36128 33508 36156
rect 33459 36125 33471 36128
rect 33413 36119 33471 36125
rect 33502 36116 33508 36128
rect 33560 36156 33566 36168
rect 34241 36159 34299 36165
rect 34241 36156 34253 36159
rect 33560 36128 34253 36156
rect 33560 36116 33566 36128
rect 34241 36125 34253 36128
rect 34287 36125 34299 36159
rect 34241 36119 34299 36125
rect 36906 36116 36912 36168
rect 36964 36116 36970 36168
rect 37090 36116 37096 36168
rect 37148 36116 37154 36168
rect 39574 36116 39580 36168
rect 39632 36156 39638 36168
rect 39853 36159 39911 36165
rect 39853 36156 39865 36159
rect 39632 36128 39865 36156
rect 39632 36116 39638 36128
rect 39853 36125 39865 36128
rect 39899 36125 39911 36159
rect 39853 36119 39911 36125
rect 39942 36116 39948 36168
rect 40000 36116 40006 36168
rect 42702 36116 42708 36168
rect 42760 36116 42766 36168
rect 42797 36159 42855 36165
rect 42797 36125 42809 36159
rect 42843 36156 42855 36159
rect 42981 36159 43039 36165
rect 42981 36156 42993 36159
rect 42843 36128 42993 36156
rect 42843 36125 42855 36128
rect 42797 36119 42855 36125
rect 42981 36125 42993 36128
rect 43027 36156 43039 36159
rect 43070 36156 43076 36168
rect 43027 36128 43076 36156
rect 43027 36125 43039 36128
rect 42981 36119 43039 36125
rect 43070 36116 43076 36128
rect 43128 36116 43134 36168
rect 43165 36159 43223 36165
rect 43165 36125 43177 36159
rect 43211 36156 43223 36159
rect 43211 36128 43300 36156
rect 43211 36125 43223 36128
rect 43165 36119 43223 36125
rect 33594 36048 33600 36100
rect 33652 36048 33658 36100
rect 34057 36091 34115 36097
rect 34057 36057 34069 36091
rect 34103 36088 34115 36091
rect 34146 36088 34152 36100
rect 34103 36060 34152 36088
rect 34103 36057 34115 36060
rect 34057 36051 34115 36057
rect 31168 35992 31754 36020
rect 31168 35980 31174 35992
rect 32122 35980 32128 36032
rect 32180 35980 32186 36032
rect 32490 35980 32496 36032
rect 32548 36020 32554 36032
rect 32769 36023 32827 36029
rect 32769 36020 32781 36023
rect 32548 35992 32781 36020
rect 32548 35980 32554 35992
rect 32769 35989 32781 35992
rect 32815 35989 32827 36023
rect 32769 35983 32827 35989
rect 33134 35980 33140 36032
rect 33192 36020 33198 36032
rect 34072 36020 34100 36051
rect 34146 36048 34152 36060
rect 34204 36048 34210 36100
rect 36924 36088 36952 36116
rect 36924 36060 37858 36088
rect 33192 35992 34100 36020
rect 37752 36020 37780 36060
rect 38838 36020 38844 36032
rect 37752 35992 38844 36020
rect 33192 35980 33198 35992
rect 38838 35980 38844 35992
rect 38896 35980 38902 36032
rect 39758 35980 39764 36032
rect 39816 36020 39822 36032
rect 39853 36023 39911 36029
rect 39853 36020 39865 36023
rect 39816 35992 39865 36020
rect 39816 35980 39822 35992
rect 39853 35989 39865 35992
rect 39899 35989 39911 36023
rect 39853 35983 39911 35989
rect 42242 35980 42248 36032
rect 42300 36020 42306 36032
rect 43272 36020 43300 36128
rect 42300 35992 43300 36020
rect 42300 35980 42306 35992
rect 1104 35930 44620 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 44620 35930
rect 1104 35856 44620 35878
rect 2869 35819 2927 35825
rect 2869 35785 2881 35819
rect 2915 35816 2927 35819
rect 4062 35816 4068 35828
rect 2915 35788 4068 35816
rect 2915 35785 2927 35788
rect 2869 35779 2927 35785
rect 4062 35776 4068 35788
rect 4120 35776 4126 35828
rect 5813 35819 5871 35825
rect 5813 35785 5825 35819
rect 5859 35816 5871 35819
rect 6086 35816 6092 35828
rect 5859 35788 6092 35816
rect 5859 35785 5871 35788
rect 5813 35779 5871 35785
rect 6086 35776 6092 35788
rect 6144 35776 6150 35828
rect 7190 35776 7196 35828
rect 7248 35816 7254 35828
rect 7469 35819 7527 35825
rect 7469 35816 7481 35819
rect 7248 35788 7481 35816
rect 7248 35776 7254 35788
rect 7469 35785 7481 35788
rect 7515 35785 7527 35819
rect 7469 35779 7527 35785
rect 12434 35776 12440 35828
rect 12492 35816 12498 35828
rect 12529 35819 12587 35825
rect 12529 35816 12541 35819
rect 12492 35788 12541 35816
rect 12492 35776 12498 35788
rect 12529 35785 12541 35788
rect 12575 35785 12587 35819
rect 12529 35779 12587 35785
rect 13354 35776 13360 35828
rect 13412 35776 13418 35828
rect 13449 35819 13507 35825
rect 13449 35785 13461 35819
rect 13495 35816 13507 35819
rect 14090 35816 14096 35828
rect 13495 35788 14096 35816
rect 13495 35785 13507 35788
rect 13449 35779 13507 35785
rect 14090 35776 14096 35788
rect 14148 35776 14154 35828
rect 14829 35819 14887 35825
rect 14829 35785 14841 35819
rect 14875 35816 14887 35819
rect 15194 35816 15200 35828
rect 14875 35788 15200 35816
rect 14875 35785 14887 35788
rect 14829 35779 14887 35785
rect 15194 35776 15200 35788
rect 15252 35776 15258 35828
rect 15381 35819 15439 35825
rect 15381 35785 15393 35819
rect 15427 35816 15439 35819
rect 16758 35816 16764 35828
rect 15427 35788 16764 35816
rect 15427 35785 15439 35788
rect 15381 35779 15439 35785
rect 16758 35776 16764 35788
rect 16816 35776 16822 35828
rect 16850 35776 16856 35828
rect 16908 35816 16914 35828
rect 17313 35819 17371 35825
rect 17313 35816 17325 35819
rect 16908 35788 17325 35816
rect 16908 35776 16914 35788
rect 17313 35785 17325 35788
rect 17359 35785 17371 35819
rect 17313 35779 17371 35785
rect 20530 35776 20536 35828
rect 20588 35776 20594 35828
rect 22554 35816 22560 35828
rect 21836 35788 22560 35816
rect 5445 35751 5503 35757
rect 5445 35717 5457 35751
rect 5491 35717 5503 35751
rect 5445 35711 5503 35717
rect 2222 35640 2228 35692
rect 2280 35680 2286 35692
rect 2685 35683 2743 35689
rect 2685 35680 2697 35683
rect 2280 35652 2697 35680
rect 2280 35640 2286 35652
rect 2685 35649 2697 35652
rect 2731 35649 2743 35683
rect 5460 35680 5488 35711
rect 5534 35708 5540 35760
rect 5592 35748 5598 35760
rect 5645 35751 5703 35757
rect 5645 35748 5657 35751
rect 5592 35720 5657 35748
rect 5592 35708 5598 35720
rect 5645 35717 5657 35720
rect 5691 35717 5703 35751
rect 13372 35748 13400 35776
rect 13541 35751 13599 35757
rect 13541 35748 13553 35751
rect 13372 35720 13553 35748
rect 5645 35711 5703 35717
rect 13541 35717 13553 35720
rect 13587 35717 13599 35751
rect 13541 35711 13599 35717
rect 15473 35751 15531 35757
rect 15473 35717 15485 35751
rect 15519 35748 15531 35751
rect 15930 35748 15936 35760
rect 15519 35720 15936 35748
rect 15519 35717 15531 35720
rect 15473 35711 15531 35717
rect 15930 35708 15936 35720
rect 15988 35708 15994 35760
rect 20254 35748 20260 35760
rect 17144 35720 20260 35748
rect 6914 35680 6920 35692
rect 5460 35652 6920 35680
rect 2685 35643 2743 35649
rect 6914 35640 6920 35652
rect 6972 35680 6978 35692
rect 7558 35680 7564 35692
rect 6972 35652 7564 35680
rect 6972 35640 6978 35652
rect 7558 35640 7564 35652
rect 7616 35640 7622 35692
rect 7650 35640 7656 35692
rect 7708 35640 7714 35692
rect 12066 35640 12072 35692
rect 12124 35640 12130 35692
rect 12713 35683 12771 35689
rect 12713 35649 12725 35683
rect 12759 35680 12771 35683
rect 14645 35683 14703 35689
rect 12759 35652 13124 35680
rect 12759 35649 12771 35652
rect 12713 35643 12771 35649
rect 13096 35553 13124 35652
rect 14645 35649 14657 35683
rect 14691 35649 14703 35683
rect 14645 35643 14703 35649
rect 13725 35615 13783 35621
rect 13725 35581 13737 35615
rect 13771 35581 13783 35615
rect 13725 35575 13783 35581
rect 13081 35547 13139 35553
rect 13081 35513 13093 35547
rect 13127 35513 13139 35547
rect 13081 35507 13139 35513
rect 5626 35436 5632 35488
rect 5684 35436 5690 35488
rect 12161 35479 12219 35485
rect 12161 35445 12173 35479
rect 12207 35476 12219 35479
rect 12802 35476 12808 35488
rect 12207 35448 12808 35476
rect 12207 35445 12219 35448
rect 12161 35439 12219 35445
rect 12802 35436 12808 35448
rect 12860 35436 12866 35488
rect 13740 35476 13768 35575
rect 14660 35544 14688 35643
rect 16758 35640 16764 35692
rect 16816 35680 16822 35692
rect 17144 35689 17172 35720
rect 20254 35708 20260 35720
rect 20312 35708 20318 35760
rect 17129 35683 17187 35689
rect 17129 35680 17141 35683
rect 16816 35652 17141 35680
rect 16816 35640 16822 35652
rect 17129 35649 17141 35652
rect 17175 35649 17187 35683
rect 17129 35643 17187 35649
rect 20441 35683 20499 35689
rect 20441 35649 20453 35683
rect 20487 35680 20499 35683
rect 20548 35680 20576 35776
rect 20487 35652 20576 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 15565 35615 15623 35621
rect 15565 35612 15577 35615
rect 15488 35584 15577 35612
rect 15013 35547 15071 35553
rect 15013 35544 15025 35547
rect 14660 35516 15025 35544
rect 15013 35513 15025 35516
rect 15059 35513 15071 35547
rect 15013 35507 15071 35513
rect 15488 35476 15516 35584
rect 15565 35581 15577 35584
rect 15611 35581 15623 35615
rect 15565 35575 15623 35581
rect 18598 35572 18604 35624
rect 18656 35572 18662 35624
rect 19242 35612 19248 35624
rect 18892 35584 19248 35612
rect 18892 35544 18920 35584
rect 19242 35572 19248 35584
rect 19300 35572 19306 35624
rect 21836 35553 21864 35788
rect 22554 35776 22560 35788
rect 22612 35776 22618 35828
rect 24946 35776 24952 35828
rect 25004 35816 25010 35828
rect 25501 35819 25559 35825
rect 25501 35816 25513 35819
rect 25004 35788 25513 35816
rect 25004 35776 25010 35788
rect 25501 35785 25513 35788
rect 25547 35785 25559 35819
rect 25501 35779 25559 35785
rect 27062 35776 27068 35828
rect 27120 35816 27126 35828
rect 27157 35819 27215 35825
rect 27157 35816 27169 35819
rect 27120 35788 27169 35816
rect 27120 35776 27126 35788
rect 27157 35785 27169 35788
rect 27203 35785 27215 35819
rect 27157 35779 27215 35785
rect 27325 35819 27383 35825
rect 27325 35785 27337 35819
rect 27371 35816 27383 35819
rect 28074 35816 28080 35828
rect 27371 35788 28080 35816
rect 27371 35785 27383 35788
rect 27325 35779 27383 35785
rect 28074 35776 28080 35788
rect 28132 35776 28138 35828
rect 29638 35816 29644 35828
rect 28920 35788 29644 35816
rect 21928 35720 22126 35748
rect 21821 35547 21879 35553
rect 21821 35544 21833 35547
rect 18064 35516 18920 35544
rect 18984 35516 21833 35544
rect 18064 35488 18092 35516
rect 18984 35488 19012 35516
rect 21821 35513 21833 35516
rect 21867 35513 21879 35547
rect 21821 35507 21879 35513
rect 18046 35476 18052 35488
rect 13740 35448 18052 35476
rect 18046 35436 18052 35448
rect 18104 35436 18110 35488
rect 18966 35436 18972 35488
rect 19024 35436 19030 35488
rect 19153 35479 19211 35485
rect 19153 35445 19165 35479
rect 19199 35476 19211 35479
rect 19242 35476 19248 35488
rect 19199 35448 19248 35476
rect 19199 35445 19211 35448
rect 19153 35439 19211 35445
rect 19242 35436 19248 35448
rect 19300 35436 19306 35488
rect 20349 35479 20407 35485
rect 20349 35445 20361 35479
rect 20395 35476 20407 35479
rect 20438 35476 20444 35488
rect 20395 35448 20444 35476
rect 20395 35445 20407 35448
rect 20349 35439 20407 35445
rect 20438 35436 20444 35448
rect 20496 35436 20502 35488
rect 20622 35436 20628 35488
rect 20680 35476 20686 35488
rect 21928 35476 21956 35720
rect 25958 35708 25964 35760
rect 26016 35748 26022 35760
rect 26329 35751 26387 35757
rect 26329 35748 26341 35751
rect 26016 35720 26341 35748
rect 26016 35708 26022 35720
rect 26329 35717 26341 35720
rect 26375 35717 26387 35751
rect 26329 35711 26387 35717
rect 26418 35708 26424 35760
rect 26476 35748 26482 35760
rect 27525 35751 27583 35757
rect 27525 35748 27537 35751
rect 26476 35720 27537 35748
rect 26476 35708 26482 35720
rect 27525 35717 27537 35720
rect 27571 35717 27583 35751
rect 27890 35748 27896 35760
rect 27525 35711 27583 35717
rect 27816 35720 27896 35748
rect 23566 35640 23572 35692
rect 23624 35640 23630 35692
rect 22094 35572 22100 35624
rect 22152 35612 22158 35624
rect 23293 35615 23351 35621
rect 23293 35612 23305 35615
rect 22152 35584 23305 35612
rect 22152 35572 22158 35584
rect 23293 35581 23305 35584
rect 23339 35581 23351 35615
rect 23293 35575 23351 35581
rect 26050 35572 26056 35624
rect 26108 35572 26114 35624
rect 27540 35544 27568 35711
rect 27816 35689 27844 35720
rect 27890 35708 27896 35720
rect 27948 35708 27954 35760
rect 28920 35757 28948 35788
rect 29638 35776 29644 35788
rect 29696 35776 29702 35828
rect 30377 35819 30435 35825
rect 30377 35785 30389 35819
rect 30423 35816 30435 35819
rect 30558 35816 30564 35828
rect 30423 35788 30564 35816
rect 30423 35785 30435 35788
rect 30377 35779 30435 35785
rect 30558 35776 30564 35788
rect 30616 35776 30622 35828
rect 30650 35776 30656 35828
rect 30708 35776 30714 35828
rect 31389 35819 31447 35825
rect 31389 35816 31401 35819
rect 30760 35788 31401 35816
rect 28905 35751 28963 35757
rect 28905 35717 28917 35751
rect 28951 35717 28963 35751
rect 28905 35711 28963 35717
rect 29362 35708 29368 35760
rect 29420 35708 29426 35760
rect 30760 35748 30788 35788
rect 31389 35785 31401 35788
rect 31435 35816 31447 35819
rect 31754 35816 31760 35828
rect 31435 35788 31760 35816
rect 31435 35785 31447 35788
rect 31389 35779 31447 35785
rect 31754 35776 31760 35788
rect 31812 35816 31818 35828
rect 32122 35816 32128 35828
rect 31812 35788 32128 35816
rect 31812 35776 31818 35788
rect 32122 35776 32128 35788
rect 32180 35776 32186 35828
rect 39758 35816 39764 35828
rect 32692 35788 33364 35816
rect 30668 35720 30788 35748
rect 30929 35751 30987 35757
rect 27801 35683 27859 35689
rect 27801 35649 27813 35683
rect 27847 35649 27859 35683
rect 27801 35643 27859 35649
rect 27985 35683 28043 35689
rect 27985 35649 27997 35683
rect 28031 35680 28043 35683
rect 28166 35680 28172 35692
rect 28031 35652 28172 35680
rect 28031 35649 28043 35652
rect 27985 35643 28043 35649
rect 28166 35640 28172 35652
rect 28224 35640 28230 35692
rect 28445 35683 28503 35689
rect 28445 35649 28457 35683
rect 28491 35680 28503 35683
rect 28534 35680 28540 35692
rect 28491 35652 28540 35680
rect 28491 35649 28503 35652
rect 28445 35643 28503 35649
rect 28534 35640 28540 35652
rect 28592 35640 28598 35692
rect 30668 35689 30696 35720
rect 30929 35717 30941 35751
rect 30975 35748 30987 35751
rect 31110 35748 31116 35760
rect 30975 35720 31116 35748
rect 30975 35717 30987 35720
rect 30929 35711 30987 35717
rect 31110 35708 31116 35720
rect 31168 35708 31174 35760
rect 31202 35708 31208 35760
rect 31260 35708 31266 35760
rect 31662 35708 31668 35760
rect 31720 35748 31726 35760
rect 31720 35720 32168 35748
rect 31720 35708 31726 35720
rect 30653 35683 30711 35689
rect 30653 35649 30665 35683
rect 30699 35649 30711 35683
rect 30653 35643 30711 35649
rect 30745 35683 30803 35689
rect 30745 35649 30757 35683
rect 30791 35680 30803 35683
rect 31220 35680 31248 35708
rect 30791 35652 31248 35680
rect 31297 35683 31355 35689
rect 30791 35649 30803 35652
rect 30745 35643 30803 35649
rect 31297 35649 31309 35683
rect 31343 35649 31355 35683
rect 31297 35643 31355 35649
rect 27890 35572 27896 35624
rect 27948 35572 27954 35624
rect 28077 35615 28135 35621
rect 28077 35581 28089 35615
rect 28123 35612 28135 35615
rect 28353 35615 28411 35621
rect 28353 35612 28365 35615
rect 28123 35584 28365 35612
rect 28123 35581 28135 35584
rect 28077 35575 28135 35581
rect 28353 35581 28365 35584
rect 28399 35581 28411 35615
rect 28353 35575 28411 35581
rect 28626 35572 28632 35624
rect 28684 35572 28690 35624
rect 31312 35612 31340 35643
rect 31386 35640 31392 35692
rect 31444 35680 31450 35692
rect 32140 35689 32168 35720
rect 32582 35708 32588 35760
rect 32640 35708 32646 35760
rect 32306 35689 32312 35692
rect 31481 35683 31539 35689
rect 31481 35680 31493 35683
rect 31444 35652 31493 35680
rect 31444 35640 31450 35652
rect 31481 35649 31493 35652
rect 31527 35680 31539 35683
rect 31573 35683 31631 35689
rect 31573 35680 31585 35683
rect 31527 35652 31585 35680
rect 31527 35649 31539 35652
rect 31481 35643 31539 35649
rect 31573 35649 31585 35652
rect 31619 35649 31631 35683
rect 31573 35643 31631 35649
rect 31757 35683 31815 35689
rect 31757 35649 31769 35683
rect 31803 35649 31815 35683
rect 31757 35643 31815 35649
rect 32125 35683 32183 35689
rect 32125 35649 32137 35683
rect 32171 35649 32183 35683
rect 32290 35683 32312 35689
rect 32290 35680 32302 35683
rect 32125 35643 32183 35649
rect 32232 35652 32302 35680
rect 31772 35612 31800 35643
rect 32232 35612 32260 35652
rect 32290 35649 32302 35652
rect 32290 35643 32312 35649
rect 32306 35640 32312 35643
rect 32364 35640 32370 35692
rect 32692 35689 32720 35788
rect 33336 35760 33364 35788
rect 39684 35788 39764 35816
rect 33226 35708 33232 35760
rect 33284 35708 33290 35760
rect 33318 35708 33324 35760
rect 33376 35708 33382 35760
rect 36906 35748 36912 35760
rect 35650 35720 36912 35748
rect 36906 35708 36912 35720
rect 36964 35708 36970 35760
rect 39684 35757 39712 35788
rect 39758 35776 39764 35788
rect 39816 35776 39822 35828
rect 39669 35751 39727 35757
rect 39669 35717 39681 35751
rect 39715 35717 39727 35751
rect 39669 35711 39727 35717
rect 32677 35683 32735 35689
rect 32677 35680 32689 35683
rect 32416 35652 32689 35680
rect 31312 35584 32260 35612
rect 27540 35516 27752 35544
rect 20680 35448 21956 35476
rect 26605 35479 26663 35485
rect 20680 35436 20686 35448
rect 26605 35445 26617 35479
rect 26651 35476 26663 35479
rect 26786 35476 26792 35488
rect 26651 35448 26792 35476
rect 26651 35445 26663 35448
rect 26605 35439 26663 35445
rect 26786 35436 26792 35448
rect 26844 35436 26850 35488
rect 27341 35479 27399 35485
rect 27341 35445 27353 35479
rect 27387 35476 27399 35479
rect 27522 35476 27528 35488
rect 27387 35448 27528 35476
rect 27387 35445 27399 35448
rect 27341 35439 27399 35445
rect 27522 35436 27528 35448
rect 27580 35436 27586 35488
rect 27614 35436 27620 35488
rect 27672 35436 27678 35488
rect 27724 35476 27752 35516
rect 31386 35504 31392 35556
rect 31444 35544 31450 35556
rect 32416 35544 32444 35652
rect 32677 35649 32689 35652
rect 32723 35649 32735 35683
rect 32677 35643 32735 35649
rect 33413 35683 33471 35689
rect 33413 35649 33425 35683
rect 33459 35649 33471 35683
rect 33413 35643 33471 35649
rect 33428 35612 33456 35643
rect 33502 35640 33508 35692
rect 33560 35640 33566 35692
rect 40802 35666 42656 35680
rect 40788 35652 42656 35666
rect 33594 35612 33600 35624
rect 32508 35584 33600 35612
rect 32508 35553 32536 35584
rect 33594 35572 33600 35584
rect 33652 35612 33658 35624
rect 33652 35584 34468 35612
rect 33652 35572 33658 35584
rect 31444 35516 32444 35544
rect 32493 35547 32551 35553
rect 31444 35504 31450 35516
rect 32493 35513 32505 35547
rect 32539 35513 32551 35547
rect 32493 35507 32551 35513
rect 34440 35488 34468 35584
rect 36078 35572 36084 35624
rect 36136 35572 36142 35624
rect 36354 35572 36360 35624
rect 36412 35612 36418 35624
rect 37090 35612 37096 35624
rect 36412 35584 37096 35612
rect 36412 35572 36418 35584
rect 37090 35572 37096 35584
rect 37148 35612 37154 35624
rect 39390 35612 39396 35624
rect 37148 35584 39396 35612
rect 37148 35572 37154 35584
rect 39390 35572 39396 35584
rect 39448 35572 39454 35624
rect 40788 35612 40816 35652
rect 39500 35584 40816 35612
rect 38838 35504 38844 35556
rect 38896 35544 38902 35556
rect 39500 35544 39528 35584
rect 40954 35572 40960 35624
rect 41012 35612 41018 35624
rect 41141 35615 41199 35621
rect 41141 35612 41153 35615
rect 41012 35584 41153 35612
rect 41012 35572 41018 35584
rect 41141 35581 41153 35584
rect 41187 35612 41199 35615
rect 41785 35615 41843 35621
rect 41785 35612 41797 35615
rect 41187 35584 41797 35612
rect 41187 35581 41199 35584
rect 41141 35575 41199 35581
rect 41785 35581 41797 35584
rect 41831 35581 41843 35615
rect 41785 35575 41843 35581
rect 38896 35516 39528 35544
rect 38896 35504 38902 35516
rect 42628 35488 42656 35652
rect 31846 35476 31852 35488
rect 27724 35448 31852 35476
rect 31846 35436 31852 35448
rect 31904 35436 31910 35488
rect 31938 35436 31944 35488
rect 31996 35436 32002 35488
rect 32401 35479 32459 35485
rect 32401 35445 32413 35479
rect 32447 35476 32459 35479
rect 33134 35476 33140 35488
rect 32447 35448 33140 35476
rect 32447 35445 32459 35448
rect 32401 35439 32459 35445
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 34422 35436 34428 35488
rect 34480 35476 34486 35488
rect 34609 35479 34667 35485
rect 34609 35476 34621 35479
rect 34480 35448 34621 35476
rect 34480 35436 34486 35448
rect 34609 35445 34621 35448
rect 34655 35445 34667 35479
rect 34609 35439 34667 35445
rect 39390 35436 39396 35488
rect 39448 35476 39454 35488
rect 39850 35476 39856 35488
rect 39448 35448 39856 35476
rect 39448 35436 39454 35448
rect 39850 35436 39856 35448
rect 39908 35436 39914 35488
rect 40126 35436 40132 35488
rect 40184 35476 40190 35488
rect 41233 35479 41291 35485
rect 41233 35476 41245 35479
rect 40184 35448 41245 35476
rect 40184 35436 40190 35448
rect 41233 35445 41245 35448
rect 41279 35445 41291 35479
rect 41233 35439 41291 35445
rect 42610 35436 42616 35488
rect 42668 35436 42674 35488
rect 1104 35386 44620 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 44620 35386
rect 1104 35312 44620 35334
rect 5534 35272 5540 35284
rect 5368 35244 5540 35272
rect 5074 35028 5080 35080
rect 5132 35068 5138 35080
rect 5368 35077 5396 35244
rect 5534 35232 5540 35244
rect 5592 35272 5598 35284
rect 6086 35272 6092 35284
rect 5592 35244 6092 35272
rect 5592 35232 5598 35244
rect 6086 35232 6092 35244
rect 6144 35232 6150 35284
rect 7650 35232 7656 35284
rect 7708 35232 7714 35284
rect 7837 35275 7895 35281
rect 7837 35241 7849 35275
rect 7883 35272 7895 35275
rect 8113 35275 8171 35281
rect 8113 35272 8125 35275
rect 7883 35244 8125 35272
rect 7883 35241 7895 35244
rect 7837 35235 7895 35241
rect 8113 35241 8125 35244
rect 8159 35241 8171 35275
rect 14274 35272 14280 35284
rect 8113 35235 8171 35241
rect 8404 35244 14280 35272
rect 5442 35164 5448 35216
rect 5500 35204 5506 35216
rect 5500 35176 5672 35204
rect 5500 35164 5506 35176
rect 5241 35071 5299 35077
rect 5241 35068 5253 35071
rect 5132 35040 5253 35068
rect 5132 35028 5138 35040
rect 5241 35037 5253 35040
rect 5287 35037 5299 35071
rect 5241 35031 5299 35037
rect 5353 35071 5411 35077
rect 5353 35037 5365 35071
rect 5399 35037 5411 35071
rect 5353 35031 5411 35037
rect 5445 35071 5503 35077
rect 5445 35037 5457 35071
rect 5491 35068 5503 35071
rect 5534 35068 5540 35080
rect 5491 35040 5540 35068
rect 5491 35037 5503 35040
rect 5445 35031 5503 35037
rect 5534 35028 5540 35040
rect 5592 35028 5598 35080
rect 5644 35077 5672 35176
rect 7466 35164 7472 35216
rect 7524 35204 7530 35216
rect 8404 35204 8432 35244
rect 14274 35232 14280 35244
rect 14332 35272 14338 35284
rect 15562 35272 15568 35284
rect 14332 35244 15568 35272
rect 14332 35232 14338 35244
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 16206 35232 16212 35284
rect 16264 35232 16270 35284
rect 16945 35275 17003 35281
rect 16945 35241 16957 35275
rect 16991 35272 17003 35275
rect 16991 35244 18552 35272
rect 16991 35241 17003 35244
rect 16945 35235 17003 35241
rect 7524 35176 8432 35204
rect 7524 35164 7530 35176
rect 8478 35164 8484 35216
rect 8536 35204 8542 35216
rect 11425 35207 11483 35213
rect 8536 35176 9352 35204
rect 8536 35164 8542 35176
rect 5721 35139 5779 35145
rect 5721 35105 5733 35139
rect 5767 35136 5779 35139
rect 6730 35136 6736 35148
rect 5767 35108 6736 35136
rect 5767 35105 5779 35108
rect 5721 35099 5779 35105
rect 6730 35096 6736 35108
rect 6788 35096 6794 35148
rect 8294 35096 8300 35148
rect 8352 35136 8358 35148
rect 9324 35136 9352 35176
rect 11425 35173 11437 35207
rect 11471 35204 11483 35207
rect 11471 35176 12434 35204
rect 11471 35173 11483 35176
rect 11425 35167 11483 35173
rect 12250 35136 12256 35148
rect 8352 35108 9168 35136
rect 8352 35096 8358 35108
rect 5629 35071 5687 35077
rect 5629 35037 5641 35071
rect 5675 35037 5687 35071
rect 7374 35068 7380 35080
rect 7130 35040 7380 35068
rect 5629 35031 5687 35037
rect 7374 35028 7380 35040
rect 7432 35028 7438 35080
rect 8481 35071 8539 35077
rect 8481 35068 8493 35071
rect 7484 35040 8493 35068
rect 4985 35003 5043 35009
rect 4985 34969 4997 35003
rect 5031 35000 5043 35003
rect 5997 35003 6055 35009
rect 5997 35000 6009 35003
rect 5031 34972 6009 35000
rect 5031 34969 5043 34972
rect 4985 34963 5043 34969
rect 5997 34969 6009 34972
rect 6043 34969 6055 35003
rect 5997 34963 6055 34969
rect 6730 34892 6736 34944
rect 6788 34932 6794 34944
rect 7484 34932 7512 35040
rect 8481 35037 8493 35040
rect 8527 35070 8539 35071
rect 8573 35071 8631 35077
rect 8573 35070 8585 35071
rect 8527 35042 8585 35070
rect 8527 35037 8539 35042
rect 8481 35031 8539 35037
rect 8573 35037 8585 35042
rect 8619 35037 8631 35071
rect 8757 35071 8815 35077
rect 8757 35068 8769 35071
rect 8573 35031 8631 35037
rect 8680 35040 8769 35068
rect 7558 34960 7564 35012
rect 7616 35000 7622 35012
rect 8021 35003 8079 35009
rect 8021 35000 8033 35003
rect 7616 34972 8033 35000
rect 7616 34960 7622 34972
rect 8021 34969 8033 34972
rect 8067 34969 8079 35003
rect 8021 34963 8079 34969
rect 8297 35003 8355 35009
rect 8297 34969 8309 35003
rect 8343 35000 8355 35003
rect 8680 35000 8708 35040
rect 8757 35037 8769 35040
rect 8803 35068 8815 35071
rect 8846 35068 8852 35080
rect 8803 35040 8852 35068
rect 8803 35037 8815 35040
rect 8757 35031 8815 35037
rect 8846 35028 8852 35040
rect 8904 35028 8910 35080
rect 8938 35028 8944 35080
rect 8996 35028 9002 35080
rect 9140 35077 9168 35108
rect 9324 35108 12256 35136
rect 9324 35077 9352 35108
rect 12250 35096 12256 35108
rect 12308 35096 12314 35148
rect 12406 35136 12434 35176
rect 16224 35136 16252 35232
rect 18524 35204 18552 35244
rect 18598 35232 18604 35284
rect 18656 35272 18662 35284
rect 18785 35275 18843 35281
rect 18785 35272 18797 35275
rect 18656 35244 18797 35272
rect 18656 35232 18662 35244
rect 18785 35241 18797 35244
rect 18831 35241 18843 35275
rect 23750 35272 23756 35284
rect 18785 35235 18843 35241
rect 19352 35244 23756 35272
rect 19352 35204 19380 35244
rect 23750 35232 23756 35244
rect 23808 35232 23814 35284
rect 25958 35232 25964 35284
rect 26016 35272 26022 35284
rect 26053 35275 26111 35281
rect 26053 35272 26065 35275
rect 26016 35244 26065 35272
rect 26016 35232 26022 35244
rect 26053 35241 26065 35244
rect 26099 35241 26111 35275
rect 26053 35235 26111 35241
rect 31938 35232 31944 35284
rect 31996 35232 32002 35284
rect 36354 35272 36360 35284
rect 35912 35244 36360 35272
rect 18524 35176 19380 35204
rect 12406 35108 16252 35136
rect 9125 35071 9183 35077
rect 9125 35037 9137 35071
rect 9171 35037 9183 35071
rect 9125 35031 9183 35037
rect 9217 35071 9275 35077
rect 9217 35037 9229 35071
rect 9263 35037 9275 35071
rect 9217 35031 9275 35037
rect 9309 35071 9367 35077
rect 9309 35037 9321 35071
rect 9355 35037 9367 35071
rect 9309 35031 9367 35037
rect 8343 34972 8708 35000
rect 8343 34969 8355 34972
rect 8297 34963 8355 34969
rect 6788 34904 7512 34932
rect 7821 34935 7879 34941
rect 6788 34892 6794 34904
rect 7821 34901 7833 34935
rect 7867 34932 7879 34935
rect 8662 34932 8668 34944
rect 7867 34904 8668 34932
rect 7867 34901 7879 34904
rect 7821 34895 7879 34901
rect 8662 34892 8668 34904
rect 8720 34932 8726 34944
rect 8757 34935 8815 34941
rect 8757 34932 8769 34935
rect 8720 34904 8769 34932
rect 8720 34892 8726 34904
rect 8757 34901 8769 34904
rect 8803 34932 8815 34935
rect 9232 34932 9260 35031
rect 9398 35028 9404 35080
rect 9456 35068 9462 35080
rect 9677 35071 9735 35077
rect 9677 35068 9689 35071
rect 9456 35040 9689 35068
rect 9456 35028 9462 35040
rect 9677 35037 9689 35040
rect 9723 35037 9735 35071
rect 9677 35031 9735 35037
rect 11054 35028 11060 35080
rect 11112 35068 11118 35080
rect 12618 35068 12624 35080
rect 11112 35040 12624 35068
rect 11112 35028 11118 35040
rect 12618 35028 12624 35040
rect 12676 35028 12682 35080
rect 14568 35077 14596 35108
rect 16850 35096 16856 35148
rect 16908 35096 16914 35148
rect 16942 35096 16948 35148
rect 17000 35136 17006 35148
rect 17037 35139 17095 35145
rect 17037 35136 17049 35139
rect 17000 35108 17049 35136
rect 17000 35096 17006 35108
rect 17037 35105 17049 35108
rect 17083 35136 17095 35139
rect 19245 35139 19303 35145
rect 19245 35136 19257 35139
rect 17083 35108 19257 35136
rect 17083 35105 17095 35108
rect 17037 35099 17095 35105
rect 19245 35105 19257 35108
rect 19291 35105 19303 35139
rect 19245 35099 19303 35105
rect 20254 35096 20260 35148
rect 20312 35136 20318 35148
rect 26418 35136 26424 35148
rect 20312 35108 25728 35136
rect 20312 35096 20318 35108
rect 14553 35071 14611 35077
rect 14553 35037 14565 35071
rect 14599 35037 14611 35071
rect 16301 35071 16359 35077
rect 16301 35068 16313 35071
rect 14553 35031 14611 35037
rect 16224 35040 16313 35068
rect 9585 35003 9643 35009
rect 9585 34969 9597 35003
rect 9631 35000 9643 35003
rect 9953 35003 10011 35009
rect 9953 35000 9965 35003
rect 9631 34972 9965 35000
rect 9631 34969 9643 34972
rect 9585 34963 9643 34969
rect 9953 34969 9965 34972
rect 9999 34969 10011 35003
rect 9953 34963 10011 34969
rect 16224 34944 16252 35040
rect 16301 35037 16313 35040
rect 16347 35068 16359 35071
rect 16577 35071 16635 35077
rect 16577 35068 16589 35071
rect 16347 35040 16589 35068
rect 16347 35037 16359 35040
rect 16301 35031 16359 35037
rect 16577 35037 16589 35040
rect 16623 35037 16635 35071
rect 16577 35031 16635 35037
rect 16761 35071 16819 35077
rect 16761 35037 16773 35071
rect 16807 35068 16819 35071
rect 16868 35068 16896 35096
rect 16807 35040 16896 35068
rect 16807 35037 16819 35040
rect 16761 35031 16819 35037
rect 18414 35028 18420 35080
rect 18472 35028 18478 35080
rect 18874 35028 18880 35080
rect 18932 35028 18938 35080
rect 20622 35028 20628 35080
rect 20680 35028 20686 35080
rect 23482 35077 23510 35108
rect 25700 35080 25728 35108
rect 26160 35108 26424 35136
rect 22557 35071 22615 35077
rect 22557 35037 22569 35071
rect 22603 35068 22615 35071
rect 23477 35071 23535 35077
rect 22603 35040 23428 35068
rect 22603 35037 22615 35040
rect 22557 35031 22615 35037
rect 17310 34960 17316 35012
rect 17368 34960 17374 35012
rect 19521 35003 19579 35009
rect 19521 35000 19533 35003
rect 19076 34972 19533 35000
rect 8803 34904 9260 34932
rect 8803 34901 8815 34904
rect 8757 34895 8815 34901
rect 12250 34892 12256 34944
rect 12308 34932 12314 34944
rect 14461 34935 14519 34941
rect 14461 34932 14473 34935
rect 12308 34904 14473 34932
rect 12308 34892 12314 34904
rect 14461 34901 14473 34904
rect 14507 34932 14519 34935
rect 14826 34932 14832 34944
rect 14507 34904 14832 34932
rect 14507 34901 14519 34904
rect 14461 34895 14519 34901
rect 14826 34892 14832 34904
rect 14884 34892 14890 34944
rect 15746 34892 15752 34944
rect 15804 34892 15810 34944
rect 16206 34892 16212 34944
rect 16264 34892 16270 34944
rect 19076 34941 19104 34972
rect 19521 34969 19533 34972
rect 19567 34969 19579 35003
rect 22738 35000 22744 35012
rect 19521 34963 19579 34969
rect 22572 34972 22744 35000
rect 22572 34944 22600 34972
rect 22738 34960 22744 34972
rect 22796 35000 22802 35012
rect 23201 35003 23259 35009
rect 23201 35000 23213 35003
rect 22796 34972 23213 35000
rect 22796 34960 22802 34972
rect 23201 34969 23213 34972
rect 23247 34969 23259 35003
rect 23400 35000 23428 35040
rect 23477 35037 23489 35071
rect 23523 35037 23535 35071
rect 23477 35031 23535 35037
rect 25038 35028 25044 35080
rect 25096 35028 25102 35080
rect 25682 35028 25688 35080
rect 25740 35028 25746 35080
rect 26160 35000 26188 35108
rect 26418 35096 26424 35108
rect 26476 35096 26482 35148
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35068 26295 35071
rect 26283 35040 27660 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 23400 34972 26188 35000
rect 23201 34963 23259 34969
rect 27632 34944 27660 35040
rect 31754 35028 31760 35080
rect 31812 35028 31818 35080
rect 31956 35077 31984 35232
rect 34422 35096 34428 35148
rect 34480 35136 34486 35148
rect 35912 35145 35940 35244
rect 36354 35232 36360 35244
rect 36412 35232 36418 35284
rect 39574 35232 39580 35284
rect 39632 35232 39638 35284
rect 39669 35275 39727 35281
rect 39669 35241 39681 35275
rect 39715 35272 39727 35275
rect 39942 35272 39948 35284
rect 39715 35244 39948 35272
rect 39715 35241 39727 35244
rect 39669 35235 39727 35241
rect 39942 35232 39948 35244
rect 40000 35232 40006 35284
rect 40037 35275 40095 35281
rect 40037 35241 40049 35275
rect 40083 35272 40095 35275
rect 40954 35272 40960 35284
rect 40083 35244 40960 35272
rect 40083 35241 40095 35244
rect 40037 35235 40095 35241
rect 40954 35232 40960 35244
rect 41012 35232 41018 35284
rect 41138 35232 41144 35284
rect 41196 35232 41202 35284
rect 39592 35204 39620 35232
rect 39850 35204 39856 35216
rect 39592 35176 39856 35204
rect 39850 35164 39856 35176
rect 39908 35164 39914 35216
rect 40126 35164 40132 35216
rect 40184 35164 40190 35216
rect 40405 35207 40463 35213
rect 40405 35204 40417 35207
rect 40236 35176 40417 35204
rect 34977 35139 35035 35145
rect 34977 35136 34989 35139
rect 34480 35108 34989 35136
rect 34480 35096 34486 35108
rect 34977 35105 34989 35108
rect 35023 35105 35035 35139
rect 34977 35099 35035 35105
rect 35897 35139 35955 35145
rect 35897 35105 35909 35139
rect 35943 35105 35955 35139
rect 35897 35099 35955 35105
rect 38746 35096 38752 35148
rect 38804 35096 38810 35148
rect 39209 35139 39267 35145
rect 39209 35105 39221 35139
rect 39255 35136 39267 35139
rect 40144 35136 40172 35164
rect 39255 35108 39436 35136
rect 39255 35105 39267 35108
rect 39209 35099 39267 35105
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35037 31999 35071
rect 31941 35031 31999 35037
rect 32030 35028 32036 35080
rect 32088 35068 32094 35080
rect 35802 35068 35808 35080
rect 32088 35040 35808 35068
rect 32088 35028 32094 35040
rect 35802 35028 35808 35040
rect 35860 35028 35866 35080
rect 39114 35028 39120 35080
rect 39172 35028 39178 35080
rect 39408 35077 39436 35108
rect 39684 35108 40172 35136
rect 39684 35077 39712 35108
rect 39393 35071 39451 35077
rect 39393 35037 39405 35071
rect 39439 35037 39451 35071
rect 39393 35031 39451 35037
rect 39672 35071 39730 35077
rect 39672 35037 39684 35071
rect 39718 35037 39730 35071
rect 39672 35031 39730 35037
rect 31849 35003 31907 35009
rect 31849 34969 31861 35003
rect 31895 35000 31907 35003
rect 32398 35000 32404 35012
rect 31895 34972 32404 35000
rect 31895 34969 31907 34972
rect 31849 34963 31907 34969
rect 32398 34960 32404 34972
rect 32456 34960 32462 35012
rect 32508 34972 35894 35000
rect 19061 34935 19119 34941
rect 19061 34901 19073 34935
rect 19107 34901 19119 34935
rect 19061 34895 19119 34901
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 20993 34935 21051 34941
rect 20993 34932 21005 34935
rect 19392 34904 21005 34932
rect 19392 34892 19398 34904
rect 20993 34901 21005 34904
rect 21039 34901 21051 34935
rect 20993 34895 21051 34901
rect 22554 34892 22560 34944
rect 22612 34892 22618 34944
rect 22833 34935 22891 34941
rect 22833 34901 22845 34935
rect 22879 34932 22891 34935
rect 24026 34932 24032 34944
rect 22879 34904 24032 34932
rect 22879 34901 22891 34904
rect 22833 34895 22891 34901
rect 24026 34892 24032 34904
rect 24084 34892 24090 34944
rect 24486 34892 24492 34944
rect 24544 34892 24550 34944
rect 27614 34892 27620 34944
rect 27672 34932 27678 34944
rect 32508 34932 32536 34972
rect 27672 34904 32536 34932
rect 27672 34892 27678 34904
rect 35342 34892 35348 34944
rect 35400 34932 35406 34944
rect 35621 34935 35679 34941
rect 35621 34932 35633 34935
rect 35400 34904 35633 34932
rect 35400 34892 35406 34904
rect 35621 34901 35633 34904
rect 35667 34901 35679 34935
rect 35866 34932 35894 34972
rect 36170 34960 36176 35012
rect 36228 34960 36234 35012
rect 36906 34960 36912 35012
rect 36964 34960 36970 35012
rect 39408 35000 39436 35031
rect 39758 35028 39764 35080
rect 39816 35068 39822 35080
rect 40236 35068 40264 35176
rect 40405 35173 40417 35176
rect 40451 35173 40463 35207
rect 40405 35167 40463 35173
rect 40972 35145 41000 35232
rect 40957 35139 41015 35145
rect 40957 35105 40969 35139
rect 41003 35105 41015 35139
rect 40957 35099 41015 35105
rect 42702 35096 42708 35148
rect 42760 35096 42766 35148
rect 39816 35040 40264 35068
rect 39816 35028 39822 35040
rect 40236 35009 40264 35040
rect 40862 35028 40868 35080
rect 40920 35028 40926 35080
rect 42242 35028 42248 35080
rect 42300 35068 42306 35080
rect 43349 35071 43407 35077
rect 43349 35068 43361 35071
rect 42300 35040 43361 35068
rect 42300 35028 42306 35040
rect 43349 35037 43361 35040
rect 43395 35037 43407 35071
rect 43349 35031 43407 35037
rect 43438 35028 43444 35080
rect 43496 35068 43502 35080
rect 43533 35071 43591 35077
rect 43533 35068 43545 35071
rect 43496 35040 43545 35068
rect 43496 35028 43502 35040
rect 43533 35037 43545 35040
rect 43579 35037 43591 35071
rect 43533 35031 43591 35037
rect 40221 35003 40279 35009
rect 39408 34972 39620 35000
rect 36538 34932 36544 34944
rect 35866 34904 36544 34932
rect 35621 34895 35679 34901
rect 36538 34892 36544 34904
rect 36596 34892 36602 34944
rect 37642 34892 37648 34944
rect 37700 34892 37706 34944
rect 39482 34892 39488 34944
rect 39540 34892 39546 34944
rect 39592 34932 39620 34972
rect 40221 34969 40233 35003
rect 40267 34969 40279 35003
rect 40221 34963 40279 34969
rect 40405 35003 40463 35009
rect 40405 34969 40417 35003
rect 40451 35000 40463 35003
rect 42058 35000 42064 35012
rect 40451 34972 42064 35000
rect 40451 34969 40463 34972
rect 40405 34963 40463 34969
rect 42058 34960 42064 34972
rect 42116 34960 42122 35012
rect 40021 34935 40079 34941
rect 40021 34932 40033 34935
rect 39592 34904 40033 34932
rect 40021 34901 40033 34904
rect 40067 34932 40079 34935
rect 42150 34932 42156 34944
rect 40067 34904 42156 34932
rect 40067 34901 40079 34904
rect 40021 34895 40079 34901
rect 42150 34892 42156 34904
rect 42208 34892 42214 34944
rect 43254 34892 43260 34944
rect 43312 34892 43318 34944
rect 43441 34935 43499 34941
rect 43441 34901 43453 34935
rect 43487 34932 43499 34935
rect 43714 34932 43720 34944
rect 43487 34904 43720 34932
rect 43487 34901 43499 34904
rect 43441 34895 43499 34901
rect 43714 34892 43720 34904
rect 43772 34892 43778 34944
rect 1104 34842 44620 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 44620 34842
rect 1104 34768 44620 34790
rect 5626 34688 5632 34740
rect 5684 34688 5690 34740
rect 5994 34728 6000 34740
rect 5828 34700 6000 34728
rect 5828 34669 5856 34700
rect 5994 34688 6000 34700
rect 6052 34688 6058 34740
rect 6086 34688 6092 34740
rect 6144 34728 6150 34740
rect 6457 34731 6515 34737
rect 6457 34728 6469 34731
rect 6144 34700 6469 34728
rect 6144 34688 6150 34700
rect 6457 34697 6469 34700
rect 6503 34728 6515 34731
rect 6638 34728 6644 34740
rect 6503 34700 6644 34728
rect 6503 34697 6515 34700
rect 6457 34691 6515 34697
rect 6638 34688 6644 34700
rect 6696 34688 6702 34740
rect 6730 34688 6736 34740
rect 6788 34688 6794 34740
rect 7466 34688 7472 34740
rect 7524 34688 7530 34740
rect 8294 34688 8300 34740
rect 8352 34688 8358 34740
rect 8662 34688 8668 34740
rect 8720 34688 8726 34740
rect 9398 34688 9404 34740
rect 9456 34688 9462 34740
rect 13446 34688 13452 34740
rect 13504 34688 13510 34740
rect 15654 34728 15660 34740
rect 14476 34700 15660 34728
rect 5813 34663 5871 34669
rect 5813 34629 5825 34663
rect 5859 34629 5871 34663
rect 6178 34660 6184 34672
rect 5813 34623 5871 34629
rect 5936 34632 6184 34660
rect 5936 34592 5964 34632
rect 6178 34620 6184 34632
rect 6236 34660 6242 34672
rect 6236 34632 6868 34660
rect 6236 34620 6242 34632
rect 5092 34564 5964 34592
rect 5997 34595 6055 34601
rect 5092 34536 5120 34564
rect 5997 34561 6009 34595
rect 6043 34592 6055 34595
rect 6362 34592 6368 34604
rect 6043 34564 6368 34592
rect 6043 34561 6055 34564
rect 5997 34555 6055 34561
rect 6362 34552 6368 34564
rect 6420 34552 6426 34604
rect 6454 34552 6460 34604
rect 6512 34592 6518 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6512 34564 6561 34592
rect 6512 34552 6518 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 6638 34552 6644 34604
rect 6696 34552 6702 34604
rect 6840 34601 6868 34632
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 7101 34595 7159 34601
rect 7101 34592 7113 34595
rect 6871 34564 7113 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 7101 34561 7113 34564
rect 7147 34561 7159 34595
rect 7101 34555 7159 34561
rect 7193 34595 7251 34601
rect 7193 34561 7205 34595
rect 7239 34592 7251 34595
rect 7484 34592 7512 34688
rect 8680 34660 8708 34688
rect 9416 34660 9444 34688
rect 11054 34660 11060 34672
rect 8128 34632 8708 34660
rect 8128 34601 8156 34632
rect 7239 34564 7512 34592
rect 8113 34595 8171 34601
rect 7239 34561 7251 34564
rect 7193 34555 7251 34561
rect 8113 34561 8125 34595
rect 8159 34561 8171 34595
rect 8113 34555 8171 34561
rect 8297 34595 8355 34601
rect 8297 34561 8309 34595
rect 8343 34592 8355 34595
rect 8389 34595 8447 34601
rect 8389 34592 8401 34595
rect 8343 34564 8401 34592
rect 8343 34561 8355 34564
rect 8297 34555 8355 34561
rect 8389 34561 8401 34564
rect 8435 34592 8447 34595
rect 8478 34592 8484 34604
rect 8435 34564 8484 34592
rect 8435 34561 8447 34564
rect 8389 34555 8447 34561
rect 8478 34552 8484 34564
rect 8536 34552 8542 34604
rect 8573 34595 8631 34601
rect 8573 34561 8585 34595
rect 8619 34592 8631 34595
rect 8680 34592 8708 34632
rect 9048 34632 9444 34660
rect 10534 34632 11060 34660
rect 8619 34564 8708 34592
rect 8619 34561 8631 34564
rect 8573 34555 8631 34561
rect 8846 34552 8852 34604
rect 8904 34552 8910 34604
rect 8938 34552 8944 34604
rect 8996 34552 9002 34604
rect 9048 34601 9076 34632
rect 11054 34620 11060 34632
rect 11112 34620 11118 34672
rect 12618 34660 12624 34672
rect 12452 34632 12624 34660
rect 9033 34595 9091 34601
rect 9033 34561 9045 34595
rect 9079 34561 9091 34595
rect 9033 34555 9091 34561
rect 11514 34552 11520 34604
rect 11572 34552 11578 34604
rect 12452 34601 12480 34632
rect 12618 34620 12624 34632
rect 12676 34660 12682 34672
rect 13464 34660 13492 34688
rect 12676 34632 13492 34660
rect 12676 34620 12682 34632
rect 12437 34595 12495 34601
rect 12437 34561 12449 34595
rect 12483 34561 12495 34595
rect 12437 34555 12495 34561
rect 12526 34552 12532 34604
rect 12584 34552 12590 34604
rect 12710 34552 12716 34604
rect 12768 34552 12774 34604
rect 12802 34552 12808 34604
rect 12860 34592 12866 34604
rect 12989 34595 13047 34601
rect 12989 34592 13001 34595
rect 12860 34564 13001 34592
rect 12860 34552 12866 34564
rect 12989 34561 13001 34564
rect 13035 34561 13047 34595
rect 12989 34555 13047 34561
rect 13078 34552 13084 34604
rect 13136 34592 13142 34604
rect 14476 34601 14504 34700
rect 15654 34688 15660 34700
rect 15712 34688 15718 34740
rect 16206 34688 16212 34740
rect 16264 34688 16270 34740
rect 16850 34688 16856 34740
rect 16908 34688 16914 34740
rect 17310 34688 17316 34740
rect 17368 34728 17374 34740
rect 17589 34731 17647 34737
rect 17589 34728 17601 34731
rect 17368 34700 17601 34728
rect 17368 34688 17374 34700
rect 17589 34697 17601 34700
rect 17635 34697 17647 34731
rect 18782 34728 18788 34740
rect 17589 34691 17647 34697
rect 18524 34700 18788 34728
rect 16482 34660 16488 34672
rect 15962 34632 16488 34660
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 16574 34620 16580 34672
rect 16632 34660 16638 34672
rect 16868 34660 16896 34688
rect 17497 34663 17555 34669
rect 16632 34632 17356 34660
rect 16632 34620 16638 34632
rect 13173 34595 13231 34601
rect 13173 34592 13185 34595
rect 13136 34564 13185 34592
rect 13136 34552 13142 34564
rect 13173 34561 13185 34564
rect 13219 34561 13231 34595
rect 13173 34555 13231 34561
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34561 14519 34595
rect 14461 34555 14519 34561
rect 17126 34552 17132 34604
rect 17184 34552 17190 34604
rect 17218 34552 17224 34604
rect 17276 34552 17282 34604
rect 17328 34601 17356 34632
rect 17497 34629 17509 34663
rect 17543 34660 17555 34663
rect 18524 34660 18552 34700
rect 18782 34688 18788 34700
rect 18840 34688 18846 34740
rect 18874 34688 18880 34740
rect 18932 34688 18938 34740
rect 19242 34688 19248 34740
rect 19300 34728 19306 34740
rect 19337 34731 19395 34737
rect 19337 34728 19349 34731
rect 19300 34700 19349 34728
rect 19300 34688 19306 34700
rect 19337 34697 19349 34700
rect 19383 34697 19395 34731
rect 25961 34731 26019 34737
rect 19337 34691 19395 34697
rect 22066 34700 24072 34728
rect 17543 34632 18552 34660
rect 17543 34629 17555 34632
rect 17497 34623 17555 34629
rect 18524 34601 18552 34632
rect 18693 34663 18751 34669
rect 18693 34629 18705 34663
rect 18739 34660 18751 34663
rect 19260 34660 19288 34688
rect 22066 34660 22094 34700
rect 23937 34663 23995 34669
rect 23937 34660 23949 34663
rect 18739 34632 19288 34660
rect 19352 34632 22094 34660
rect 23492 34632 23949 34660
rect 18739 34629 18751 34632
rect 18693 34623 18751 34629
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 18509 34595 18567 34601
rect 17313 34555 17371 34561
rect 17604 34564 18460 34592
rect 5074 34484 5080 34536
rect 5132 34484 5138 34536
rect 5442 34484 5448 34536
rect 5500 34524 5506 34536
rect 8662 34524 8668 34536
rect 5500 34496 8668 34524
rect 5500 34484 5506 34496
rect 8662 34484 8668 34496
rect 8720 34524 8726 34536
rect 8864 34524 8892 34552
rect 8720 34496 8892 34524
rect 12897 34527 12955 34533
rect 8720 34484 8726 34496
rect 12897 34493 12909 34527
rect 12943 34524 12955 34527
rect 13354 34524 13360 34536
rect 12943 34496 13360 34524
rect 12943 34493 12955 34496
rect 12897 34487 12955 34493
rect 13354 34484 13360 34496
rect 13412 34484 13418 34536
rect 14734 34484 14740 34536
rect 14792 34484 14798 34536
rect 17144 34524 17172 34552
rect 17604 34524 17632 34564
rect 17144 34496 17632 34524
rect 18046 34484 18052 34536
rect 18104 34484 18110 34536
rect 18233 34527 18291 34533
rect 18233 34493 18245 34527
rect 18279 34524 18291 34527
rect 18325 34527 18383 34533
rect 18325 34524 18337 34527
rect 18279 34496 18337 34524
rect 18279 34493 18291 34496
rect 18233 34487 18291 34493
rect 18325 34493 18337 34496
rect 18371 34493 18383 34527
rect 18432 34524 18460 34564
rect 18509 34561 18521 34595
rect 18555 34561 18567 34595
rect 18509 34555 18567 34561
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18800 34524 18828 34555
rect 19242 34552 19248 34604
rect 19300 34552 19306 34604
rect 19352 34524 19380 34632
rect 18432 34496 19380 34524
rect 19429 34527 19487 34533
rect 18325 34487 18383 34493
rect 19429 34493 19441 34527
rect 19475 34493 19487 34527
rect 19429 34487 19487 34493
rect 8573 34459 8631 34465
rect 8573 34425 8585 34459
rect 8619 34456 8631 34459
rect 8846 34456 8852 34468
rect 8619 34428 8852 34456
rect 8619 34425 8631 34428
rect 8573 34419 8631 34425
rect 8846 34416 8852 34428
rect 8904 34416 8910 34468
rect 18064 34456 18092 34484
rect 19058 34456 19064 34468
rect 18064 34428 19064 34456
rect 19058 34416 19064 34428
rect 19116 34456 19122 34468
rect 19444 34456 19472 34487
rect 22002 34484 22008 34536
rect 22060 34524 22066 34536
rect 22833 34527 22891 34533
rect 22833 34524 22845 34527
rect 22060 34496 22845 34524
rect 22060 34484 22066 34496
rect 22833 34493 22845 34496
rect 22879 34493 22891 34527
rect 22833 34487 22891 34493
rect 22554 34456 22560 34468
rect 19116 34428 22560 34456
rect 19116 34416 19122 34428
rect 22554 34416 22560 34428
rect 22612 34416 22618 34468
rect 23492 34400 23520 34632
rect 23937 34629 23949 34632
rect 23983 34629 23995 34663
rect 23937 34623 23995 34629
rect 24044 34604 24072 34700
rect 25961 34697 25973 34731
rect 26007 34728 26019 34731
rect 26050 34728 26056 34740
rect 26007 34700 26056 34728
rect 26007 34697 26019 34700
rect 25961 34691 26019 34697
rect 26050 34688 26056 34700
rect 26108 34688 26114 34740
rect 27890 34688 27896 34740
rect 27948 34688 27954 34740
rect 30190 34688 30196 34740
rect 30248 34728 30254 34740
rect 33502 34728 33508 34740
rect 30248 34700 33508 34728
rect 30248 34688 30254 34700
rect 33502 34688 33508 34700
rect 33560 34688 33566 34740
rect 35621 34731 35679 34737
rect 35268 34700 35572 34728
rect 24486 34620 24492 34672
rect 24544 34620 24550 34672
rect 25222 34620 25228 34672
rect 25280 34620 25286 34672
rect 27433 34663 27491 34669
rect 27433 34629 27445 34663
rect 27479 34660 27491 34663
rect 27801 34663 27859 34669
rect 27801 34660 27813 34663
rect 27479 34632 27813 34660
rect 27479 34629 27491 34632
rect 27433 34623 27491 34629
rect 27801 34629 27813 34632
rect 27847 34629 27859 34663
rect 27908 34660 27936 34688
rect 28442 34660 28448 34672
rect 27908 34632 28448 34660
rect 27801 34623 27859 34629
rect 28442 34620 28448 34632
rect 28500 34660 28506 34672
rect 34606 34660 34612 34672
rect 28500 34632 28764 34660
rect 28500 34620 28506 34632
rect 23566 34552 23572 34604
rect 23624 34552 23630 34604
rect 23658 34552 23664 34604
rect 23716 34592 23722 34604
rect 23753 34595 23811 34601
rect 23753 34592 23765 34595
rect 23716 34564 23765 34592
rect 23716 34552 23722 34564
rect 23753 34561 23765 34564
rect 23799 34561 23811 34595
rect 23753 34555 23811 34561
rect 24026 34552 24032 34604
rect 24084 34552 24090 34604
rect 27246 34552 27252 34604
rect 27304 34552 27310 34604
rect 27522 34552 27528 34604
rect 27580 34552 27586 34604
rect 28736 34601 28764 34632
rect 28828 34632 34612 34660
rect 27893 34595 27951 34601
rect 27893 34561 27905 34595
rect 27939 34592 27951 34595
rect 28169 34595 28227 34601
rect 28169 34592 28181 34595
rect 27939 34564 28181 34592
rect 27939 34561 27951 34564
rect 27893 34555 27951 34561
rect 28169 34561 28181 34564
rect 28215 34561 28227 34595
rect 28169 34555 28227 34561
rect 28721 34595 28779 34601
rect 28721 34561 28733 34595
rect 28767 34561 28779 34595
rect 28721 34555 28779 34561
rect 23584 34524 23612 34552
rect 24213 34527 24271 34533
rect 24213 34524 24225 34527
rect 23584 34496 24225 34524
rect 24213 34493 24225 34496
rect 24259 34493 24271 34527
rect 24213 34487 24271 34493
rect 26786 34484 26792 34536
rect 26844 34524 26850 34536
rect 28828 34524 28856 34632
rect 34606 34620 34612 34632
rect 34664 34620 34670 34672
rect 35268 34669 35296 34700
rect 35253 34663 35311 34669
rect 35253 34629 35265 34663
rect 35299 34629 35311 34663
rect 35253 34623 35311 34629
rect 35342 34620 35348 34672
rect 35400 34620 35406 34672
rect 35544 34660 35572 34700
rect 35621 34697 35633 34731
rect 35667 34728 35679 34731
rect 36078 34728 36084 34740
rect 35667 34700 36084 34728
rect 35667 34697 35679 34700
rect 35621 34691 35679 34697
rect 36078 34688 36084 34700
rect 36136 34688 36142 34740
rect 37642 34728 37648 34740
rect 36464 34700 37648 34728
rect 36170 34660 36176 34672
rect 35544 34632 36176 34660
rect 36170 34620 36176 34632
rect 36228 34620 36234 34672
rect 36464 34669 36492 34700
rect 37642 34688 37648 34700
rect 37700 34688 37706 34740
rect 37918 34688 37924 34740
rect 37976 34728 37982 34740
rect 38013 34731 38071 34737
rect 38013 34728 38025 34731
rect 37976 34700 38025 34728
rect 37976 34688 37982 34700
rect 38013 34697 38025 34700
rect 38059 34697 38071 34731
rect 38013 34691 38071 34697
rect 39114 34688 39120 34740
rect 39172 34728 39178 34740
rect 40221 34731 40279 34737
rect 40221 34728 40233 34731
rect 39172 34700 40233 34728
rect 39172 34688 39178 34700
rect 40221 34697 40233 34700
rect 40267 34697 40279 34731
rect 42058 34728 42064 34740
rect 40221 34691 40279 34697
rect 41892 34700 42064 34728
rect 36449 34663 36507 34669
rect 36449 34629 36461 34663
rect 36495 34629 36507 34663
rect 36449 34623 36507 34629
rect 36538 34620 36544 34672
rect 36596 34660 36602 34672
rect 41892 34669 41920 34700
rect 42058 34688 42064 34700
rect 42116 34688 42122 34740
rect 42242 34688 42248 34740
rect 42300 34688 42306 34740
rect 42521 34731 42579 34737
rect 42521 34697 42533 34731
rect 42567 34728 42579 34731
rect 42702 34728 42708 34740
rect 42567 34700 42708 34728
rect 42567 34697 42579 34700
rect 42521 34691 42579 34697
rect 36649 34663 36707 34669
rect 36649 34660 36661 34663
rect 36596 34632 36661 34660
rect 36596 34620 36602 34632
rect 36649 34629 36661 34632
rect 36695 34629 36707 34663
rect 36649 34623 36707 34629
rect 41877 34663 41935 34669
rect 41877 34629 41889 34663
rect 41923 34629 41935 34663
rect 41877 34623 41935 34629
rect 42107 34629 42165 34635
rect 42107 34626 42119 34629
rect 30742 34552 30748 34604
rect 30800 34552 30806 34604
rect 30926 34552 30932 34604
rect 30984 34552 30990 34604
rect 35069 34595 35127 34601
rect 35069 34561 35081 34595
rect 35115 34561 35127 34595
rect 35069 34555 35127 34561
rect 26844 34496 28856 34524
rect 30837 34527 30895 34533
rect 26844 34484 26850 34496
rect 30837 34493 30849 34527
rect 30883 34524 30895 34527
rect 32306 34524 32312 34536
rect 30883 34496 32312 34524
rect 30883 34493 30895 34496
rect 30837 34487 30895 34493
rect 32306 34484 32312 34496
rect 32364 34484 32370 34536
rect 35084 34524 35112 34555
rect 35434 34552 35440 34604
rect 35492 34552 35498 34604
rect 36188 34592 36216 34620
rect 37461 34595 37519 34601
rect 36188 34564 36584 34592
rect 36556 34536 36584 34564
rect 37461 34561 37473 34595
rect 37507 34561 37519 34595
rect 37921 34595 37979 34601
rect 37921 34592 37933 34595
rect 37461 34555 37519 34561
rect 37568 34564 37933 34592
rect 35342 34524 35348 34536
rect 35084 34496 35348 34524
rect 35342 34484 35348 34496
rect 35400 34484 35406 34536
rect 35802 34484 35808 34536
rect 35860 34524 35866 34536
rect 36262 34524 36268 34536
rect 35860 34496 36268 34524
rect 35860 34484 35866 34496
rect 36262 34484 36268 34496
rect 36320 34484 36326 34536
rect 36538 34484 36544 34536
rect 36596 34484 36602 34536
rect 31018 34456 31024 34468
rect 26896 34428 31024 34456
rect 26896 34400 26924 34428
rect 31018 34416 31024 34428
rect 31076 34456 31082 34468
rect 37476 34456 37504 34555
rect 31076 34428 37504 34456
rect 31076 34416 31082 34428
rect 8757 34391 8815 34397
rect 8757 34357 8769 34391
rect 8803 34388 8815 34391
rect 9030 34388 9036 34400
rect 8803 34360 9036 34388
rect 8803 34357 8815 34360
rect 8757 34351 8815 34357
rect 9030 34348 9036 34360
rect 9088 34348 9094 34400
rect 9306 34397 9312 34400
rect 9296 34391 9312 34397
rect 9296 34357 9308 34391
rect 9296 34351 9312 34357
rect 9306 34348 9312 34351
rect 9364 34348 9370 34400
rect 10778 34348 10784 34400
rect 10836 34348 10842 34400
rect 11606 34348 11612 34400
rect 11664 34348 11670 34400
rect 12986 34348 12992 34400
rect 13044 34348 13050 34400
rect 23474 34348 23480 34400
rect 23532 34348 23538 34400
rect 23566 34348 23572 34400
rect 23624 34348 23630 34400
rect 26878 34348 26884 34400
rect 26936 34348 26942 34400
rect 27062 34348 27068 34400
rect 27120 34388 27126 34400
rect 27249 34391 27307 34397
rect 27249 34388 27261 34391
rect 27120 34360 27261 34388
rect 27120 34348 27126 34360
rect 27249 34357 27261 34360
rect 27295 34357 27307 34391
rect 27249 34351 27307 34357
rect 36262 34348 36268 34400
rect 36320 34388 36326 34400
rect 36633 34391 36691 34397
rect 36633 34388 36645 34391
rect 36320 34360 36645 34388
rect 36320 34348 36326 34360
rect 36633 34357 36645 34360
rect 36679 34357 36691 34391
rect 36633 34351 36691 34357
rect 36817 34391 36875 34397
rect 36817 34357 36829 34391
rect 36863 34388 36875 34391
rect 37568 34388 37596 34564
rect 37921 34561 37933 34564
rect 37967 34561 37979 34595
rect 37921 34555 37979 34561
rect 38010 34552 38016 34604
rect 38068 34592 38074 34604
rect 38378 34592 38384 34604
rect 38068 34564 38384 34592
rect 38068 34552 38074 34564
rect 38378 34552 38384 34564
rect 38436 34552 38442 34604
rect 39482 34552 39488 34604
rect 39540 34592 39546 34604
rect 40773 34595 40831 34601
rect 40773 34592 40785 34595
rect 39540 34564 40785 34592
rect 39540 34552 39546 34564
rect 40773 34561 40785 34564
rect 40819 34561 40831 34595
rect 40773 34555 40831 34561
rect 41414 34552 41420 34604
rect 41472 34592 41478 34604
rect 42092 34595 42119 34626
rect 42153 34604 42165 34629
rect 42153 34595 42156 34604
rect 42092 34592 42156 34595
rect 41472 34564 42156 34592
rect 41472 34552 41478 34564
rect 42150 34552 42156 34564
rect 42208 34552 42214 34604
rect 42536 34456 42564 34691
rect 42702 34688 42708 34700
rect 42760 34688 42766 34740
rect 42610 34620 42616 34672
rect 42668 34660 42674 34672
rect 42668 34632 42826 34660
rect 42668 34620 42674 34632
rect 43714 34620 43720 34672
rect 43772 34660 43778 34672
rect 43993 34663 44051 34669
rect 43993 34660 44005 34663
rect 43772 34632 44005 34660
rect 43772 34620 43778 34632
rect 43993 34629 44005 34632
rect 44039 34629 44051 34663
rect 43993 34623 44051 34629
rect 44266 34552 44272 34604
rect 44324 34552 44330 34604
rect 42076 34428 42564 34456
rect 36863 34360 37596 34388
rect 36863 34357 36875 34360
rect 36817 34351 36875 34357
rect 37642 34348 37648 34400
rect 37700 34348 37706 34400
rect 38470 34348 38476 34400
rect 38528 34388 38534 34400
rect 39390 34388 39396 34400
rect 38528 34360 39396 34388
rect 38528 34348 38534 34360
rect 39390 34348 39396 34360
rect 39448 34388 39454 34400
rect 42076 34397 42104 34428
rect 39669 34391 39727 34397
rect 39669 34388 39681 34391
rect 39448 34360 39681 34388
rect 39448 34348 39454 34360
rect 39669 34357 39681 34360
rect 39715 34357 39727 34391
rect 39669 34351 39727 34357
rect 42061 34391 42119 34397
rect 42061 34357 42073 34391
rect 42107 34357 42119 34391
rect 42061 34351 42119 34357
rect 1104 34298 44620 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 44620 34298
rect 1104 34224 44620 34246
rect 5534 34144 5540 34196
rect 5592 34184 5598 34196
rect 6181 34187 6239 34193
rect 6181 34184 6193 34187
rect 5592 34156 6193 34184
rect 5592 34144 5598 34156
rect 6181 34153 6193 34156
rect 6227 34153 6239 34187
rect 6181 34147 6239 34153
rect 9217 34187 9275 34193
rect 9217 34153 9229 34187
rect 9263 34184 9275 34187
rect 9306 34184 9312 34196
rect 9263 34156 9312 34184
rect 9263 34153 9275 34156
rect 9217 34147 9275 34153
rect 9306 34144 9312 34156
rect 9364 34144 9370 34196
rect 12345 34187 12403 34193
rect 12345 34153 12357 34187
rect 12391 34184 12403 34187
rect 12710 34184 12716 34196
rect 12391 34156 12716 34184
rect 12391 34153 12403 34156
rect 12345 34147 12403 34153
rect 12710 34144 12716 34156
rect 12768 34144 12774 34196
rect 12894 34144 12900 34196
rect 12952 34184 12958 34196
rect 14277 34187 14335 34193
rect 14277 34184 14289 34187
rect 12952 34156 14289 34184
rect 12952 34144 12958 34156
rect 6086 34076 6092 34128
rect 6144 34076 6150 34128
rect 12618 34076 12624 34128
rect 12676 34076 12682 34128
rect 13372 34125 13400 34156
rect 14277 34153 14289 34156
rect 14323 34153 14335 34187
rect 14277 34147 14335 34153
rect 14734 34144 14740 34196
rect 14792 34144 14798 34196
rect 15654 34144 15660 34196
rect 15712 34184 15718 34196
rect 15933 34187 15991 34193
rect 15933 34184 15945 34187
rect 15712 34156 15945 34184
rect 15712 34144 15718 34156
rect 15933 34153 15945 34156
rect 15979 34153 15991 34187
rect 15933 34147 15991 34153
rect 17773 34187 17831 34193
rect 17773 34153 17785 34187
rect 17819 34184 17831 34187
rect 17954 34184 17960 34196
rect 17819 34156 17960 34184
rect 17819 34153 17831 34156
rect 17773 34147 17831 34153
rect 17954 34144 17960 34156
rect 18012 34184 18018 34196
rect 21542 34184 21548 34196
rect 18012 34156 21548 34184
rect 18012 34144 18018 34156
rect 21542 34144 21548 34156
rect 21600 34144 21606 34196
rect 25038 34144 25044 34196
rect 25096 34144 25102 34196
rect 28442 34144 28448 34196
rect 28500 34144 28506 34196
rect 30377 34187 30435 34193
rect 30377 34153 30389 34187
rect 30423 34184 30435 34187
rect 30742 34184 30748 34196
rect 30423 34156 30748 34184
rect 30423 34153 30435 34156
rect 30377 34147 30435 34153
rect 30742 34144 30748 34156
rect 30800 34144 30806 34196
rect 30926 34144 30932 34196
rect 30984 34184 30990 34196
rect 31110 34184 31116 34196
rect 30984 34156 31116 34184
rect 30984 34144 30990 34156
rect 31110 34144 31116 34156
rect 31168 34144 31174 34196
rect 31386 34144 31392 34196
rect 31444 34144 31450 34196
rect 32858 34144 32864 34196
rect 32916 34144 32922 34196
rect 33318 34144 33324 34196
rect 33376 34184 33382 34196
rect 33778 34184 33784 34196
rect 33376 34156 33784 34184
rect 33376 34144 33382 34156
rect 33778 34144 33784 34156
rect 33836 34144 33842 34196
rect 34054 34144 34060 34196
rect 34112 34144 34118 34196
rect 35161 34187 35219 34193
rect 35161 34153 35173 34187
rect 35207 34184 35219 34187
rect 35342 34184 35348 34196
rect 35207 34156 35348 34184
rect 35207 34153 35219 34156
rect 35161 34147 35219 34153
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 39482 34144 39488 34196
rect 39540 34184 39546 34196
rect 39577 34187 39635 34193
rect 39577 34184 39589 34187
rect 39540 34156 39589 34184
rect 39540 34144 39546 34156
rect 39577 34153 39589 34156
rect 39623 34153 39635 34187
rect 39577 34147 39635 34153
rect 42981 34187 43039 34193
rect 42981 34153 42993 34187
rect 43027 34184 43039 34187
rect 43438 34184 43444 34196
rect 43027 34156 43444 34184
rect 43027 34153 43039 34156
rect 42981 34147 43039 34153
rect 43438 34144 43444 34156
rect 43496 34144 43502 34196
rect 13265 34119 13323 34125
rect 13265 34116 13277 34119
rect 12728 34088 13277 34116
rect 6104 34048 6132 34076
rect 10597 34051 10655 34057
rect 6104 34020 6316 34048
rect 5721 33983 5779 33989
rect 5721 33949 5733 33983
rect 5767 33949 5779 33983
rect 5721 33943 5779 33949
rect 6089 33983 6147 33989
rect 6089 33949 6101 33983
rect 6135 33980 6147 33983
rect 6178 33980 6184 33992
rect 6135 33952 6184 33980
rect 6135 33949 6147 33952
rect 6089 33943 6147 33949
rect 5736 33912 5764 33943
rect 6178 33940 6184 33952
rect 6236 33940 6242 33992
rect 6288 33989 6316 34020
rect 10597 34017 10609 34051
rect 10643 34048 10655 34051
rect 10778 34048 10784 34060
rect 10643 34020 10784 34048
rect 10643 34017 10655 34020
rect 10597 34011 10655 34017
rect 10778 34008 10784 34020
rect 10836 34048 10842 34060
rect 11330 34048 11336 34060
rect 10836 34020 11336 34048
rect 10836 34008 10842 34020
rect 11330 34008 11336 34020
rect 11388 34008 11394 34060
rect 12342 34048 12348 34060
rect 11532 34020 12348 34048
rect 6273 33983 6331 33989
rect 6273 33949 6285 33983
rect 6319 33949 6331 33983
rect 6273 33943 6331 33949
rect 6362 33940 6368 33992
rect 6420 33940 6426 33992
rect 8846 33940 8852 33992
rect 8904 33980 8910 33992
rect 8941 33983 8999 33989
rect 8941 33980 8953 33983
rect 8904 33952 8953 33980
rect 8904 33940 8910 33952
rect 8941 33949 8953 33952
rect 8987 33949 8999 33983
rect 8941 33943 8999 33949
rect 9030 33940 9036 33992
rect 9088 33980 9094 33992
rect 11532 33989 11560 34020
rect 12342 34008 12348 34020
rect 12400 34008 12406 34060
rect 9217 33983 9275 33989
rect 9217 33980 9229 33983
rect 9088 33952 9229 33980
rect 9088 33940 9094 33952
rect 9217 33949 9229 33952
rect 9263 33949 9275 33983
rect 9217 33943 9275 33949
rect 11425 33983 11483 33989
rect 11425 33949 11437 33983
rect 11471 33949 11483 33983
rect 11425 33943 11483 33949
rect 11517 33983 11575 33989
rect 11517 33949 11529 33983
rect 11563 33949 11575 33983
rect 11517 33943 11575 33949
rect 6380 33912 6408 33940
rect 5736 33884 6408 33912
rect 5534 33804 5540 33856
rect 5592 33844 5598 33856
rect 5629 33847 5687 33853
rect 5629 33844 5641 33847
rect 5592 33816 5641 33844
rect 5592 33804 5598 33816
rect 5629 33813 5641 33816
rect 5675 33813 5687 33847
rect 5629 33807 5687 33813
rect 8938 33804 8944 33856
rect 8996 33844 9002 33856
rect 9033 33847 9091 33853
rect 9033 33844 9045 33847
rect 8996 33816 9045 33844
rect 8996 33804 9002 33816
rect 9033 33813 9045 33816
rect 9079 33844 9091 33847
rect 9953 33847 10011 33853
rect 9953 33844 9965 33847
rect 9079 33816 9965 33844
rect 9079 33813 9091 33816
rect 9033 33807 9091 33813
rect 9953 33813 9965 33816
rect 9999 33813 10011 33847
rect 11440 33844 11468 33943
rect 11606 33940 11612 33992
rect 11664 33940 11670 33992
rect 11701 33983 11759 33989
rect 11701 33949 11713 33983
rect 11747 33980 11759 33983
rect 11790 33980 11796 33992
rect 11747 33952 11796 33980
rect 11747 33949 11759 33952
rect 11701 33943 11759 33949
rect 11790 33940 11796 33952
rect 11848 33940 11854 33992
rect 12066 33940 12072 33992
rect 12124 33980 12130 33992
rect 12250 33980 12256 33992
rect 12124 33952 12256 33980
rect 12124 33940 12130 33952
rect 12250 33940 12256 33952
rect 12308 33940 12314 33992
rect 12526 33940 12532 33992
rect 12584 33940 12590 33992
rect 12636 33989 12664 34076
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33949 12679 33983
rect 12621 33943 12679 33949
rect 11624 33912 11652 33940
rect 11885 33915 11943 33921
rect 11885 33912 11897 33915
rect 11624 33884 11897 33912
rect 11885 33881 11897 33884
rect 11931 33881 11943 33915
rect 11885 33875 11943 33881
rect 11974 33872 11980 33924
rect 12032 33872 12038 33924
rect 12728 33912 12756 34088
rect 13265 34085 13277 34088
rect 13311 34085 13323 34119
rect 13265 34079 13323 34085
rect 13357 34119 13415 34125
rect 13357 34085 13369 34119
rect 13403 34085 13415 34119
rect 13357 34079 13415 34085
rect 13633 34119 13691 34125
rect 13633 34085 13645 34119
rect 13679 34116 13691 34119
rect 19334 34116 19340 34128
rect 13679 34088 19340 34116
rect 13679 34085 13691 34088
rect 13633 34079 13691 34085
rect 19334 34076 19340 34088
rect 19392 34076 19398 34128
rect 20806 34076 20812 34128
rect 20864 34116 20870 34128
rect 22278 34116 22284 34128
rect 20864 34088 22284 34116
rect 20864 34076 20870 34088
rect 22278 34076 22284 34088
rect 22336 34076 22342 34128
rect 25133 34119 25191 34125
rect 25133 34116 25145 34119
rect 24688 34088 25145 34116
rect 24688 34060 24716 34088
rect 25133 34085 25145 34088
rect 25179 34085 25191 34119
rect 25133 34079 25191 34085
rect 30558 34076 30564 34128
rect 30616 34076 30622 34128
rect 31018 34076 31024 34128
rect 31076 34076 31082 34128
rect 12986 34008 12992 34060
rect 13044 34048 13050 34060
rect 20898 34048 20904 34060
rect 13044 34020 13952 34048
rect 13044 34008 13050 34020
rect 13170 33940 13176 33992
rect 13228 33940 13234 33992
rect 13446 33940 13452 33992
rect 13504 33940 13510 33992
rect 13924 33989 13952 34020
rect 14108 34020 14504 34048
rect 14108 33989 14136 34020
rect 14476 33992 14504 34020
rect 20272 34020 20904 34048
rect 13725 33983 13783 33989
rect 13725 33979 13737 33983
rect 13648 33951 13737 33979
rect 12176 33884 12756 33912
rect 12176 33856 12204 33884
rect 12802 33872 12808 33924
rect 12860 33912 12866 33924
rect 12897 33915 12955 33921
rect 12897 33912 12909 33915
rect 12860 33884 12909 33912
rect 12860 33872 12866 33884
rect 12897 33881 12909 33884
rect 12943 33881 12955 33915
rect 12897 33875 12955 33881
rect 12989 33915 13047 33921
rect 12989 33881 13001 33915
rect 13035 33912 13047 33915
rect 13078 33912 13084 33924
rect 13035 33884 13084 33912
rect 13035 33881 13047 33884
rect 12989 33875 13047 33881
rect 13078 33872 13084 33884
rect 13136 33872 13142 33924
rect 11790 33844 11796 33856
rect 11440 33816 11796 33844
rect 9953 33807 10011 33813
rect 11790 33804 11796 33816
rect 11848 33804 11854 33856
rect 12158 33804 12164 33856
rect 12216 33804 12222 33856
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 12434 33804 12440 33856
rect 12492 33844 12498 33856
rect 13648 33844 13676 33951
rect 13725 33949 13737 33951
rect 13771 33949 13783 33983
rect 13725 33943 13783 33949
rect 13909 33983 13967 33989
rect 13909 33949 13921 33983
rect 13955 33949 13967 33983
rect 13909 33943 13967 33949
rect 14093 33983 14151 33989
rect 14093 33949 14105 33983
rect 14139 33949 14151 33983
rect 14093 33943 14151 33949
rect 14182 33940 14188 33992
rect 14240 33980 14246 33992
rect 14277 33983 14335 33989
rect 14277 33980 14289 33983
rect 14240 33952 14289 33980
rect 14240 33940 14246 33952
rect 14277 33949 14289 33952
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 14458 33940 14464 33992
rect 14516 33940 14522 33992
rect 14918 33940 14924 33992
rect 14976 33940 14982 33992
rect 15838 33940 15844 33992
rect 15896 33980 15902 33992
rect 20272 33989 20300 34020
rect 20898 34008 20904 34020
rect 20956 34008 20962 34060
rect 22554 34008 22560 34060
rect 22612 34008 22618 34060
rect 22649 34051 22707 34057
rect 22649 34017 22661 34051
rect 22695 34048 22707 34051
rect 23474 34048 23480 34060
rect 22695 34020 23480 34048
rect 22695 34017 22707 34020
rect 22649 34011 22707 34017
rect 23474 34008 23480 34020
rect 23532 34008 23538 34060
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 23937 34051 23995 34057
rect 23937 34048 23949 34051
rect 23624 34020 23949 34048
rect 23624 34008 23630 34020
rect 23937 34017 23949 34020
rect 23983 34017 23995 34051
rect 23937 34011 23995 34017
rect 24670 34008 24676 34060
rect 24728 34008 24734 34060
rect 24762 34008 24768 34060
rect 24820 34048 24826 34060
rect 25685 34051 25743 34057
rect 25685 34048 25697 34051
rect 24820 34020 25697 34048
rect 24820 34008 24826 34020
rect 25685 34017 25697 34020
rect 25731 34017 25743 34051
rect 25685 34011 25743 34017
rect 26973 34051 27031 34057
rect 26973 34017 26985 34051
rect 27019 34048 27031 34051
rect 27062 34048 27068 34060
rect 27019 34020 27068 34048
rect 27019 34017 27031 34020
rect 26973 34011 27031 34017
rect 27062 34008 27068 34020
rect 27120 34008 27126 34060
rect 17405 33983 17463 33989
rect 17405 33980 17417 33983
rect 15896 33952 17417 33980
rect 15896 33940 15902 33952
rect 17405 33949 17417 33952
rect 17451 33980 17463 33983
rect 20257 33983 20315 33989
rect 17451 33952 19196 33980
rect 17451 33949 17463 33952
rect 17405 33943 17463 33949
rect 19168 33924 19196 33952
rect 20257 33949 20269 33983
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 21450 33980 21456 33992
rect 20487 33952 21456 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 24394 33940 24400 33992
rect 24452 33940 24458 33992
rect 24545 33983 24603 33989
rect 24545 33949 24557 33983
rect 24591 33980 24603 33983
rect 24688 33980 24716 34008
rect 24591 33952 24716 33980
rect 24591 33949 24603 33952
rect 24545 33943 24603 33949
rect 24854 33940 24860 33992
rect 24912 33989 24918 33992
rect 24912 33980 24920 33989
rect 24912 33952 24957 33980
rect 24912 33943 24920 33952
rect 24912 33940 24918 33943
rect 26050 33940 26056 33992
rect 26108 33940 26114 33992
rect 26602 33940 26608 33992
rect 26660 33980 26666 33992
rect 26697 33983 26755 33989
rect 26697 33980 26709 33983
rect 26660 33952 26709 33980
rect 26660 33940 26666 33952
rect 26697 33949 26709 33952
rect 26743 33949 26755 33983
rect 26697 33943 26755 33949
rect 30193 33983 30251 33989
rect 30193 33949 30205 33983
rect 30239 33980 30251 33983
rect 30576 33980 30604 34076
rect 31036 34048 31064 34076
rect 31404 34048 31432 34144
rect 37274 34116 37280 34128
rect 33704 34088 37280 34116
rect 31036 34020 31156 34048
rect 31021 33983 31079 33989
rect 31021 33980 31033 33983
rect 30239 33952 31033 33980
rect 30239 33949 30251 33952
rect 30193 33943 30251 33949
rect 31021 33949 31033 33952
rect 31067 33949 31079 33983
rect 31021 33943 31079 33949
rect 17586 33872 17592 33924
rect 17644 33912 17650 33924
rect 17865 33915 17923 33921
rect 17865 33912 17877 33915
rect 17644 33884 17877 33912
rect 17644 33872 17650 33884
rect 17865 33881 17877 33884
rect 17911 33881 17923 33915
rect 17865 33875 17923 33881
rect 19150 33872 19156 33924
rect 19208 33912 19214 33924
rect 23014 33912 23020 33924
rect 19208 33884 23020 33912
rect 19208 33872 19214 33884
rect 23014 33872 23020 33884
rect 23072 33872 23078 33924
rect 23566 33912 23572 33924
rect 23124 33884 23572 33912
rect 12492 33816 13676 33844
rect 12492 33804 12498 33816
rect 13814 33804 13820 33856
rect 13872 33804 13878 33856
rect 20346 33804 20352 33856
rect 20404 33804 20410 33856
rect 22738 33804 22744 33856
rect 22796 33804 22802 33856
rect 23124 33853 23152 33884
rect 23566 33872 23572 33884
rect 23624 33872 23630 33924
rect 24673 33915 24731 33921
rect 24673 33912 24685 33915
rect 24596 33884 24685 33912
rect 24596 33856 24624 33884
rect 24673 33881 24685 33884
rect 24719 33881 24731 33915
rect 24673 33875 24731 33881
rect 24765 33915 24823 33921
rect 24765 33881 24777 33915
rect 24811 33912 24823 33915
rect 26068 33912 26096 33940
rect 24811 33884 26096 33912
rect 24811 33881 24823 33884
rect 24765 33875 24823 33881
rect 26418 33872 26424 33924
rect 26476 33912 26482 33924
rect 27430 33912 27436 33924
rect 26476 33884 27436 33912
rect 26476 33872 26482 33884
rect 27430 33872 27436 33884
rect 27488 33872 27494 33924
rect 30009 33915 30067 33921
rect 30009 33881 30021 33915
rect 30055 33912 30067 33915
rect 30837 33915 30895 33921
rect 30055 33884 30788 33912
rect 30055 33881 30067 33884
rect 30009 33875 30067 33881
rect 23109 33847 23167 33853
rect 23109 33813 23121 33847
rect 23155 33813 23167 33847
rect 23109 33807 23167 33813
rect 23382 33804 23388 33856
rect 23440 33804 23446 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 29822 33804 29828 33856
rect 29880 33844 29886 33856
rect 30561 33847 30619 33853
rect 30561 33844 30573 33847
rect 29880 33816 30573 33844
rect 29880 33804 29886 33816
rect 30561 33813 30573 33816
rect 30607 33813 30619 33847
rect 30760 33844 30788 33884
rect 30837 33881 30849 33915
rect 30883 33912 30895 33915
rect 31128 33912 31156 34020
rect 31220 34020 31432 34048
rect 31220 33989 31248 34020
rect 33502 34008 33508 34060
rect 33560 34048 33566 34060
rect 33597 34051 33655 34057
rect 33597 34048 33609 34051
rect 33560 34020 33609 34048
rect 33560 34008 33566 34020
rect 33597 34017 33609 34020
rect 33643 34017 33655 34051
rect 33597 34011 33655 34017
rect 33704 33992 33732 34088
rect 37274 34076 37280 34088
rect 37332 34116 37338 34128
rect 37332 34088 37504 34116
rect 37332 34076 37338 34088
rect 34149 34051 34207 34057
rect 34149 34048 34161 34051
rect 33980 34020 34161 34048
rect 31205 33983 31263 33989
rect 31205 33949 31217 33983
rect 31251 33949 31263 33983
rect 31205 33943 31263 33949
rect 30883 33884 31156 33912
rect 30883 33881 30895 33884
rect 30837 33875 30895 33881
rect 31220 33856 31248 33943
rect 31386 33940 31392 33992
rect 31444 33940 31450 33992
rect 32306 33940 32312 33992
rect 32364 33940 32370 33992
rect 32490 33940 32496 33992
rect 32548 33940 32554 33992
rect 32582 33940 32588 33992
rect 32640 33940 32646 33992
rect 33686 33940 33692 33992
rect 33744 33940 33750 33992
rect 32766 33872 32772 33924
rect 32824 33872 32830 33924
rect 33980 33912 34008 34020
rect 34149 34017 34161 34020
rect 34195 34017 34207 34051
rect 34149 34011 34207 34017
rect 34790 34008 34796 34060
rect 34848 34008 34854 34060
rect 37476 34057 37504 34088
rect 37461 34051 37519 34057
rect 37461 34017 37473 34051
rect 37507 34017 37519 34051
rect 37461 34011 37519 34017
rect 37829 34051 37887 34057
rect 37829 34017 37841 34051
rect 37875 34048 37887 34051
rect 38470 34048 38476 34060
rect 37875 34020 38476 34048
rect 37875 34017 37887 34020
rect 37829 34011 37887 34017
rect 38470 34008 38476 34020
rect 38528 34008 38534 34060
rect 40862 34048 40868 34060
rect 40512 34020 40868 34048
rect 34057 33983 34115 33989
rect 34057 33949 34069 33983
rect 34103 33949 34115 33983
rect 34057 33943 34115 33949
rect 34885 33983 34943 33989
rect 34885 33949 34897 33983
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 33060 33884 34008 33912
rect 34072 33912 34100 33943
rect 34900 33912 34928 33943
rect 39850 33940 39856 33992
rect 39908 33980 39914 33992
rect 40512 33989 40540 34020
rect 40862 34008 40868 34020
rect 40920 34048 40926 34060
rect 40957 34051 41015 34057
rect 40957 34048 40969 34051
rect 40920 34020 40969 34048
rect 40920 34008 40926 34020
rect 40957 34017 40969 34020
rect 41003 34017 41015 34051
rect 40957 34011 41015 34017
rect 41414 34008 41420 34060
rect 41472 34008 41478 34060
rect 41877 34051 41935 34057
rect 41877 34017 41889 34051
rect 41923 34048 41935 34051
rect 41923 34020 43944 34048
rect 41923 34017 41935 34020
rect 41877 34011 41935 34017
rect 40313 33983 40371 33989
rect 40313 33980 40325 33983
rect 39908 33952 40325 33980
rect 39908 33940 39914 33952
rect 40313 33949 40325 33952
rect 40359 33949 40371 33983
rect 40313 33943 40371 33949
rect 40497 33983 40555 33989
rect 40497 33949 40509 33983
rect 40543 33949 40555 33983
rect 40497 33943 40555 33949
rect 40773 33983 40831 33989
rect 40773 33949 40785 33983
rect 40819 33949 40831 33983
rect 41432 33980 41460 34008
rect 40773 33943 40831 33949
rect 41386 33952 41460 33980
rect 41509 33983 41567 33989
rect 34072 33884 34928 33912
rect 38105 33915 38163 33921
rect 33060 33856 33088 33884
rect 31202 33844 31208 33856
rect 30760 33816 31208 33844
rect 30561 33807 30619 33813
rect 31202 33804 31208 33816
rect 31260 33804 31266 33856
rect 32030 33804 32036 33856
rect 32088 33804 32094 33856
rect 32122 33804 32128 33856
rect 32180 33804 32186 33856
rect 33042 33804 33048 33856
rect 33100 33804 33106 33856
rect 33226 33804 33232 33856
rect 33284 33844 33290 33856
rect 33321 33847 33379 33853
rect 33321 33844 33333 33847
rect 33284 33816 33333 33844
rect 33284 33804 33290 33816
rect 33321 33813 33333 33816
rect 33367 33844 33379 33847
rect 34072 33844 34100 33884
rect 38105 33881 38117 33915
rect 38151 33881 38163 33915
rect 40328 33912 40356 33943
rect 40788 33912 40816 33943
rect 39330 33884 39804 33912
rect 40328 33884 40816 33912
rect 38105 33875 38163 33881
rect 33367 33816 34100 33844
rect 33367 33813 33379 33816
rect 33321 33807 33379 33813
rect 34422 33804 34428 33856
rect 34480 33804 34486 33856
rect 36906 33804 36912 33856
rect 36964 33804 36970 33856
rect 38120 33844 38148 33875
rect 39776 33856 39804 33884
rect 38746 33844 38752 33856
rect 38120 33816 38752 33844
rect 38746 33804 38752 33816
rect 38804 33804 38810 33856
rect 39758 33804 39764 33856
rect 39816 33804 39822 33856
rect 40402 33804 40408 33856
rect 40460 33804 40466 33856
rect 40586 33804 40592 33856
rect 40644 33844 40650 33856
rect 41386 33844 41414 33952
rect 41509 33949 41521 33983
rect 41555 33949 41567 33983
rect 41509 33943 41567 33949
rect 41524 33912 41552 33943
rect 42058 33940 42064 33992
rect 42116 33940 42122 33992
rect 42150 33940 42156 33992
rect 42208 33980 42214 33992
rect 42705 33983 42763 33989
rect 42705 33980 42717 33983
rect 42208 33952 42717 33980
rect 42208 33940 42214 33952
rect 42705 33949 42717 33952
rect 42751 33949 42763 33983
rect 42705 33943 42763 33949
rect 42981 33983 43039 33989
rect 42981 33949 42993 33983
rect 43027 33980 43039 33983
rect 43254 33980 43260 33992
rect 43027 33952 43260 33980
rect 43027 33949 43039 33952
rect 42981 33943 43039 33949
rect 43254 33940 43260 33952
rect 43312 33940 43318 33992
rect 42613 33915 42671 33921
rect 42613 33912 42625 33915
rect 41524 33884 42625 33912
rect 42613 33881 42625 33884
rect 42659 33912 42671 33915
rect 42797 33915 42855 33921
rect 42797 33912 42809 33915
rect 42659 33884 42809 33912
rect 42659 33881 42671 33884
rect 42613 33875 42671 33881
rect 42797 33881 42809 33884
rect 42843 33881 42855 33915
rect 42797 33875 42855 33881
rect 43916 33856 43944 34020
rect 44634 34008 44640 34060
rect 44692 34008 44698 34060
rect 44269 33983 44327 33989
rect 44269 33949 44281 33983
rect 44315 33980 44327 33983
rect 44652 33980 44680 34008
rect 44315 33952 44680 33980
rect 44315 33949 44327 33952
rect 44269 33943 44327 33949
rect 40644 33816 41414 33844
rect 40644 33804 40650 33816
rect 43898 33804 43904 33856
rect 43956 33804 43962 33856
rect 44082 33804 44088 33856
rect 44140 33804 44146 33856
rect 1104 33754 44620 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 44620 33754
rect 1104 33680 44620 33702
rect 6362 33600 6368 33652
rect 6420 33600 6426 33652
rect 8386 33600 8392 33652
rect 8444 33600 8450 33652
rect 11974 33600 11980 33652
rect 12032 33600 12038 33652
rect 12161 33643 12219 33649
rect 12161 33609 12173 33643
rect 12207 33640 12219 33643
rect 12710 33640 12716 33652
rect 12207 33612 12716 33640
rect 12207 33609 12219 33612
rect 12161 33603 12219 33609
rect 12710 33600 12716 33612
rect 12768 33600 12774 33652
rect 13814 33640 13820 33652
rect 12820 33612 13820 33640
rect 5166 33464 5172 33516
rect 5224 33504 5230 33516
rect 5997 33507 6055 33513
rect 5224 33476 5290 33504
rect 5224 33464 5230 33476
rect 5997 33473 6009 33507
rect 6043 33473 6055 33507
rect 5997 33467 6055 33473
rect 6181 33507 6239 33513
rect 6181 33473 6193 33507
rect 6227 33504 6239 33507
rect 6549 33507 6607 33513
rect 6549 33504 6561 33507
rect 6227 33476 6561 33504
rect 6227 33473 6239 33476
rect 6181 33467 6239 33473
rect 6549 33473 6561 33476
rect 6595 33504 6607 33507
rect 8404 33504 8432 33600
rect 11992 33572 12020 33600
rect 12820 33572 12848 33612
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 14829 33643 14887 33649
rect 14829 33609 14841 33643
rect 14875 33640 14887 33643
rect 14918 33640 14924 33652
rect 14875 33612 14924 33640
rect 14875 33609 14887 33612
rect 14829 33603 14887 33609
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 15197 33643 15255 33649
rect 15197 33609 15209 33643
rect 15243 33640 15255 33643
rect 15746 33640 15752 33652
rect 15243 33612 15752 33640
rect 15243 33609 15255 33612
rect 15197 33603 15255 33609
rect 15746 33600 15752 33612
rect 15804 33600 15810 33652
rect 20254 33600 20260 33652
rect 20312 33600 20318 33652
rect 20714 33600 20720 33652
rect 20772 33640 20778 33652
rect 21082 33640 21088 33652
rect 20772 33612 21088 33640
rect 20772 33600 20778 33612
rect 21082 33600 21088 33612
rect 21140 33600 21146 33652
rect 22002 33600 22008 33652
rect 22060 33600 22066 33652
rect 25038 33640 25044 33652
rect 22204 33612 25044 33640
rect 11808 33544 12020 33572
rect 12084 33544 12848 33572
rect 14737 33575 14795 33581
rect 9309 33507 9367 33513
rect 9309 33504 9321 33507
rect 6595 33476 8064 33504
rect 8404 33476 9321 33504
rect 6595 33473 6607 33476
rect 6549 33467 6607 33473
rect 3878 33396 3884 33448
rect 3936 33396 3942 33448
rect 4157 33439 4215 33445
rect 4157 33405 4169 33439
rect 4203 33436 4215 33439
rect 4614 33436 4620 33448
rect 4203 33408 4620 33436
rect 4203 33405 4215 33408
rect 4157 33399 4215 33405
rect 4614 33396 4620 33408
rect 4672 33396 4678 33448
rect 5629 33439 5687 33445
rect 5629 33405 5641 33439
rect 5675 33436 5687 33439
rect 6012 33436 6040 33467
rect 8036 33448 8064 33476
rect 9309 33473 9321 33476
rect 9355 33473 9367 33507
rect 9309 33467 9367 33473
rect 11606 33464 11612 33516
rect 11664 33504 11670 33516
rect 11808 33513 11836 33544
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 11664 33476 11805 33504
rect 11664 33464 11670 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 11882 33464 11888 33516
rect 11940 33464 11946 33516
rect 11974 33464 11980 33516
rect 12032 33464 12038 33516
rect 12084 33513 12112 33544
rect 14737 33541 14749 33575
rect 14783 33572 14795 33575
rect 22204 33572 22232 33612
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 26234 33640 26240 33652
rect 25792 33612 26240 33640
rect 14783 33544 22232 33572
rect 14783 33541 14795 33544
rect 14737 33535 14795 33541
rect 23382 33532 23388 33584
rect 23440 33572 23446 33584
rect 23477 33575 23535 33581
rect 23477 33572 23489 33575
rect 23440 33544 23489 33572
rect 23440 33532 23446 33544
rect 23477 33541 23489 33544
rect 23523 33541 23535 33575
rect 23477 33535 23535 33541
rect 23566 33532 23572 33584
rect 23624 33572 23630 33584
rect 25792 33572 25820 33612
rect 26234 33600 26240 33612
rect 26292 33640 26298 33652
rect 26418 33640 26424 33652
rect 26292 33612 26424 33640
rect 26292 33600 26298 33612
rect 26418 33600 26424 33612
rect 26476 33600 26482 33652
rect 27890 33640 27896 33652
rect 27264 33612 27896 33640
rect 23624 33544 24072 33572
rect 25622 33544 25820 33572
rect 26053 33575 26111 33581
rect 23624 33532 23630 33544
rect 12069 33507 12127 33513
rect 12069 33473 12081 33507
rect 12115 33473 12127 33507
rect 12069 33467 12127 33473
rect 12250 33464 12256 33516
rect 12308 33504 12314 33516
rect 12345 33507 12403 33513
rect 12345 33504 12357 33507
rect 12308 33476 12357 33504
rect 12308 33464 12314 33476
rect 12345 33473 12357 33476
rect 12391 33473 12403 33507
rect 12345 33467 12403 33473
rect 12437 33507 12495 33513
rect 12437 33473 12449 33507
rect 12483 33504 12495 33507
rect 12618 33504 12624 33516
rect 12483 33476 12624 33504
rect 12483 33473 12495 33476
rect 12437 33467 12495 33473
rect 12618 33464 12624 33476
rect 12676 33464 12682 33516
rect 12713 33507 12771 33513
rect 12713 33473 12725 33507
rect 12759 33504 12771 33507
rect 12986 33504 12992 33516
rect 12759 33476 12992 33504
rect 12759 33473 12771 33476
rect 12713 33467 12771 33473
rect 12986 33464 12992 33476
rect 13044 33464 13050 33516
rect 15838 33504 15844 33516
rect 15212 33476 15844 33504
rect 6733 33439 6791 33445
rect 6733 33436 6745 33439
rect 5675 33408 6745 33436
rect 5675 33405 5687 33408
rect 5629 33399 5687 33405
rect 6733 33405 6745 33408
rect 6779 33405 6791 33439
rect 6733 33399 6791 33405
rect 6748 33368 6776 33399
rect 8018 33396 8024 33448
rect 8076 33396 8082 33448
rect 11900 33436 11928 33464
rect 12529 33439 12587 33445
rect 12529 33436 12541 33439
rect 11900 33408 12541 33436
rect 12529 33405 12541 33408
rect 12575 33405 12587 33439
rect 12529 33399 12587 33405
rect 9766 33368 9772 33380
rect 6748 33340 9772 33368
rect 9766 33328 9772 33340
rect 9824 33328 9830 33380
rect 12158 33328 12164 33380
rect 12216 33368 12222 33380
rect 12345 33371 12403 33377
rect 12345 33368 12357 33371
rect 12216 33340 12357 33368
rect 12216 33328 12222 33340
rect 12345 33337 12357 33340
rect 12391 33337 12403 33371
rect 12345 33331 12403 33337
rect 12434 33328 12440 33380
rect 12492 33368 12498 33380
rect 12492 33340 12572 33368
rect 12492 33328 12498 33340
rect 5810 33260 5816 33312
rect 5868 33260 5874 33312
rect 9401 33303 9459 33309
rect 9401 33269 9413 33303
rect 9447 33300 9459 33303
rect 12066 33300 12072 33312
rect 9447 33272 12072 33300
rect 9447 33269 9459 33272
rect 9401 33263 9459 33269
rect 12066 33260 12072 33272
rect 12124 33260 12130 33312
rect 12544 33309 12572 33340
rect 13262 33328 13268 33380
rect 13320 33368 13326 33380
rect 13449 33371 13507 33377
rect 13449 33368 13461 33371
rect 13320 33340 13461 33368
rect 13320 33328 13326 33340
rect 13449 33337 13461 33340
rect 13495 33368 13507 33371
rect 15212 33368 15240 33476
rect 15838 33464 15844 33476
rect 15896 33464 15902 33516
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 17037 33507 17095 33513
rect 16071 33476 16712 33504
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 15289 33439 15347 33445
rect 15289 33405 15301 33439
rect 15335 33405 15347 33439
rect 15289 33399 15347 33405
rect 15473 33439 15531 33445
rect 15473 33405 15485 33439
rect 15519 33436 15531 33439
rect 15519 33408 16620 33436
rect 15519 33405 15531 33408
rect 15473 33399 15531 33405
rect 13495 33340 15240 33368
rect 15304 33368 15332 33399
rect 16022 33368 16028 33380
rect 15304 33340 16028 33368
rect 13495 33337 13507 33340
rect 13449 33331 13507 33337
rect 16022 33328 16028 33340
rect 16080 33328 16086 33380
rect 12529 33303 12587 33309
rect 12529 33269 12541 33303
rect 12575 33269 12587 33303
rect 12529 33263 12587 33269
rect 12894 33260 12900 33312
rect 12952 33260 12958 33312
rect 13170 33260 13176 33312
rect 13228 33300 13234 33312
rect 13814 33300 13820 33312
rect 13228 33272 13820 33300
rect 13228 33260 13234 33272
rect 13814 33260 13820 33272
rect 13872 33260 13878 33312
rect 15841 33303 15899 33309
rect 15841 33269 15853 33303
rect 15887 33300 15899 33303
rect 15930 33300 15936 33312
rect 15887 33272 15936 33300
rect 15887 33269 15899 33272
rect 15841 33263 15899 33269
rect 15930 33260 15936 33272
rect 15988 33260 15994 33312
rect 16592 33300 16620 33408
rect 16684 33377 16712 33476
rect 17037 33473 17049 33507
rect 17083 33504 17095 33507
rect 17497 33507 17555 33513
rect 17497 33504 17509 33507
rect 17083 33476 17509 33504
rect 17083 33473 17095 33476
rect 17037 33467 17095 33473
rect 17497 33473 17509 33476
rect 17543 33473 17555 33507
rect 17497 33467 17555 33473
rect 18414 33464 18420 33516
rect 18472 33464 18478 33516
rect 18877 33507 18935 33513
rect 18877 33504 18889 33507
rect 18524 33476 18889 33504
rect 18524 33448 18552 33476
rect 18877 33473 18889 33476
rect 18923 33473 18935 33507
rect 18877 33467 18935 33473
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33473 19303 33507
rect 19245 33467 19303 33473
rect 17126 33396 17132 33448
rect 17184 33396 17190 33448
rect 17221 33439 17279 33445
rect 17221 33405 17233 33439
rect 17267 33436 17279 33439
rect 17310 33436 17316 33448
rect 17267 33408 17316 33436
rect 17267 33405 17279 33408
rect 17221 33399 17279 33405
rect 16669 33371 16727 33377
rect 16669 33337 16681 33371
rect 16715 33337 16727 33371
rect 17236 33368 17264 33399
rect 17310 33396 17316 33408
rect 17368 33396 17374 33448
rect 18049 33439 18107 33445
rect 18049 33405 18061 33439
rect 18095 33405 18107 33439
rect 18049 33399 18107 33405
rect 16669 33331 16727 33337
rect 17144 33340 17264 33368
rect 17144 33300 17172 33340
rect 16592 33272 17172 33300
rect 17218 33260 17224 33312
rect 17276 33300 17282 33312
rect 18064 33300 18092 33399
rect 18506 33396 18512 33448
rect 18564 33396 18570 33448
rect 19260 33436 19288 33467
rect 19334 33464 19340 33516
rect 19392 33464 19398 33516
rect 19426 33464 19432 33516
rect 19484 33464 19490 33516
rect 19705 33507 19763 33513
rect 19705 33473 19717 33507
rect 19751 33504 19763 33507
rect 19751 33476 20116 33504
rect 19751 33473 19763 33476
rect 19705 33467 19763 33473
rect 19444 33436 19472 33464
rect 19260 33408 19472 33436
rect 19260 33368 19288 33408
rect 20088 33377 20116 33476
rect 20162 33464 20168 33516
rect 20220 33504 20226 33516
rect 20254 33507 20312 33513
rect 20254 33504 20266 33507
rect 20220 33476 20266 33504
rect 20220 33464 20226 33476
rect 20254 33473 20266 33476
rect 20300 33504 20312 33507
rect 21085 33507 21143 33513
rect 20300 33476 20852 33504
rect 20300 33473 20312 33476
rect 20254 33467 20312 33473
rect 20622 33436 20628 33448
rect 20180 33408 20628 33436
rect 18616 33340 19288 33368
rect 20073 33371 20131 33377
rect 18616 33309 18644 33340
rect 20073 33337 20085 33371
rect 20119 33337 20131 33371
rect 20073 33331 20131 33337
rect 17276 33272 18092 33300
rect 18601 33303 18659 33309
rect 17276 33260 17282 33272
rect 18601 33269 18613 33303
rect 18647 33269 18659 33303
rect 18601 33263 18659 33269
rect 18785 33303 18843 33309
rect 18785 33269 18797 33303
rect 18831 33300 18843 33303
rect 19518 33300 19524 33312
rect 18831 33272 19524 33300
rect 18831 33269 18843 33272
rect 18785 33263 18843 33269
rect 19518 33260 19524 33272
rect 19576 33260 19582 33312
rect 19705 33303 19763 33309
rect 19705 33269 19717 33303
rect 19751 33300 19763 33303
rect 20180 33300 20208 33408
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 20717 33439 20775 33445
rect 20717 33405 20729 33439
rect 20763 33405 20775 33439
rect 20717 33399 20775 33405
rect 19751 33272 20208 33300
rect 19751 33269 19763 33272
rect 19705 33263 19763 33269
rect 20622 33260 20628 33312
rect 20680 33260 20686 33312
rect 20732 33300 20760 33399
rect 20824 33377 20852 33476
rect 21085 33473 21097 33507
rect 21131 33504 21143 33507
rect 21266 33504 21272 33516
rect 21131 33476 21272 33504
rect 21131 33473 21143 33476
rect 21085 33467 21143 33473
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 21450 33464 21456 33516
rect 21508 33464 21514 33516
rect 21542 33464 21548 33516
rect 21600 33504 21606 33516
rect 24044 33513 24072 33544
rect 26053 33541 26065 33575
rect 26099 33572 26111 33575
rect 26510 33572 26516 33584
rect 26099 33544 26516 33572
rect 26099 33541 26111 33544
rect 26053 33535 26111 33541
rect 26510 33532 26516 33544
rect 26568 33532 26574 33584
rect 27264 33581 27292 33612
rect 27890 33600 27896 33612
rect 27948 33600 27954 33652
rect 28534 33600 28540 33652
rect 28592 33640 28598 33652
rect 28721 33643 28779 33649
rect 28721 33640 28733 33643
rect 28592 33612 28733 33640
rect 28592 33600 28598 33612
rect 28721 33609 28733 33612
rect 28767 33609 28779 33643
rect 28721 33603 28779 33609
rect 31021 33643 31079 33649
rect 31021 33609 31033 33643
rect 31067 33640 31079 33643
rect 31386 33640 31392 33652
rect 31067 33612 31392 33640
rect 31067 33609 31079 33612
rect 31021 33603 31079 33609
rect 31386 33600 31392 33612
rect 31444 33600 31450 33652
rect 32030 33600 32036 33652
rect 32088 33600 32094 33652
rect 32306 33649 32312 33652
rect 32293 33643 32312 33649
rect 32293 33609 32305 33643
rect 32293 33603 32312 33609
rect 32306 33600 32312 33603
rect 32364 33600 32370 33652
rect 33410 33600 33416 33652
rect 33468 33640 33474 33652
rect 33468 33612 33640 33640
rect 33468 33600 33474 33612
rect 27249 33575 27307 33581
rect 27249 33541 27261 33575
rect 27295 33541 27307 33575
rect 27249 33535 27307 33541
rect 27522 33532 27528 33584
rect 27580 33572 27586 33584
rect 29822 33572 29828 33584
rect 27580 33544 27738 33572
rect 29012 33544 29828 33572
rect 27580 33532 27586 33544
rect 29012 33516 29040 33544
rect 29822 33532 29828 33544
rect 29880 33572 29886 33584
rect 31757 33575 31815 33581
rect 29880 33544 30038 33572
rect 29880 33532 29886 33544
rect 31757 33541 31769 33575
rect 31803 33572 31815 33575
rect 32048 33572 32076 33600
rect 31803 33544 32076 33572
rect 31803 33541 31815 33544
rect 31757 33535 31815 33541
rect 32122 33532 32128 33584
rect 32180 33532 32186 33584
rect 32490 33532 32496 33584
rect 32548 33532 32554 33584
rect 33612 33581 33640 33612
rect 33686 33600 33692 33652
rect 33744 33600 33750 33652
rect 33965 33643 34023 33649
rect 33965 33609 33977 33643
rect 34011 33609 34023 33643
rect 33965 33603 34023 33609
rect 33137 33575 33195 33581
rect 33137 33541 33149 33575
rect 33183 33572 33195 33575
rect 33597 33575 33655 33581
rect 33183 33544 33456 33572
rect 33183 33541 33195 33544
rect 33137 33535 33195 33541
rect 24029 33507 24087 33513
rect 21600 33476 22402 33504
rect 21600 33464 21606 33476
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 26697 33507 26755 33513
rect 26697 33473 26709 33507
rect 26743 33504 26755 33507
rect 26878 33504 26884 33516
rect 26743 33476 26884 33504
rect 26743 33473 26755 33476
rect 26697 33467 26755 33473
rect 26878 33464 26884 33476
rect 26936 33464 26942 33516
rect 28994 33464 29000 33516
rect 29052 33464 29058 33516
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33504 31447 33507
rect 32140 33504 32168 33532
rect 32585 33507 32643 33513
rect 32585 33504 32597 33507
rect 31435 33476 31984 33504
rect 32140 33476 32597 33504
rect 31435 33473 31447 33476
rect 31389 33467 31447 33473
rect 20898 33396 20904 33448
rect 20956 33396 20962 33448
rect 20990 33396 20996 33448
rect 21048 33396 21054 33448
rect 21361 33439 21419 33445
rect 21361 33405 21373 33439
rect 21407 33405 21419 33439
rect 21361 33399 21419 33405
rect 23753 33439 23811 33445
rect 23753 33405 23765 33439
rect 23799 33436 23811 33439
rect 26329 33439 26387 33445
rect 23799 33408 25084 33436
rect 23799 33405 23811 33408
rect 23753 33399 23811 33405
rect 20809 33371 20867 33377
rect 20809 33337 20821 33371
rect 20855 33337 20867 33371
rect 20916 33368 20944 33396
rect 21376 33368 21404 33399
rect 20916 33340 21404 33368
rect 24581 33371 24639 33377
rect 20809 33331 20867 33337
rect 24581 33337 24593 33371
rect 24627 33368 24639 33371
rect 24762 33368 24768 33380
rect 24627 33340 24768 33368
rect 24627 33337 24639 33340
rect 24581 33331 24639 33337
rect 24762 33328 24768 33340
rect 24820 33328 24826 33380
rect 21174 33300 21180 33312
rect 20732 33272 21180 33300
rect 21174 33260 21180 33272
rect 21232 33260 21238 33312
rect 23842 33260 23848 33312
rect 23900 33260 23906 33312
rect 25056 33300 25084 33408
rect 26329 33405 26341 33439
rect 26375 33436 26387 33439
rect 26602 33436 26608 33448
rect 26375 33408 26608 33436
rect 26375 33405 26387 33408
rect 26329 33399 26387 33405
rect 26344 33300 26372 33399
rect 26602 33396 26608 33408
rect 26660 33436 26666 33448
rect 26973 33439 27031 33445
rect 26973 33436 26985 33439
rect 26660 33408 26985 33436
rect 26660 33396 26666 33408
rect 26973 33405 26985 33408
rect 27019 33436 27031 33439
rect 28626 33436 28632 33448
rect 27019 33408 28632 33436
rect 27019 33405 27031 33408
rect 26973 33399 27031 33405
rect 28626 33396 28632 33408
rect 28684 33436 28690 33448
rect 29273 33439 29331 33445
rect 29273 33436 29285 33439
rect 28684 33408 29285 33436
rect 28684 33396 28690 33408
rect 29273 33405 29285 33408
rect 29319 33405 29331 33439
rect 29273 33399 29331 33405
rect 29549 33439 29607 33445
rect 29549 33405 29561 33439
rect 29595 33436 29607 33439
rect 31297 33439 31355 33445
rect 29595 33408 31156 33436
rect 29595 33405 29607 33408
rect 29549 33399 29607 33405
rect 26418 33328 26424 33380
rect 26476 33328 26482 33380
rect 31128 33377 31156 33408
rect 31297 33405 31309 33439
rect 31343 33405 31355 33439
rect 31297 33399 31355 33405
rect 31113 33371 31171 33377
rect 31113 33337 31125 33371
rect 31159 33337 31171 33371
rect 31312 33368 31340 33399
rect 31570 33396 31576 33448
rect 31628 33436 31634 33448
rect 31665 33439 31723 33445
rect 31665 33436 31677 33439
rect 31628 33408 31677 33436
rect 31628 33396 31634 33408
rect 31665 33405 31677 33408
rect 31711 33405 31723 33439
rect 31956 33436 31984 33476
rect 32585 33473 32597 33476
rect 32631 33473 32643 33507
rect 32585 33467 32643 33473
rect 32766 33464 32772 33516
rect 32824 33464 32830 33516
rect 33042 33464 33048 33516
rect 33100 33464 33106 33516
rect 33226 33464 33232 33516
rect 33284 33464 33290 33516
rect 33318 33464 33324 33516
rect 33376 33464 33382 33516
rect 33428 33513 33456 33544
rect 33597 33541 33609 33575
rect 33643 33541 33655 33575
rect 33597 33535 33655 33541
rect 33704 33513 33732 33600
rect 33414 33507 33472 33513
rect 33414 33473 33426 33507
rect 33460 33473 33472 33507
rect 33414 33467 33472 33473
rect 33689 33507 33747 33513
rect 33689 33473 33701 33507
rect 33735 33473 33747 33507
rect 33689 33467 33747 33473
rect 33778 33464 33784 33516
rect 33836 33513 33842 33516
rect 33836 33504 33844 33513
rect 33980 33504 34008 33603
rect 34422 33600 34428 33652
rect 34480 33600 34486 33652
rect 34514 33600 34520 33652
rect 34572 33600 34578 33652
rect 36538 33640 36544 33652
rect 36372 33612 36544 33640
rect 34241 33507 34299 33513
rect 34241 33504 34253 33507
rect 33836 33476 33881 33504
rect 33980 33476 34253 33504
rect 33836 33467 33844 33476
rect 34241 33473 34253 33476
rect 34287 33473 34299 33507
rect 34440 33504 34468 33600
rect 34532 33572 34560 33600
rect 36372 33581 36400 33612
rect 36538 33600 36544 33612
rect 36596 33600 36602 33652
rect 36906 33600 36912 33652
rect 36964 33600 36970 33652
rect 37274 33600 37280 33652
rect 37332 33600 37338 33652
rect 39758 33600 39764 33652
rect 39816 33600 39822 33652
rect 40862 33600 40868 33652
rect 40920 33640 40926 33652
rect 41049 33643 41107 33649
rect 41049 33640 41061 33643
rect 40920 33612 41061 33640
rect 40920 33600 40926 33612
rect 41049 33609 41061 33612
rect 41095 33609 41107 33643
rect 41049 33603 41107 33609
rect 42058 33600 42064 33652
rect 42116 33640 42122 33652
rect 42429 33643 42487 33649
rect 42429 33640 42441 33643
rect 42116 33612 42441 33640
rect 42116 33600 42122 33612
rect 42429 33609 42441 33612
rect 42475 33609 42487 33643
rect 42429 33603 42487 33609
rect 42536 33612 43576 33640
rect 36357 33575 36415 33581
rect 34532 33544 34744 33572
rect 34716 33513 34744 33544
rect 35452 33544 36308 33572
rect 35452 33516 35480 33544
rect 34517 33507 34575 33513
rect 34517 33504 34529 33507
rect 34440 33476 34529 33504
rect 34241 33467 34299 33473
rect 34517 33473 34529 33476
rect 34563 33473 34575 33507
rect 34517 33467 34575 33473
rect 34701 33507 34759 33513
rect 34701 33473 34713 33507
rect 34747 33473 34759 33507
rect 35161 33507 35219 33513
rect 35161 33504 35173 33507
rect 34701 33467 34759 33473
rect 34808 33476 35173 33504
rect 33836 33464 33842 33467
rect 32677 33439 32735 33445
rect 32677 33436 32689 33439
rect 31956 33408 32689 33436
rect 31665 33399 31723 33405
rect 32677 33405 32689 33408
rect 32723 33405 32735 33439
rect 32677 33399 32735 33405
rect 32125 33371 32183 33377
rect 32125 33368 32137 33371
rect 31312 33340 32137 33368
rect 31113 33331 31171 33337
rect 32125 33337 32137 33340
rect 32171 33337 32183 33371
rect 32784 33368 32812 33464
rect 33060 33436 33088 33464
rect 34808 33436 34836 33476
rect 35161 33473 35173 33476
rect 35207 33504 35219 33507
rect 35342 33504 35348 33516
rect 35207 33476 35348 33504
rect 35207 33473 35219 33476
rect 35161 33467 35219 33473
rect 35342 33464 35348 33476
rect 35400 33464 35406 33516
rect 35434 33464 35440 33516
rect 35492 33464 35498 33516
rect 36173 33507 36231 33513
rect 36173 33504 36185 33507
rect 35866 33476 36185 33504
rect 33060 33408 34836 33436
rect 35069 33439 35127 33445
rect 35069 33405 35081 33439
rect 35115 33405 35127 33439
rect 35069 33399 35127 33405
rect 35529 33439 35587 33445
rect 35529 33405 35541 33439
rect 35575 33436 35587 33439
rect 35866 33436 35894 33476
rect 36173 33473 36185 33476
rect 36219 33473 36231 33507
rect 36280 33504 36308 33544
rect 36357 33541 36369 33575
rect 36403 33541 36415 33575
rect 36357 33535 36415 33541
rect 36449 33575 36507 33581
rect 36449 33541 36461 33575
rect 36495 33572 36507 33575
rect 36924 33572 36952 33600
rect 36495 33544 36952 33572
rect 36495 33541 36507 33544
rect 36449 33535 36507 33541
rect 38286 33532 38292 33584
rect 38344 33572 38350 33584
rect 39776 33572 39804 33600
rect 42536 33572 42564 33612
rect 38344 33544 39804 33572
rect 40802 33558 42564 33572
rect 40788 33544 42564 33558
rect 38344 33532 38350 33544
rect 36541 33507 36599 33513
rect 36541 33504 36553 33507
rect 36280 33476 36553 33504
rect 36173 33467 36231 33473
rect 36541 33473 36553 33476
rect 36587 33504 36599 33507
rect 36814 33504 36820 33516
rect 36587 33476 36820 33504
rect 36587 33473 36599 33476
rect 36541 33467 36599 33473
rect 36814 33464 36820 33476
rect 36872 33464 36878 33516
rect 38749 33439 38807 33445
rect 38749 33436 38761 33439
rect 35575 33408 35894 33436
rect 36740 33408 38761 33436
rect 35575 33405 35587 33408
rect 35529 33399 35587 33405
rect 32784 33340 33088 33368
rect 32125 33331 32183 33337
rect 25056 33272 26372 33300
rect 26436 33300 26464 33328
rect 33060 33312 33088 33340
rect 33870 33328 33876 33380
rect 33928 33368 33934 33380
rect 34057 33371 34115 33377
rect 34057 33368 34069 33371
rect 33928 33340 34069 33368
rect 33928 33328 33934 33340
rect 34057 33337 34069 33340
rect 34103 33337 34115 33371
rect 34057 33331 34115 33337
rect 34698 33328 34704 33380
rect 34756 33368 34762 33380
rect 35084 33368 35112 33399
rect 36740 33377 36768 33408
rect 38749 33405 38761 33408
rect 38795 33405 38807 33439
rect 38749 33399 38807 33405
rect 39025 33439 39083 33445
rect 39025 33405 39037 33439
rect 39071 33436 39083 33439
rect 39301 33439 39359 33445
rect 39301 33436 39313 33439
rect 39071 33408 39313 33436
rect 39071 33405 39083 33408
rect 39025 33399 39083 33405
rect 39301 33405 39313 33408
rect 39347 33405 39359 33439
rect 39301 33399 39359 33405
rect 39577 33439 39635 33445
rect 39577 33405 39589 33439
rect 39623 33436 39635 33439
rect 40126 33436 40132 33448
rect 39623 33408 40132 33436
rect 39623 33405 39635 33408
rect 39577 33399 39635 33405
rect 34756 33340 35112 33368
rect 36725 33371 36783 33377
rect 34756 33328 34762 33340
rect 36725 33337 36737 33371
rect 36771 33337 36783 33371
rect 36725 33331 36783 33337
rect 26513 33303 26571 33309
rect 26513 33300 26525 33303
rect 26436 33272 26525 33300
rect 26513 33269 26525 33272
rect 26559 33269 26571 33303
rect 26513 33263 26571 33269
rect 32309 33303 32367 33309
rect 32309 33269 32321 33303
rect 32355 33300 32367 33303
rect 32582 33300 32588 33312
rect 32355 33272 32588 33300
rect 32355 33269 32367 33272
rect 32309 33263 32367 33269
rect 32582 33260 32588 33272
rect 32640 33260 32646 33312
rect 33042 33260 33048 33312
rect 33100 33260 33106 33312
rect 38378 33260 38384 33312
rect 38436 33300 38442 33312
rect 39040 33300 39068 33399
rect 40126 33396 40132 33408
rect 40184 33396 40190 33448
rect 38436 33272 39068 33300
rect 38436 33260 38442 33272
rect 39758 33260 39764 33312
rect 39816 33300 39822 33312
rect 40788 33300 40816 33544
rect 43438 33532 43444 33584
rect 43496 33572 43502 33584
rect 43548 33572 43576 33612
rect 43496 33544 43576 33572
rect 43496 33532 43502 33544
rect 43898 33532 43904 33584
rect 43956 33532 43962 33584
rect 44177 33439 44235 33445
rect 44177 33405 44189 33439
rect 44223 33405 44235 33439
rect 44177 33399 44235 33405
rect 39816 33272 40816 33300
rect 39816 33260 39822 33272
rect 42518 33260 42524 33312
rect 42576 33300 42582 33312
rect 44192 33300 44220 33399
rect 42576 33272 44220 33300
rect 42576 33260 42582 33272
rect 1104 33210 44620 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 44620 33210
rect 1104 33136 44620 33158
rect 4614 33056 4620 33108
rect 4672 33056 4678 33108
rect 5445 33099 5503 33105
rect 5445 33065 5457 33099
rect 5491 33096 5503 33099
rect 5810 33096 5816 33108
rect 5491 33068 5816 33096
rect 5491 33065 5503 33068
rect 5445 33059 5503 33065
rect 5810 33056 5816 33068
rect 5868 33056 5874 33108
rect 8294 33056 8300 33108
rect 8352 33096 8358 33108
rect 8665 33099 8723 33105
rect 8665 33096 8677 33099
rect 8352 33068 8677 33096
rect 8352 33056 8358 33068
rect 8665 33065 8677 33068
rect 8711 33096 8723 33099
rect 9122 33096 9128 33108
rect 8711 33068 9128 33096
rect 8711 33065 8723 33068
rect 8665 33059 8723 33065
rect 9122 33056 9128 33068
rect 9180 33056 9186 33108
rect 12066 33056 12072 33108
rect 12124 33096 12130 33108
rect 12618 33096 12624 33108
rect 12124 33068 12624 33096
rect 12124 33056 12130 33068
rect 12618 33056 12624 33068
rect 12676 33056 12682 33108
rect 13449 33099 13507 33105
rect 13449 33065 13461 33099
rect 13495 33096 13507 33099
rect 14093 33099 14151 33105
rect 14093 33096 14105 33099
rect 13495 33068 14105 33096
rect 13495 33065 13507 33068
rect 13449 33059 13507 33065
rect 13814 32988 13820 33040
rect 13872 32988 13878 33040
rect 6914 32960 6920 32972
rect 3896 32932 6920 32960
rect 3896 32904 3924 32932
rect 6914 32920 6920 32932
rect 6972 32920 6978 32972
rect 12434 32920 12440 32972
rect 12492 32960 12498 32972
rect 13265 32963 13323 32969
rect 13265 32960 13277 32963
rect 12492 32932 13277 32960
rect 12492 32920 12498 32932
rect 13265 32929 13277 32932
rect 13311 32929 13323 32963
rect 13265 32923 13323 32929
rect 3878 32852 3884 32904
rect 3936 32852 3942 32904
rect 4801 32895 4859 32901
rect 4801 32861 4813 32895
rect 4847 32892 4859 32895
rect 4847 32864 5304 32892
rect 4847 32861 4859 32864
rect 4801 32855 4859 32861
rect 5276 32765 5304 32864
rect 5534 32852 5540 32904
rect 5592 32852 5598 32904
rect 5718 32852 5724 32904
rect 5776 32892 5782 32904
rect 5776 32864 6960 32892
rect 5776 32852 5782 32864
rect 5429 32827 5487 32833
rect 5429 32793 5441 32827
rect 5475 32824 5487 32827
rect 5552 32824 5580 32852
rect 5475 32796 5580 32824
rect 5629 32827 5687 32833
rect 5475 32793 5487 32796
rect 5429 32787 5487 32793
rect 5629 32793 5641 32827
rect 5675 32824 5687 32827
rect 6822 32824 6828 32836
rect 5675 32796 6828 32824
rect 5675 32793 5687 32796
rect 5629 32787 5687 32793
rect 6822 32784 6828 32796
rect 6880 32784 6886 32836
rect 5261 32759 5319 32765
rect 5261 32725 5273 32759
rect 5307 32725 5319 32759
rect 6932 32756 6960 32864
rect 12894 32852 12900 32904
rect 12952 32892 12958 32904
rect 13173 32895 13231 32901
rect 13173 32892 13185 32895
rect 12952 32864 13185 32892
rect 12952 32852 12958 32864
rect 13173 32861 13185 32864
rect 13219 32861 13231 32895
rect 13173 32855 13231 32861
rect 13354 32852 13360 32904
rect 13412 32892 13418 32904
rect 13924 32901 13952 33068
rect 14093 33065 14105 33068
rect 14139 33065 14151 33099
rect 14550 33096 14556 33108
rect 14093 33059 14151 33065
rect 14292 33068 14556 33096
rect 13449 32895 13507 32901
rect 13449 32892 13461 32895
rect 13412 32864 13461 32892
rect 13412 32852 13418 32864
rect 13449 32861 13461 32864
rect 13495 32861 13507 32895
rect 13449 32855 13507 32861
rect 13909 32895 13967 32901
rect 13909 32861 13921 32895
rect 13955 32861 13967 32895
rect 13909 32855 13967 32861
rect 14182 32852 14188 32904
rect 14240 32852 14246 32904
rect 14292 32901 14320 33068
rect 14550 33056 14556 33068
rect 14608 33096 14614 33108
rect 14608 33068 16988 33096
rect 14608 33056 14614 33068
rect 16960 33028 16988 33068
rect 17218 33056 17224 33108
rect 17276 33096 17282 33108
rect 17405 33099 17463 33105
rect 17405 33096 17417 33099
rect 17276 33068 17417 33096
rect 17276 33056 17282 33068
rect 17405 33065 17417 33068
rect 17451 33065 17463 33099
rect 17405 33059 17463 33065
rect 17586 33056 17592 33108
rect 17644 33096 17650 33108
rect 17957 33099 18015 33105
rect 17644 33068 17908 33096
rect 17644 33056 17650 33068
rect 17880 33028 17908 33068
rect 17957 33065 17969 33099
rect 18003 33096 18015 33099
rect 18506 33096 18512 33108
rect 18003 33068 18512 33096
rect 18003 33065 18015 33068
rect 17957 33059 18015 33065
rect 18506 33056 18512 33068
rect 18564 33056 18570 33108
rect 19426 33056 19432 33108
rect 19484 33056 19490 33108
rect 19889 33099 19947 33105
rect 19889 33065 19901 33099
rect 19935 33096 19947 33099
rect 20162 33096 20168 33108
rect 19935 33068 20168 33096
rect 19935 33065 19947 33068
rect 19889 33059 19947 33065
rect 20162 33056 20168 33068
rect 20220 33056 20226 33108
rect 21821 33099 21879 33105
rect 20917 33068 21772 33096
rect 20917 33028 20945 33068
rect 14384 33000 15792 33028
rect 16960 33000 17632 33028
rect 17880 33000 20945 33028
rect 14384 32901 14412 33000
rect 14458 32920 14464 32972
rect 14516 32960 14522 32972
rect 14645 32963 14703 32969
rect 14645 32960 14657 32963
rect 14516 32932 14657 32960
rect 14516 32920 14522 32932
rect 14645 32929 14657 32932
rect 14691 32929 14703 32963
rect 14645 32923 14703 32929
rect 15654 32920 15660 32972
rect 15712 32920 15718 32972
rect 15764 32960 15792 33000
rect 17604 32969 17632 33000
rect 20990 32988 20996 33040
rect 21048 32988 21054 33040
rect 21266 32988 21272 33040
rect 21324 32988 21330 33040
rect 17589 32963 17647 32969
rect 15764 32932 17356 32960
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 14369 32895 14427 32901
rect 14369 32861 14381 32895
rect 14415 32861 14427 32895
rect 14369 32855 14427 32861
rect 7190 32784 7196 32836
rect 7248 32784 7254 32836
rect 8478 32824 8484 32836
rect 8418 32796 8484 32824
rect 8478 32784 8484 32796
rect 8536 32824 8542 32836
rect 9306 32824 9312 32836
rect 8536 32796 9312 32824
rect 8536 32784 8542 32796
rect 9306 32784 9312 32796
rect 9364 32784 9370 32836
rect 14200 32824 14228 32852
rect 14737 32827 14795 32833
rect 14737 32824 14749 32827
rect 14200 32796 14749 32824
rect 14737 32793 14749 32796
rect 14783 32793 14795 32827
rect 14737 32787 14795 32793
rect 15930 32784 15936 32836
rect 15988 32784 15994 32836
rect 17218 32824 17224 32836
rect 17158 32796 17224 32824
rect 17218 32784 17224 32796
rect 17276 32784 17282 32836
rect 17328 32824 17356 32932
rect 17589 32929 17601 32963
rect 17635 32960 17647 32963
rect 19705 32963 19763 32969
rect 17635 32932 18920 32960
rect 17635 32929 17647 32932
rect 17589 32923 17647 32929
rect 18892 32904 18920 32932
rect 19705 32929 19717 32963
rect 19751 32960 19763 32963
rect 20346 32960 20352 32972
rect 19751 32932 20352 32960
rect 19751 32929 19763 32932
rect 19705 32923 19763 32929
rect 20346 32920 20352 32932
rect 20404 32920 20410 32972
rect 21008 32960 21036 32988
rect 20548 32932 21036 32960
rect 17773 32895 17831 32901
rect 17773 32861 17785 32895
rect 17819 32892 17831 32895
rect 17862 32892 17868 32904
rect 17819 32864 17868 32892
rect 17819 32861 17831 32864
rect 17773 32855 17831 32861
rect 17788 32824 17816 32855
rect 17862 32852 17868 32864
rect 17920 32852 17926 32904
rect 18874 32852 18880 32904
rect 18932 32852 18938 32904
rect 19981 32895 20039 32901
rect 19981 32861 19993 32895
rect 20027 32861 20039 32895
rect 19981 32855 20039 32861
rect 17328 32796 17816 32824
rect 18414 32784 18420 32836
rect 18472 32784 18478 32836
rect 11698 32756 11704 32768
rect 6932 32728 11704 32756
rect 5261 32719 5319 32725
rect 11698 32716 11704 32728
rect 11756 32716 11762 32768
rect 13633 32759 13691 32765
rect 13633 32725 13645 32759
rect 13679 32756 13691 32759
rect 18432 32756 18460 32784
rect 13679 32728 18460 32756
rect 19996 32756 20024 32855
rect 20070 32852 20076 32904
rect 20128 32892 20134 32904
rect 20548 32901 20576 32932
rect 20257 32895 20315 32901
rect 20257 32892 20269 32895
rect 20128 32864 20269 32892
rect 20128 32852 20134 32864
rect 20257 32861 20269 32864
rect 20303 32861 20315 32895
rect 20533 32895 20591 32901
rect 20533 32892 20545 32895
rect 20257 32855 20315 32861
rect 20364 32864 20545 32892
rect 20364 32833 20392 32864
rect 20533 32861 20545 32864
rect 20579 32861 20591 32895
rect 20533 32855 20591 32861
rect 20717 32895 20775 32901
rect 20717 32861 20729 32895
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 20349 32827 20407 32833
rect 20349 32793 20361 32827
rect 20395 32793 20407 32827
rect 20732 32824 20760 32855
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 20993 32895 21051 32901
rect 20993 32892 21005 32895
rect 20864 32864 21005 32892
rect 20864 32852 20870 32864
rect 20993 32861 21005 32864
rect 21039 32861 21051 32895
rect 20993 32855 21051 32861
rect 21269 32895 21327 32901
rect 21269 32861 21281 32895
rect 21315 32892 21327 32895
rect 21634 32892 21640 32904
rect 21315 32864 21640 32892
rect 21315 32861 21327 32864
rect 21269 32855 21327 32861
rect 21634 32852 21640 32864
rect 21692 32852 21698 32904
rect 21358 32824 21364 32836
rect 20732 32796 21364 32824
rect 20349 32787 20407 32793
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 21744 32824 21772 33068
rect 21821 33065 21833 33099
rect 21867 33096 21879 33099
rect 22278 33096 22284 33108
rect 21867 33068 22284 33096
rect 21867 33065 21879 33068
rect 21821 33059 21879 33065
rect 22278 33056 22284 33068
rect 22336 33096 22342 33108
rect 22738 33096 22744 33108
rect 22336 33068 22744 33096
rect 22336 33056 22342 33068
rect 22738 33056 22744 33068
rect 22796 33056 22802 33108
rect 23842 33056 23848 33108
rect 23900 33056 23906 33108
rect 24670 33056 24676 33108
rect 24728 33056 24734 33108
rect 26510 33056 26516 33108
rect 26568 33056 26574 33108
rect 28626 33056 28632 33108
rect 28684 33056 28690 33108
rect 34698 33056 34704 33108
rect 34756 33056 34762 33108
rect 34790 33056 34796 33108
rect 34848 33096 34854 33108
rect 34885 33099 34943 33105
rect 34885 33096 34897 33099
rect 34848 33068 34897 33096
rect 34848 33056 34854 33068
rect 34885 33065 34897 33068
rect 34931 33065 34943 33099
rect 34885 33059 34943 33065
rect 35161 33099 35219 33105
rect 35161 33065 35173 33099
rect 35207 33096 35219 33099
rect 35342 33096 35348 33108
rect 35207 33068 35348 33096
rect 35207 33065 35219 33068
rect 35161 33059 35219 33065
rect 23293 32963 23351 32969
rect 23293 32929 23305 32963
rect 23339 32960 23351 32963
rect 23860 32960 23888 33056
rect 23339 32932 23888 32960
rect 23339 32929 23351 32932
rect 23293 32923 23351 32929
rect 23566 32852 23572 32904
rect 23624 32852 23630 32904
rect 23658 32852 23664 32904
rect 23716 32892 23722 32904
rect 24397 32895 24455 32901
rect 24397 32892 24409 32895
rect 23716 32864 24409 32892
rect 23716 32852 23722 32864
rect 24397 32861 24409 32864
rect 24443 32861 24455 32895
rect 24397 32855 24455 32861
rect 24545 32895 24603 32901
rect 24545 32861 24557 32895
rect 24591 32892 24603 32895
rect 24688 32892 24716 33056
rect 25041 33031 25099 33037
rect 25041 32997 25053 33031
rect 25087 33028 25099 33031
rect 25087 33000 25912 33028
rect 25087 32997 25099 33000
rect 25041 32991 25099 32997
rect 25884 32969 25912 33000
rect 26326 32988 26332 33040
rect 26384 33028 26390 33040
rect 33870 33028 33876 33040
rect 26384 33000 33876 33028
rect 26384 32988 26390 33000
rect 33870 32988 33876 33000
rect 33928 32988 33934 33040
rect 34333 33031 34391 33037
rect 34333 32997 34345 33031
rect 34379 33028 34391 33031
rect 34716 33028 34744 33056
rect 35176 33028 35204 33059
rect 35342 33056 35348 33068
rect 35400 33056 35406 33108
rect 37921 33099 37979 33105
rect 37921 33065 37933 33099
rect 37967 33096 37979 33099
rect 38286 33096 38292 33108
rect 37967 33068 38292 33096
rect 37967 33065 37979 33068
rect 37921 33059 37979 33065
rect 38286 33056 38292 33068
rect 38344 33056 38350 33108
rect 40126 33056 40132 33108
rect 40184 33056 40190 33108
rect 34379 33000 34744 33028
rect 34379 32997 34391 33000
rect 34333 32991 34391 32997
rect 25869 32963 25927 32969
rect 25869 32929 25881 32963
rect 25915 32929 25927 32963
rect 25869 32923 25927 32929
rect 26881 32963 26939 32969
rect 26881 32929 26893 32963
rect 26927 32960 26939 32963
rect 27246 32960 27252 32972
rect 26927 32932 27252 32960
rect 26927 32929 26939 32932
rect 26881 32923 26939 32929
rect 27246 32920 27252 32932
rect 27304 32920 27310 32972
rect 34514 32960 34520 32972
rect 33704 32932 34520 32960
rect 24765 32895 24823 32901
rect 24765 32892 24777 32895
rect 24591 32861 24624 32892
rect 24688 32864 24777 32892
rect 24545 32855 24624 32861
rect 24765 32861 24777 32864
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 21744 32796 22126 32824
rect 20254 32756 20260 32768
rect 19996 32728 20260 32756
rect 13679 32725 13691 32728
rect 13633 32719 13691 32725
rect 20254 32716 20260 32728
rect 20312 32756 20318 32768
rect 20533 32759 20591 32765
rect 20533 32756 20545 32759
rect 20312 32728 20545 32756
rect 20312 32716 20318 32728
rect 20533 32725 20545 32728
rect 20579 32725 20591 32759
rect 20533 32719 20591 32725
rect 21085 32759 21143 32765
rect 21085 32725 21097 32759
rect 21131 32756 21143 32759
rect 21174 32756 21180 32768
rect 21131 32728 21180 32756
rect 21131 32725 21143 32728
rect 21085 32719 21143 32725
rect 21174 32716 21180 32728
rect 21232 32716 21238 32768
rect 24596 32756 24624 32855
rect 24854 32852 24860 32904
rect 24912 32901 24918 32904
rect 24912 32892 24920 32901
rect 25777 32895 25835 32901
rect 24912 32864 24957 32892
rect 24912 32855 24920 32864
rect 25777 32861 25789 32895
rect 25823 32892 25835 32895
rect 26418 32892 26424 32904
rect 25823 32864 26424 32892
rect 25823 32861 25835 32864
rect 25777 32855 25835 32861
rect 24912 32852 24918 32855
rect 26418 32852 26424 32864
rect 26476 32852 26482 32904
rect 26605 32895 26663 32901
rect 26605 32861 26617 32895
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 24670 32784 24676 32836
rect 24728 32784 24734 32836
rect 25682 32784 25688 32836
rect 25740 32824 25746 32836
rect 26620 32824 26648 32855
rect 27154 32852 27160 32904
rect 27212 32852 27218 32904
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32892 31171 32895
rect 31386 32892 31392 32904
rect 31159 32864 31392 32892
rect 31159 32861 31171 32864
rect 31113 32855 31171 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 31573 32895 31631 32901
rect 31573 32861 31585 32895
rect 31619 32861 31631 32895
rect 31573 32855 31631 32861
rect 25740 32796 26648 32824
rect 25740 32784 25746 32796
rect 31202 32784 31208 32836
rect 31260 32824 31266 32836
rect 31297 32827 31355 32833
rect 31297 32824 31309 32827
rect 31260 32796 31309 32824
rect 31260 32784 31266 32796
rect 31297 32793 31309 32796
rect 31343 32824 31355 32827
rect 31588 32824 31616 32855
rect 33502 32852 33508 32904
rect 33560 32892 33566 32904
rect 33704 32901 33732 32932
rect 34514 32920 34520 32932
rect 34572 32920 34578 32972
rect 34716 32960 34744 33000
rect 34900 33000 35204 33028
rect 40221 33031 40279 33037
rect 34793 32963 34851 32969
rect 34793 32960 34805 32963
rect 34716 32932 34805 32960
rect 34793 32929 34805 32932
rect 34839 32929 34851 32963
rect 34793 32923 34851 32929
rect 33689 32895 33747 32901
rect 33689 32892 33701 32895
rect 33560 32864 33701 32892
rect 33560 32852 33566 32864
rect 33689 32861 33701 32864
rect 33735 32861 33747 32895
rect 33689 32855 33747 32861
rect 33873 32895 33931 32901
rect 33873 32861 33885 32895
rect 33919 32892 33931 32895
rect 34054 32892 34060 32904
rect 33919 32864 34060 32892
rect 33919 32861 33931 32864
rect 33873 32855 33931 32861
rect 34054 32852 34060 32864
rect 34112 32852 34118 32904
rect 34149 32895 34207 32901
rect 34149 32861 34161 32895
rect 34195 32861 34207 32895
rect 34149 32855 34207 32861
rect 34701 32895 34759 32901
rect 34701 32861 34713 32895
rect 34747 32892 34759 32895
rect 34900 32892 34928 33000
rect 40221 32997 40233 33031
rect 40267 33028 40279 33031
rect 40402 33028 40408 33040
rect 40267 33000 40408 33028
rect 40267 32997 40279 33000
rect 40221 32991 40279 32997
rect 40402 32988 40408 33000
rect 40460 32988 40466 33040
rect 43717 33031 43775 33037
rect 43717 32997 43729 33031
rect 43763 33028 43775 33031
rect 44082 33028 44088 33040
rect 43763 33000 44088 33028
rect 43763 32997 43775 33000
rect 43717 32991 43775 32997
rect 44082 32988 44088 33000
rect 44140 32988 44146 33040
rect 34977 32963 35035 32969
rect 34977 32929 34989 32963
rect 35023 32929 35035 32963
rect 34977 32923 35035 32929
rect 34747 32864 34928 32892
rect 34992 32892 35020 32923
rect 43346 32920 43352 32972
rect 43404 32960 43410 32972
rect 43530 32960 43536 32972
rect 43404 32932 43536 32960
rect 43404 32920 43410 32932
rect 43530 32920 43536 32932
rect 43588 32920 43594 32972
rect 35069 32895 35127 32901
rect 35069 32892 35081 32895
rect 34992 32864 35081 32892
rect 34747 32861 34759 32864
rect 34701 32855 34759 32861
rect 34164 32824 34192 32855
rect 34992 32824 35020 32864
rect 35069 32861 35081 32864
rect 35115 32861 35127 32895
rect 35069 32855 35127 32861
rect 35250 32852 35256 32904
rect 35308 32852 35314 32904
rect 37642 32852 37648 32904
rect 37700 32892 37706 32904
rect 38562 32892 38568 32904
rect 37700 32864 38568 32892
rect 37700 32852 37706 32864
rect 38562 32852 38568 32864
rect 38620 32852 38626 32904
rect 40313 32895 40371 32901
rect 40313 32861 40325 32895
rect 40359 32892 40371 32895
rect 40586 32892 40592 32904
rect 40359 32864 40592 32892
rect 40359 32861 40371 32864
rect 40313 32855 40371 32861
rect 40586 32852 40592 32864
rect 40644 32852 40650 32904
rect 31343 32796 31616 32824
rect 33428 32796 34192 32824
rect 34532 32796 35020 32824
rect 31343 32793 31355 32796
rect 31297 32787 31355 32793
rect 33428 32768 33456 32796
rect 34532 32768 34560 32796
rect 39390 32784 39396 32836
rect 39448 32824 39454 32836
rect 40034 32824 40040 32836
rect 39448 32796 40040 32824
rect 39448 32784 39454 32796
rect 40034 32784 40040 32796
rect 40092 32784 40098 32836
rect 24946 32756 24952 32768
rect 24596 32728 24952 32756
rect 24946 32716 24952 32728
rect 25004 32756 25010 32768
rect 25133 32759 25191 32765
rect 25133 32756 25145 32759
rect 25004 32728 25145 32756
rect 25004 32716 25010 32728
rect 25133 32725 25145 32728
rect 25179 32725 25191 32759
rect 25133 32719 25191 32725
rect 30926 32716 30932 32768
rect 30984 32716 30990 32768
rect 31386 32716 31392 32768
rect 31444 32716 31450 32768
rect 33410 32716 33416 32768
rect 33468 32716 33474 32768
rect 34514 32716 34520 32768
rect 34572 32716 34578 32768
rect 43806 32716 43812 32768
rect 43864 32716 43870 32768
rect 1104 32666 44620 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 44620 32666
rect 1104 32592 44620 32614
rect 7190 32512 7196 32564
rect 7248 32552 7254 32564
rect 7837 32555 7895 32561
rect 7837 32552 7849 32555
rect 7248 32524 7849 32552
rect 7248 32512 7254 32524
rect 7837 32521 7849 32524
rect 7883 32521 7895 32555
rect 7837 32515 7895 32521
rect 8018 32512 8024 32564
rect 8076 32552 8082 32564
rect 8389 32555 8447 32561
rect 8389 32552 8401 32555
rect 8076 32524 8401 32552
rect 8076 32512 8082 32524
rect 8389 32521 8401 32524
rect 8435 32521 8447 32555
rect 8389 32515 8447 32521
rect 16485 32555 16543 32561
rect 16485 32521 16497 32555
rect 16531 32521 16543 32555
rect 16485 32515 16543 32521
rect 7006 32444 7012 32496
rect 7064 32484 7070 32496
rect 7101 32487 7159 32493
rect 7101 32484 7113 32487
rect 7064 32456 7113 32484
rect 7064 32444 7070 32456
rect 7101 32453 7113 32456
rect 7147 32484 7159 32487
rect 7282 32484 7288 32496
rect 7147 32456 7288 32484
rect 7147 32453 7159 32456
rect 7101 32447 7159 32453
rect 7282 32444 7288 32456
rect 7340 32444 7346 32496
rect 16500 32484 16528 32515
rect 16574 32512 16580 32564
rect 16632 32552 16638 32564
rect 16632 32524 19472 32552
rect 16632 32512 16638 32524
rect 16945 32487 17003 32493
rect 16945 32484 16957 32487
rect 8220 32456 12434 32484
rect 16500 32456 16957 32484
rect 6178 32376 6184 32428
rect 6236 32376 6242 32428
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32385 6883 32419
rect 6825 32379 6883 32385
rect 6840 32348 6868 32379
rect 8018 32376 8024 32428
rect 8076 32376 8082 32428
rect 7285 32351 7343 32357
rect 7285 32348 7297 32351
rect 6840 32320 7297 32348
rect 7285 32317 7297 32320
rect 7331 32348 7343 32351
rect 7650 32348 7656 32360
rect 7331 32320 7656 32348
rect 7331 32317 7343 32320
rect 7285 32311 7343 32317
rect 7650 32308 7656 32320
rect 7708 32348 7714 32360
rect 8220 32348 8248 32456
rect 8297 32419 8355 32425
rect 8297 32385 8309 32419
rect 8343 32385 8355 32419
rect 8297 32379 8355 32385
rect 8481 32419 8539 32425
rect 8481 32385 8493 32419
rect 8527 32416 8539 32419
rect 9122 32416 9128 32428
rect 8527 32388 9128 32416
rect 8527 32385 8539 32388
rect 8481 32379 8539 32385
rect 7708 32320 8248 32348
rect 8312 32348 8340 32379
rect 9122 32376 9128 32388
rect 9180 32376 9186 32428
rect 10597 32419 10655 32425
rect 10597 32385 10609 32419
rect 10643 32416 10655 32419
rect 11606 32416 11612 32428
rect 10643 32388 11612 32416
rect 10643 32385 10655 32388
rect 10597 32379 10655 32385
rect 11606 32376 11612 32388
rect 11664 32376 11670 32428
rect 11698 32376 11704 32428
rect 11756 32416 11762 32428
rect 12406 32416 12434 32456
rect 16945 32453 16957 32456
rect 16991 32453 17003 32487
rect 16945 32447 17003 32453
rect 17954 32444 17960 32496
rect 18012 32444 18018 32496
rect 11756 32388 12020 32416
rect 12406 32388 15608 32416
rect 11756 32376 11762 32388
rect 8312 32320 8524 32348
rect 7708 32308 7714 32320
rect 5166 32240 5172 32292
rect 5224 32280 5230 32292
rect 6641 32283 6699 32289
rect 6641 32280 6653 32283
rect 5224 32252 6653 32280
rect 5224 32240 5230 32252
rect 6641 32249 6653 32252
rect 6687 32280 6699 32283
rect 8386 32280 8392 32292
rect 6687 32252 8392 32280
rect 6687 32249 6699 32252
rect 6641 32243 6699 32249
rect 8386 32240 8392 32252
rect 8444 32240 8450 32292
rect 8496 32224 8524 32320
rect 9766 32308 9772 32360
rect 9824 32348 9830 32360
rect 10505 32351 10563 32357
rect 10505 32348 10517 32351
rect 9824 32320 10517 32348
rect 9824 32308 9830 32320
rect 10505 32317 10517 32320
rect 10551 32317 10563 32351
rect 11992 32348 12020 32388
rect 14642 32348 14648 32360
rect 11992 32320 14648 32348
rect 10505 32311 10563 32317
rect 14642 32308 14648 32320
rect 14700 32308 14706 32360
rect 15580 32280 15608 32388
rect 15654 32376 15660 32428
rect 15712 32376 15718 32428
rect 16298 32376 16304 32428
rect 16356 32376 16362 32428
rect 19444 32425 19472 32524
rect 22278 32512 22284 32564
rect 22336 32512 22342 32564
rect 26602 32552 26608 32564
rect 24872 32524 26608 32552
rect 22296 32425 22324 32512
rect 24872 32425 24900 32524
rect 26602 32512 26608 32524
rect 26660 32512 26666 32564
rect 27890 32512 27896 32564
rect 27948 32512 27954 32564
rect 33318 32512 33324 32564
rect 33376 32552 33382 32564
rect 34057 32555 34115 32561
rect 34057 32552 34069 32555
rect 33376 32524 34069 32552
rect 33376 32512 33382 32524
rect 34057 32521 34069 32524
rect 34103 32521 34115 32555
rect 34057 32515 34115 32521
rect 35250 32512 35256 32564
rect 35308 32552 35314 32564
rect 35621 32555 35679 32561
rect 35621 32552 35633 32555
rect 35308 32524 35633 32552
rect 35308 32512 35314 32524
rect 35621 32521 35633 32524
rect 35667 32521 35679 32555
rect 35621 32515 35679 32521
rect 43806 32512 43812 32564
rect 43864 32512 43870 32564
rect 26418 32444 26424 32496
rect 26476 32444 26482 32496
rect 31202 32484 31208 32496
rect 28000 32456 31208 32484
rect 19429 32419 19487 32425
rect 19429 32385 19441 32419
rect 19475 32385 19487 32419
rect 19429 32379 19487 32385
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32385 24915 32419
rect 24857 32379 24915 32385
rect 26234 32376 26240 32428
rect 26292 32376 26298 32428
rect 15672 32348 15700 32376
rect 16669 32351 16727 32357
rect 16669 32348 16681 32351
rect 15672 32320 16681 32348
rect 16669 32317 16681 32320
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 18417 32351 18475 32357
rect 18417 32317 18429 32351
rect 18463 32348 18475 32351
rect 19061 32351 19119 32357
rect 19061 32348 19073 32351
rect 18463 32320 19073 32348
rect 18463 32317 18475 32320
rect 18417 32311 18475 32317
rect 19061 32317 19073 32320
rect 19107 32348 19119 32351
rect 19245 32351 19303 32357
rect 19245 32348 19257 32351
rect 19107 32320 19257 32348
rect 19107 32317 19119 32320
rect 19061 32311 19119 32317
rect 19245 32317 19257 32320
rect 19291 32317 19303 32351
rect 19245 32311 19303 32317
rect 19613 32351 19671 32357
rect 19613 32317 19625 32351
rect 19659 32348 19671 32351
rect 23658 32348 23664 32360
rect 19659 32320 23664 32348
rect 19659 32317 19671 32320
rect 19613 32311 19671 32317
rect 23658 32308 23664 32320
rect 23716 32308 23722 32360
rect 25130 32308 25136 32360
rect 25188 32308 25194 32360
rect 15580 32252 16805 32280
rect 5810 32172 5816 32224
rect 5868 32212 5874 32224
rect 5997 32215 6055 32221
rect 5997 32212 6009 32215
rect 5868 32184 6009 32212
rect 5868 32172 5874 32184
rect 5997 32181 6009 32184
rect 6043 32181 6055 32215
rect 5997 32175 6055 32181
rect 8478 32172 8484 32224
rect 8536 32172 8542 32224
rect 10962 32172 10968 32224
rect 11020 32172 11026 32224
rect 11330 32172 11336 32224
rect 11388 32212 11394 32224
rect 15838 32212 15844 32224
rect 11388 32184 15844 32212
rect 11388 32172 11394 32184
rect 15838 32172 15844 32184
rect 15896 32172 15902 32224
rect 16777 32212 16805 32252
rect 18690 32240 18696 32292
rect 18748 32280 18754 32292
rect 24394 32280 24400 32292
rect 18748 32252 24400 32280
rect 18748 32240 18754 32252
rect 24394 32240 24400 32252
rect 24452 32240 24458 32292
rect 26252 32280 26280 32376
rect 26436 32348 26464 32444
rect 28000 32425 28028 32456
rect 31202 32444 31208 32456
rect 31260 32444 31266 32496
rect 31386 32444 31392 32496
rect 31444 32444 31450 32496
rect 33594 32444 33600 32496
rect 33652 32444 33658 32496
rect 34514 32484 34520 32496
rect 34164 32456 34520 32484
rect 27985 32419 28043 32425
rect 27985 32385 27997 32419
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 30926 32376 30932 32428
rect 30984 32376 30990 32428
rect 31113 32419 31171 32425
rect 31113 32385 31125 32419
rect 31159 32416 31171 32419
rect 31404 32416 31432 32444
rect 31159 32388 31432 32416
rect 31159 32385 31171 32388
rect 31113 32379 31171 32385
rect 26605 32351 26663 32357
rect 26605 32348 26617 32351
rect 26436 32320 26617 32348
rect 26605 32317 26617 32320
rect 26651 32317 26663 32351
rect 26605 32311 26663 32317
rect 29730 32308 29736 32360
rect 29788 32348 29794 32360
rect 30650 32348 30656 32360
rect 29788 32320 30656 32348
rect 29788 32308 29794 32320
rect 30650 32308 30656 32320
rect 30708 32308 30714 32360
rect 31294 32308 31300 32360
rect 31352 32348 31358 32360
rect 32122 32348 32128 32360
rect 31352 32320 32128 32348
rect 31352 32308 31358 32320
rect 32122 32308 32128 32320
rect 32180 32308 32186 32360
rect 33612 32348 33640 32444
rect 34164 32425 34192 32456
rect 34514 32444 34520 32456
rect 34572 32444 34578 32496
rect 35437 32487 35495 32493
rect 35437 32484 35449 32487
rect 34624 32456 35449 32484
rect 34624 32425 34652 32456
rect 35437 32453 35449 32456
rect 35483 32484 35495 32487
rect 35483 32456 35894 32484
rect 35483 32453 35495 32456
rect 35437 32447 35495 32453
rect 34149 32419 34207 32425
rect 34149 32385 34161 32419
rect 34195 32385 34207 32419
rect 34149 32379 34207 32385
rect 34425 32419 34483 32425
rect 34425 32385 34437 32419
rect 34471 32385 34483 32419
rect 34425 32379 34483 32385
rect 34609 32419 34667 32425
rect 34609 32385 34621 32419
rect 34655 32385 34667 32419
rect 34609 32379 34667 32385
rect 34440 32348 34468 32379
rect 34698 32376 34704 32428
rect 34756 32416 34762 32428
rect 34793 32419 34851 32425
rect 34793 32416 34805 32419
rect 34756 32388 34805 32416
rect 34756 32376 34762 32388
rect 34793 32385 34805 32388
rect 34839 32385 34851 32419
rect 34793 32379 34851 32385
rect 35253 32419 35311 32425
rect 35253 32385 35265 32419
rect 35299 32385 35311 32419
rect 35253 32379 35311 32385
rect 35268 32348 35296 32379
rect 33612 32320 35296 32348
rect 35866 32348 35894 32456
rect 42061 32419 42119 32425
rect 42061 32385 42073 32419
rect 42107 32416 42119 32419
rect 42426 32416 42432 32428
rect 42107 32388 42432 32416
rect 42107 32385 42119 32388
rect 42061 32379 42119 32385
rect 42426 32376 42432 32388
rect 42484 32376 42490 32428
rect 43533 32419 43591 32425
rect 43533 32385 43545 32419
rect 43579 32416 43591 32419
rect 43824 32416 43852 32512
rect 43579 32388 43852 32416
rect 43579 32385 43591 32388
rect 43533 32379 43591 32385
rect 36170 32348 36176 32360
rect 35866 32320 36176 32348
rect 36170 32308 36176 32320
rect 36228 32308 36234 32360
rect 26878 32280 26884 32292
rect 26252 32252 26884 32280
rect 26878 32240 26884 32252
rect 26936 32240 26942 32292
rect 30576 32252 31156 32280
rect 30576 32224 30604 32252
rect 17586 32212 17592 32224
rect 16777 32184 17592 32212
rect 17586 32172 17592 32184
rect 17644 32212 17650 32224
rect 18046 32212 18052 32224
rect 17644 32184 18052 32212
rect 17644 32172 17650 32184
rect 18046 32172 18052 32184
rect 18104 32172 18110 32224
rect 18506 32172 18512 32224
rect 18564 32172 18570 32224
rect 20806 32172 20812 32224
rect 20864 32212 20870 32224
rect 21174 32212 21180 32224
rect 20864 32184 21180 32212
rect 20864 32172 20870 32184
rect 21174 32172 21180 32184
rect 21232 32172 21238 32224
rect 22186 32172 22192 32224
rect 22244 32172 22250 32224
rect 30558 32172 30564 32224
rect 30616 32172 30622 32224
rect 31018 32172 31024 32224
rect 31076 32172 31082 32224
rect 31128 32212 31156 32252
rect 31202 32240 31208 32292
rect 31260 32280 31266 32292
rect 31570 32280 31576 32292
rect 31260 32252 31576 32280
rect 31260 32240 31266 32252
rect 31570 32240 31576 32252
rect 31628 32280 31634 32292
rect 33778 32280 33784 32292
rect 31628 32252 33784 32280
rect 31628 32240 31634 32252
rect 33778 32240 33784 32252
rect 33836 32280 33842 32292
rect 34977 32283 35035 32289
rect 34977 32280 34989 32283
rect 33836 32252 34989 32280
rect 33836 32240 33842 32252
rect 34977 32249 34989 32252
rect 35023 32249 35035 32283
rect 34977 32243 35035 32249
rect 35342 32212 35348 32224
rect 31128 32184 35348 32212
rect 35342 32172 35348 32184
rect 35400 32212 35406 32224
rect 38010 32212 38016 32224
rect 35400 32184 38016 32212
rect 35400 32172 35406 32184
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 42242 32172 42248 32224
rect 42300 32172 42306 32224
rect 43346 32172 43352 32224
rect 43404 32172 43410 32224
rect 1104 32122 44620 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 44620 32122
rect 1104 32048 44620 32070
rect 7190 31968 7196 32020
rect 7248 32008 7254 32020
rect 7742 32008 7748 32020
rect 7248 31980 7748 32008
rect 7248 31968 7254 31980
rect 7742 31968 7748 31980
rect 7800 31968 7806 32020
rect 7837 32011 7895 32017
rect 7837 31977 7849 32011
rect 7883 32008 7895 32011
rect 8113 32011 8171 32017
rect 8113 32008 8125 32011
rect 7883 31980 8125 32008
rect 7883 31977 7895 31980
rect 7837 31971 7895 31977
rect 8113 31977 8125 31980
rect 8159 31977 8171 32011
rect 8113 31971 8171 31977
rect 10962 31968 10968 32020
rect 11020 31968 11026 32020
rect 11057 32011 11115 32017
rect 11057 31977 11069 32011
rect 11103 32008 11115 32011
rect 11238 32008 11244 32020
rect 11103 31980 11244 32008
rect 11103 31977 11115 31980
rect 11057 31971 11115 31977
rect 11238 31968 11244 31980
rect 11296 31968 11302 32020
rect 11330 31968 11336 32020
rect 11388 32008 11394 32020
rect 11388 31980 11744 32008
rect 11388 31968 11394 31980
rect 6932 31912 7972 31940
rect 6932 31884 6960 31912
rect 3878 31832 3884 31884
rect 3936 31872 3942 31884
rect 5445 31875 5503 31881
rect 5445 31872 5457 31875
rect 3936 31844 5457 31872
rect 3936 31832 3942 31844
rect 5445 31841 5457 31844
rect 5491 31841 5503 31875
rect 5445 31835 5503 31841
rect 5721 31875 5779 31881
rect 5721 31841 5733 31875
rect 5767 31872 5779 31875
rect 5810 31872 5816 31884
rect 5767 31844 5816 31872
rect 5767 31841 5779 31844
rect 5721 31835 5779 31841
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 6914 31832 6920 31884
rect 6972 31832 6978 31884
rect 7944 31872 7972 31912
rect 8018 31900 8024 31952
rect 8076 31900 8082 31952
rect 10980 31940 11008 31968
rect 9140 31912 9444 31940
rect 10980 31912 11652 31940
rect 7944 31844 9076 31872
rect 8570 31804 8576 31816
rect 7852 31776 8576 31804
rect 5166 31696 5172 31748
rect 5224 31736 5230 31748
rect 5224 31708 6210 31736
rect 5224 31696 5230 31708
rect 7098 31696 7104 31748
rect 7156 31736 7162 31748
rect 7653 31739 7711 31745
rect 7653 31736 7665 31739
rect 7156 31708 7665 31736
rect 7156 31696 7162 31708
rect 7653 31705 7665 31708
rect 7699 31736 7711 31739
rect 7742 31736 7748 31748
rect 7699 31708 7748 31736
rect 7699 31705 7711 31708
rect 7653 31699 7711 31705
rect 7742 31696 7748 31708
rect 7800 31696 7806 31748
rect 7852 31745 7880 31776
rect 8570 31764 8576 31776
rect 8628 31804 8634 31816
rect 8941 31807 8999 31813
rect 8941 31804 8953 31807
rect 8628 31776 8953 31804
rect 8628 31764 8634 31776
rect 8941 31773 8953 31776
rect 8987 31773 8999 31807
rect 8941 31767 8999 31773
rect 7852 31739 7911 31745
rect 7852 31708 7865 31739
rect 7853 31705 7865 31708
rect 7899 31705 7911 31739
rect 7853 31699 7911 31705
rect 8294 31696 8300 31748
rect 8352 31696 8358 31748
rect 8386 31696 8392 31748
rect 8444 31736 8450 31748
rect 8481 31739 8539 31745
rect 8481 31736 8493 31739
rect 8444 31708 8493 31736
rect 8444 31696 8450 31708
rect 8481 31705 8493 31708
rect 8527 31705 8539 31739
rect 9048 31736 9076 31844
rect 9140 31816 9168 31912
rect 9309 31875 9367 31881
rect 9309 31841 9321 31875
rect 9355 31841 9367 31875
rect 9416 31872 9444 31912
rect 9416 31844 10824 31872
rect 9309 31835 9367 31841
rect 9122 31764 9128 31816
rect 9180 31764 9186 31816
rect 9324 31804 9352 31835
rect 9232 31776 9352 31804
rect 10796 31804 10824 31844
rect 10796 31776 11100 31804
rect 9232 31736 9260 31776
rect 9048 31708 9260 31736
rect 8481 31699 8539 31705
rect 9306 31696 9312 31748
rect 9364 31696 9370 31748
rect 9582 31696 9588 31748
rect 9640 31696 9646 31748
rect 9968 31708 10074 31736
rect 8312 31668 8340 31696
rect 8570 31668 8576 31680
rect 8312 31640 8576 31668
rect 8570 31628 8576 31640
rect 8628 31628 8634 31680
rect 9030 31628 9036 31680
rect 9088 31628 9094 31680
rect 9324 31668 9352 31696
rect 9968 31668 9996 31708
rect 9324 31640 9996 31668
rect 11072 31668 11100 31776
rect 11238 31764 11244 31816
rect 11296 31764 11302 31816
rect 11624 31813 11652 31912
rect 11716 31813 11744 31980
rect 16298 31968 16304 32020
rect 16356 32008 16362 32020
rect 16761 32011 16819 32017
rect 16761 32008 16773 32011
rect 16356 31980 16773 32008
rect 16356 31968 16362 31980
rect 16761 31977 16773 31980
rect 16807 31977 16819 32011
rect 16761 31971 16819 31977
rect 19981 32011 20039 32017
rect 19981 31977 19993 32011
rect 20027 32008 20039 32011
rect 20254 32008 20260 32020
rect 20027 31980 20260 32008
rect 20027 31977 20039 31980
rect 19981 31971 20039 31977
rect 20254 31968 20260 31980
rect 20312 32008 20318 32020
rect 21269 32011 21327 32017
rect 21269 32008 21281 32011
rect 20312 31980 21281 32008
rect 20312 31968 20318 31980
rect 21269 31977 21281 31980
rect 21315 31977 21327 32011
rect 21269 31971 21327 31977
rect 24854 31968 24860 32020
rect 24912 31968 24918 32020
rect 25130 31968 25136 32020
rect 25188 32008 25194 32020
rect 25317 32011 25375 32017
rect 25317 32008 25329 32011
rect 25188 31980 25329 32008
rect 25188 31968 25194 31980
rect 25317 31977 25329 31980
rect 25363 31977 25375 32011
rect 25317 31971 25375 31977
rect 27154 31968 27160 32020
rect 27212 32008 27218 32020
rect 30558 32008 30564 32020
rect 27212 31980 30564 32008
rect 27212 31968 27218 31980
rect 30558 31968 30564 31980
rect 30616 31968 30622 32020
rect 30650 31968 30656 32020
rect 30708 32008 30714 32020
rect 31573 32011 31631 32017
rect 31573 32008 31585 32011
rect 30708 31980 31585 32008
rect 30708 31968 30714 31980
rect 31573 31977 31585 31980
rect 31619 31977 31631 32011
rect 31573 31971 31631 31977
rect 32122 31968 32128 32020
rect 32180 31968 32186 32020
rect 34054 31968 34060 32020
rect 34112 31968 34118 32020
rect 37001 32011 37059 32017
rect 37001 31977 37013 32011
rect 37047 32008 37059 32011
rect 37350 32011 37408 32017
rect 37350 32008 37362 32011
rect 37047 31980 37362 32008
rect 37047 31977 37059 31980
rect 37001 31971 37059 31977
rect 37350 31977 37362 31980
rect 37396 31977 37408 32011
rect 37350 31971 37408 31977
rect 37458 31968 37464 32020
rect 37516 32008 37522 32020
rect 39482 32008 39488 32020
rect 37516 31980 39488 32008
rect 37516 31968 37522 31980
rect 39482 31968 39488 31980
rect 39540 32008 39546 32020
rect 39853 32011 39911 32017
rect 39853 32008 39865 32011
rect 39540 31980 39865 32008
rect 39540 31968 39546 31980
rect 39853 31977 39865 31980
rect 39899 31977 39911 32011
rect 41601 32011 41659 32017
rect 41601 32008 41613 32011
rect 39853 31971 39911 31977
rect 41386 31980 41613 32008
rect 12253 31943 12311 31949
rect 12253 31909 12265 31943
rect 12299 31940 12311 31943
rect 12526 31940 12532 31952
rect 12299 31912 12532 31940
rect 12299 31909 12311 31912
rect 12253 31903 12311 31909
rect 12526 31900 12532 31912
rect 12584 31900 12590 31952
rect 15746 31940 15752 31952
rect 15028 31912 15752 31940
rect 15028 31872 15056 31912
rect 15746 31900 15752 31912
rect 15804 31900 15810 31952
rect 16390 31900 16396 31952
rect 16448 31900 16454 31952
rect 19426 31900 19432 31952
rect 19484 31940 19490 31952
rect 19613 31943 19671 31949
rect 19613 31940 19625 31943
rect 19484 31912 19625 31940
rect 19484 31900 19490 31912
rect 19613 31909 19625 31912
rect 19659 31909 19671 31943
rect 19613 31903 19671 31909
rect 20165 31943 20223 31949
rect 20165 31909 20177 31943
rect 20211 31940 20223 31943
rect 20806 31940 20812 31952
rect 20211 31912 20812 31940
rect 20211 31909 20223 31912
rect 20165 31903 20223 31909
rect 20806 31900 20812 31912
rect 20864 31900 20870 31952
rect 24872 31940 24900 31968
rect 31021 31943 31079 31949
rect 31021 31940 31033 31943
rect 24872 31912 25176 31940
rect 15194 31872 15200 31884
rect 11900 31844 15056 31872
rect 15120 31844 15200 31872
rect 11900 31813 11928 31844
rect 12158 31813 12164 31816
rect 11609 31807 11667 31813
rect 11609 31773 11621 31807
rect 11655 31773 11667 31807
rect 11609 31767 11667 31773
rect 11702 31807 11760 31813
rect 11702 31773 11714 31807
rect 11748 31773 11760 31807
rect 11702 31767 11760 31773
rect 11885 31807 11943 31813
rect 11885 31773 11897 31807
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 12115 31807 12164 31813
rect 12115 31773 12127 31807
rect 12161 31773 12164 31807
rect 12115 31767 12164 31773
rect 12158 31764 12164 31767
rect 12216 31764 12222 31816
rect 12434 31804 12440 31816
rect 12268 31776 12440 31804
rect 11974 31696 11980 31748
rect 12032 31736 12038 31748
rect 12268 31736 12296 31776
rect 12434 31764 12440 31776
rect 12492 31764 12498 31816
rect 15120 31813 15148 31844
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 16408 31872 16436 31900
rect 15396 31844 16436 31872
rect 15008 31807 15066 31813
rect 15008 31773 15020 31807
rect 15054 31773 15066 31807
rect 15008 31767 15066 31773
rect 15105 31807 15163 31813
rect 15105 31773 15117 31807
rect 15151 31773 15163 31807
rect 15105 31767 15163 31773
rect 12032 31708 12296 31736
rect 12032 31696 12038 31708
rect 11333 31671 11391 31677
rect 11333 31668 11345 31671
rect 11072 31640 11345 31668
rect 11333 31637 11345 31640
rect 11379 31668 11391 31671
rect 11698 31668 11704 31680
rect 11379 31640 11704 31668
rect 11379 31637 11391 31640
rect 11333 31631 11391 31637
rect 11698 31628 11704 31640
rect 11756 31628 11762 31680
rect 14366 31628 14372 31680
rect 14424 31668 14430 31680
rect 14829 31671 14887 31677
rect 14829 31668 14841 31671
rect 14424 31640 14841 31668
rect 14424 31628 14430 31640
rect 14829 31637 14841 31640
rect 14875 31637 14887 31671
rect 15028 31668 15056 31767
rect 15286 31764 15292 31816
rect 15344 31804 15350 31816
rect 15396 31813 15424 31844
rect 17310 31832 17316 31884
rect 17368 31832 17374 31884
rect 20714 31832 20720 31884
rect 20772 31872 20778 31884
rect 20772 31844 21036 31872
rect 20772 31832 20778 31844
rect 15380 31807 15438 31813
rect 15380 31804 15392 31807
rect 15344 31776 15392 31804
rect 15344 31764 15350 31776
rect 15380 31773 15392 31776
rect 15426 31773 15438 31807
rect 15380 31767 15438 31773
rect 15470 31764 15476 31816
rect 15528 31764 15534 31816
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 15948 31776 17233 31804
rect 15197 31739 15255 31745
rect 15197 31705 15209 31739
rect 15243 31736 15255 31739
rect 15562 31736 15568 31748
rect 15243 31708 15568 31736
rect 15243 31705 15255 31708
rect 15197 31699 15255 31705
rect 15562 31696 15568 31708
rect 15620 31696 15626 31748
rect 15102 31668 15108 31680
rect 15028 31640 15108 31668
rect 14829 31631 14887 31637
rect 15102 31628 15108 31640
rect 15160 31668 15166 31680
rect 15948 31668 15976 31776
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 18506 31764 18512 31816
rect 18564 31764 18570 31816
rect 20438 31764 20444 31816
rect 20496 31804 20502 31816
rect 20901 31807 20959 31813
rect 20901 31804 20913 31807
rect 20496 31776 20913 31804
rect 20496 31764 20502 31776
rect 20901 31773 20913 31776
rect 20947 31773 20959 31807
rect 20901 31767 20959 31773
rect 17129 31739 17187 31745
rect 17129 31705 17141 31739
rect 17175 31736 17187 31739
rect 18524 31736 18552 31764
rect 17175 31708 18552 31736
rect 17175 31705 17187 31708
rect 17129 31699 17187 31705
rect 19334 31696 19340 31748
rect 19392 31736 19398 31748
rect 19392 31708 20116 31736
rect 19392 31696 19398 31708
rect 20088 31680 20116 31708
rect 20162 31696 20168 31748
rect 20220 31736 20226 31748
rect 20625 31739 20683 31745
rect 20625 31736 20637 31739
rect 20220 31708 20637 31736
rect 20220 31696 20226 31708
rect 20625 31705 20637 31708
rect 20671 31705 20683 31739
rect 20625 31699 20683 31705
rect 20809 31739 20867 31745
rect 20809 31705 20821 31739
rect 20855 31736 20867 31739
rect 21008 31736 21036 31844
rect 24946 31832 24952 31884
rect 25004 31872 25010 31884
rect 25004 31844 25084 31872
rect 25004 31832 25010 31844
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 20855 31708 21036 31736
rect 21100 31736 21128 31767
rect 24026 31764 24032 31816
rect 24084 31804 24090 31816
rect 24854 31813 24860 31816
rect 24673 31807 24731 31813
rect 24673 31804 24685 31807
rect 24084 31776 24685 31804
rect 24084 31764 24090 31776
rect 24673 31773 24685 31776
rect 24719 31773 24731 31807
rect 24673 31767 24731 31773
rect 24821 31807 24860 31813
rect 24821 31773 24833 31807
rect 24821 31767 24860 31773
rect 24854 31764 24860 31767
rect 24912 31764 24918 31816
rect 25056 31813 25084 31844
rect 25148 31813 25176 31912
rect 29840 31912 31033 31940
rect 29734 31817 29792 31823
rect 29734 31816 29746 31817
rect 29780 31816 29792 31817
rect 25041 31807 25099 31813
rect 25041 31773 25053 31807
rect 25087 31773 25099 31807
rect 25041 31767 25099 31773
rect 25138 31807 25196 31813
rect 25138 31773 25150 31807
rect 25184 31773 25196 31807
rect 29730 31804 29736 31816
rect 29702 31776 29736 31804
rect 25138 31767 25196 31773
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 29840 31813 29868 31912
rect 31021 31909 31033 31912
rect 31067 31909 31079 31943
rect 31021 31903 31079 31909
rect 31220 31912 31524 31940
rect 30193 31875 30251 31881
rect 30193 31841 30205 31875
rect 30239 31872 30251 31875
rect 30285 31875 30343 31881
rect 30285 31872 30297 31875
rect 30239 31844 30297 31872
rect 30239 31841 30251 31844
rect 30193 31835 30251 31841
rect 30285 31841 30297 31844
rect 30331 31841 30343 31875
rect 31220 31872 31248 31912
rect 30285 31835 30343 31841
rect 31036 31844 31248 31872
rect 31496 31872 31524 31912
rect 31754 31900 31760 31952
rect 31812 31940 31818 31952
rect 32140 31940 32168 31968
rect 41046 31940 41052 31952
rect 31812 31912 32168 31940
rect 31812 31900 31818 31912
rect 31496 31844 31892 31872
rect 31036 31816 31064 31844
rect 29825 31807 29883 31813
rect 29825 31773 29837 31807
rect 29871 31773 29883 31807
rect 29825 31767 29883 31773
rect 29914 31764 29920 31816
rect 29972 31764 29978 31816
rect 30098 31813 30104 31816
rect 30055 31807 30104 31813
rect 30055 31773 30067 31807
rect 30101 31773 30104 31807
rect 30055 31767 30104 31773
rect 30098 31764 30104 31767
rect 30156 31764 30162 31816
rect 30466 31764 30472 31816
rect 30524 31804 30530 31816
rect 30837 31807 30895 31813
rect 30837 31804 30849 31807
rect 30524 31776 30849 31804
rect 30524 31764 30530 31776
rect 30837 31773 30849 31776
rect 30883 31804 30895 31807
rect 30883 31776 30917 31804
rect 30883 31773 30895 31776
rect 30837 31767 30895 31773
rect 21542 31736 21548 31748
rect 21100 31708 21548 31736
rect 20855 31705 20867 31708
rect 20809 31699 20867 31705
rect 21542 31696 21548 31708
rect 21600 31696 21606 31748
rect 24578 31696 24584 31748
rect 24636 31736 24642 31748
rect 24949 31739 25007 31745
rect 24949 31736 24961 31739
rect 24636 31708 24961 31736
rect 24636 31696 24642 31708
rect 24949 31705 24961 31708
rect 24995 31736 25007 31739
rect 26418 31736 26424 31748
rect 24995 31708 26424 31736
rect 24995 31705 25007 31708
rect 24949 31699 25007 31705
rect 26418 31696 26424 31708
rect 26476 31696 26482 31748
rect 27080 31708 29684 31736
rect 27080 31680 27108 31708
rect 15160 31640 15976 31668
rect 15160 31628 15166 31640
rect 19978 31628 19984 31680
rect 20036 31628 20042 31680
rect 20070 31628 20076 31680
rect 20128 31628 20134 31680
rect 20254 31628 20260 31680
rect 20312 31628 20318 31680
rect 20438 31628 20444 31680
rect 20496 31628 20502 31680
rect 20530 31628 20536 31680
rect 20588 31628 20594 31680
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 24486 31668 24492 31680
rect 21048 31640 24492 31668
rect 21048 31628 21054 31640
rect 24486 31628 24492 31640
rect 24544 31628 24550 31680
rect 27062 31628 27068 31680
rect 27120 31628 27126 31680
rect 29546 31628 29552 31680
rect 29604 31628 29610 31680
rect 29656 31668 29684 31708
rect 30742 31696 30748 31748
rect 30800 31736 30806 31748
rect 30852 31736 30880 31767
rect 31018 31764 31024 31816
rect 31076 31764 31082 31816
rect 31110 31764 31116 31816
rect 31168 31764 31174 31816
rect 31220 31813 31248 31844
rect 31205 31807 31263 31813
rect 31205 31773 31217 31807
rect 31251 31773 31263 31807
rect 31205 31767 31263 31773
rect 31294 31764 31300 31816
rect 31352 31804 31358 31816
rect 31404 31813 31524 31814
rect 31404 31807 31539 31813
rect 31404 31804 31493 31807
rect 31352 31786 31493 31804
rect 31352 31776 31432 31786
rect 31352 31764 31358 31776
rect 31481 31773 31493 31786
rect 31527 31773 31539 31807
rect 31481 31767 31539 31773
rect 31570 31764 31576 31816
rect 31628 31764 31634 31816
rect 31864 31813 31892 31844
rect 31938 31832 31944 31884
rect 31996 31832 32002 31884
rect 32140 31872 32168 31912
rect 38488 31912 39804 31940
rect 37093 31875 37151 31881
rect 32140 31844 32260 31872
rect 32232 31813 32260 31844
rect 37093 31841 37105 31875
rect 37139 31872 37151 31875
rect 38010 31872 38016 31884
rect 37139 31844 38016 31872
rect 37139 31841 37151 31844
rect 37093 31835 37151 31841
rect 38010 31832 38016 31844
rect 38068 31872 38074 31884
rect 38378 31872 38384 31884
rect 38068 31844 38384 31872
rect 38068 31832 38074 31844
rect 38378 31832 38384 31844
rect 38436 31832 38442 31884
rect 31849 31807 31907 31813
rect 31849 31773 31861 31807
rect 31895 31804 31907 31807
rect 32125 31807 32183 31813
rect 32125 31804 32137 31807
rect 31895 31776 32137 31804
rect 31895 31773 31907 31776
rect 31849 31767 31907 31773
rect 32125 31773 32137 31776
rect 32171 31773 32183 31807
rect 32125 31767 32183 31773
rect 32217 31807 32275 31813
rect 32217 31773 32229 31807
rect 32263 31773 32275 31807
rect 36449 31807 36507 31813
rect 36449 31804 36461 31807
rect 32217 31767 32275 31773
rect 32324 31776 36461 31804
rect 30800 31708 30880 31736
rect 31128 31736 31156 31764
rect 31389 31739 31447 31745
rect 31389 31736 31401 31739
rect 31128 31708 31401 31736
rect 30800 31696 30806 31708
rect 31389 31705 31401 31708
rect 31435 31705 31447 31739
rect 31389 31699 31447 31705
rect 31665 31739 31723 31745
rect 31665 31705 31677 31739
rect 31711 31736 31723 31739
rect 31754 31736 31760 31748
rect 31711 31708 31760 31736
rect 31711 31705 31723 31708
rect 31665 31699 31723 31705
rect 31754 31696 31760 31708
rect 31812 31696 31818 31748
rect 31941 31739 31999 31745
rect 31941 31705 31953 31739
rect 31987 31736 31999 31739
rect 32324 31736 32352 31776
rect 36449 31773 36461 31776
rect 36495 31773 36507 31807
rect 36449 31767 36507 31773
rect 36538 31764 36544 31816
rect 36596 31804 36602 31816
rect 36633 31807 36691 31813
rect 36633 31804 36645 31807
rect 36596 31776 36645 31804
rect 36596 31764 36602 31776
rect 36633 31773 36645 31776
rect 36679 31773 36691 31807
rect 36633 31767 36691 31773
rect 36725 31807 36783 31813
rect 36725 31773 36737 31807
rect 36771 31773 36783 31807
rect 36725 31767 36783 31773
rect 31987 31708 32352 31736
rect 31987 31705 31999 31708
rect 31941 31699 31999 31705
rect 33226 31696 33232 31748
rect 33284 31736 33290 31748
rect 34241 31739 34299 31745
rect 34241 31736 34253 31739
rect 33284 31708 34253 31736
rect 33284 31696 33290 31708
rect 34241 31705 34253 31708
rect 34287 31736 34299 31739
rect 34330 31736 34336 31748
rect 34287 31708 34336 31736
rect 34287 31705 34299 31708
rect 34241 31699 34299 31705
rect 34330 31696 34336 31708
rect 34388 31696 34394 31748
rect 34422 31696 34428 31748
rect 34480 31696 34486 31748
rect 36740 31736 36768 31767
rect 36814 31764 36820 31816
rect 36872 31813 36878 31816
rect 36872 31807 36899 31813
rect 36887 31773 36899 31807
rect 38488 31790 38516 31912
rect 39776 31884 39804 31912
rect 40052 31912 41052 31940
rect 40052 31884 40080 31912
rect 41046 31900 41052 31912
rect 41104 31900 41110 31952
rect 38562 31832 38568 31884
rect 38620 31872 38626 31884
rect 39666 31872 39672 31884
rect 38620 31844 39672 31872
rect 38620 31832 38626 31844
rect 39666 31832 39672 31844
rect 39724 31832 39730 31884
rect 39758 31832 39764 31884
rect 39816 31832 39822 31884
rect 40034 31832 40040 31884
rect 40092 31832 40098 31884
rect 40497 31875 40555 31881
rect 40497 31841 40509 31875
rect 40543 31872 40555 31875
rect 40543 31844 40908 31872
rect 40543 31841 40555 31844
rect 40497 31835 40555 31841
rect 40512 31804 40540 31835
rect 36872 31767 36899 31773
rect 38856 31776 40540 31804
rect 36872 31764 36878 31767
rect 37458 31736 37464 31748
rect 36740 31708 37464 31736
rect 37458 31696 37464 31708
rect 37516 31696 37522 31748
rect 36814 31668 36820 31680
rect 29656 31640 36820 31668
rect 36814 31628 36820 31640
rect 36872 31628 36878 31680
rect 38102 31628 38108 31680
rect 38160 31668 38166 31680
rect 38856 31677 38884 31776
rect 40770 31764 40776 31816
rect 40828 31764 40834 31816
rect 40880 31813 40908 31844
rect 40865 31807 40923 31813
rect 40865 31773 40877 31807
rect 40911 31773 40923 31807
rect 40865 31767 40923 31773
rect 41141 31807 41199 31813
rect 41141 31773 41153 31807
rect 41187 31804 41199 31807
rect 41386 31804 41414 31980
rect 41601 31977 41613 31980
rect 41647 32008 41659 32011
rect 42886 32008 42892 32020
rect 41647 31980 42892 32008
rect 41647 31977 41659 31980
rect 41601 31971 41659 31977
rect 42886 31968 42892 31980
rect 42944 31968 42950 32020
rect 42518 31832 42524 31884
rect 42576 31832 42582 31884
rect 42797 31875 42855 31881
rect 42797 31841 42809 31875
rect 42843 31872 42855 31875
rect 43346 31872 43352 31884
rect 42843 31844 43352 31872
rect 42843 31841 42855 31844
rect 42797 31835 42855 31841
rect 43346 31832 43352 31844
rect 43404 31832 43410 31884
rect 44266 31832 44272 31884
rect 44324 31832 44330 31884
rect 41187 31776 41414 31804
rect 41187 31773 41199 31776
rect 41141 31767 41199 31773
rect 42150 31764 42156 31816
rect 42208 31764 42214 31816
rect 39666 31696 39672 31748
rect 39724 31736 39730 31748
rect 40678 31736 40684 31748
rect 39724 31708 40684 31736
rect 39724 31696 39730 31708
rect 40678 31696 40684 31708
rect 40736 31696 40742 31748
rect 43438 31696 43444 31748
rect 43496 31696 43502 31748
rect 38841 31671 38899 31677
rect 38841 31668 38853 31671
rect 38160 31640 38853 31668
rect 38160 31628 38166 31640
rect 38841 31637 38853 31640
rect 38887 31637 38899 31671
rect 38841 31631 38899 31637
rect 39206 31628 39212 31680
rect 39264 31668 39270 31680
rect 39758 31668 39764 31680
rect 39264 31640 39764 31668
rect 39264 31628 39270 31640
rect 39758 31628 39764 31640
rect 39816 31628 39822 31680
rect 40589 31671 40647 31677
rect 40589 31637 40601 31671
rect 40635 31668 40647 31671
rect 41138 31668 41144 31680
rect 40635 31640 41144 31668
rect 40635 31637 40647 31640
rect 40589 31631 40647 31637
rect 41138 31628 41144 31640
rect 41196 31628 41202 31680
rect 1104 31578 44620 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 44620 31578
rect 1104 31504 44620 31526
rect 6181 31467 6239 31473
rect 6181 31433 6193 31467
rect 6227 31464 6239 31467
rect 6270 31464 6276 31476
rect 6227 31436 6276 31464
rect 6227 31433 6239 31436
rect 6181 31427 6239 31433
rect 6270 31424 6276 31436
rect 6328 31424 6334 31476
rect 8478 31424 8484 31476
rect 8536 31424 8542 31476
rect 9030 31424 9036 31476
rect 9088 31424 9094 31476
rect 9401 31467 9459 31473
rect 9401 31433 9413 31467
rect 9447 31464 9459 31467
rect 9582 31464 9588 31476
rect 9447 31436 9588 31464
rect 9447 31433 9459 31436
rect 9401 31427 9459 31433
rect 9582 31424 9588 31436
rect 9640 31424 9646 31476
rect 11974 31424 11980 31476
rect 12032 31424 12038 31476
rect 13998 31464 14004 31476
rect 13636 31436 14004 31464
rect 5813 31399 5871 31405
rect 5813 31365 5825 31399
rect 5859 31365 5871 31399
rect 5813 31359 5871 31365
rect 6029 31399 6087 31405
rect 6029 31365 6041 31399
rect 6075 31396 6087 31399
rect 7374 31396 7380 31408
rect 6075 31368 7380 31396
rect 6075 31365 6087 31368
rect 6029 31359 6087 31365
rect 5534 31288 5540 31340
rect 5592 31328 5598 31340
rect 5828 31328 5856 31359
rect 7374 31356 7380 31368
rect 7432 31356 7438 31408
rect 8110 31356 8116 31408
rect 8168 31356 8174 31408
rect 8496 31396 8524 31424
rect 9048 31396 9076 31424
rect 8496 31368 8892 31396
rect 7098 31328 7104 31340
rect 5592 31300 7104 31328
rect 5592 31288 5598 31300
rect 7098 31288 7104 31300
rect 7156 31288 7162 31340
rect 8297 31331 8355 31337
rect 8297 31297 8309 31331
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 8481 31331 8539 31337
rect 8481 31297 8493 31331
rect 8527 31328 8539 31331
rect 8570 31328 8576 31340
rect 8527 31300 8576 31328
rect 8527 31297 8539 31300
rect 8481 31291 8539 31297
rect 8312 31204 8340 31291
rect 8294 31152 8300 31204
rect 8352 31152 8358 31204
rect 8496 31192 8524 31291
rect 8570 31288 8576 31300
rect 8628 31288 8634 31340
rect 8662 31288 8668 31340
rect 8720 31328 8726 31340
rect 8757 31331 8815 31337
rect 8757 31328 8769 31331
rect 8720 31300 8769 31328
rect 8720 31288 8726 31300
rect 8757 31297 8769 31300
rect 8803 31297 8815 31331
rect 8757 31291 8815 31297
rect 8864 31260 8892 31368
rect 8956 31368 9076 31396
rect 8956 31337 8984 31368
rect 8941 31331 8999 31337
rect 8941 31297 8953 31331
rect 8987 31297 8999 31331
rect 8941 31291 8999 31297
rect 9033 31331 9091 31337
rect 9033 31297 9045 31331
rect 9079 31297 9091 31331
rect 9033 31291 9091 31297
rect 9048 31260 9076 31291
rect 9122 31288 9128 31340
rect 9180 31288 9186 31340
rect 11790 31288 11796 31340
rect 11848 31328 11854 31340
rect 11885 31331 11943 31337
rect 11885 31328 11897 31331
rect 11848 31300 11897 31328
rect 11848 31288 11854 31300
rect 11885 31297 11897 31300
rect 11931 31297 11943 31331
rect 11885 31291 11943 31297
rect 12618 31288 12624 31340
rect 12676 31328 12682 31340
rect 13636 31337 13664 31436
rect 13998 31424 14004 31436
rect 14056 31464 14062 31476
rect 14458 31464 14464 31476
rect 14056 31436 14464 31464
rect 14056 31424 14062 31436
rect 14458 31424 14464 31436
rect 14516 31424 14522 31476
rect 19334 31464 19340 31476
rect 14660 31436 19340 31464
rect 14660 31408 14688 31436
rect 19334 31424 19340 31436
rect 19392 31424 19398 31476
rect 19610 31424 19616 31476
rect 19668 31464 19674 31476
rect 21266 31464 21272 31476
rect 19668 31436 21272 31464
rect 19668 31424 19674 31436
rect 21266 31424 21272 31436
rect 21324 31424 21330 31476
rect 24854 31424 24860 31476
rect 24912 31424 24918 31476
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 32858 31464 32864 31476
rect 25096 31436 32864 31464
rect 25096 31424 25102 31436
rect 32858 31424 32864 31436
rect 32916 31424 32922 31476
rect 35253 31467 35311 31473
rect 33060 31436 33457 31464
rect 14550 31396 14556 31408
rect 14016 31368 14556 31396
rect 14016 31337 14044 31368
rect 14550 31356 14556 31368
rect 14608 31356 14614 31408
rect 14642 31356 14648 31408
rect 14700 31356 14706 31408
rect 15562 31396 15568 31408
rect 15212 31368 15568 31396
rect 13633 31331 13691 31337
rect 12676 31300 13492 31328
rect 12676 31288 12682 31300
rect 13170 31260 13176 31272
rect 8864 31232 9076 31260
rect 9324 31232 13176 31260
rect 9324 31192 9352 31232
rect 13170 31220 13176 31232
rect 13228 31220 13234 31272
rect 13464 31260 13492 31300
rect 13633 31297 13645 31331
rect 13679 31297 13691 31331
rect 13633 31291 13691 31297
rect 13909 31331 13967 31337
rect 13909 31297 13921 31331
rect 13955 31297 13967 31331
rect 13909 31291 13967 31297
rect 14001 31331 14059 31337
rect 14001 31297 14013 31331
rect 14047 31297 14059 31331
rect 14001 31291 14059 31297
rect 13722 31260 13728 31272
rect 13464 31232 13728 31260
rect 13722 31220 13728 31232
rect 13780 31220 13786 31272
rect 13924 31260 13952 31291
rect 14182 31288 14188 31340
rect 14240 31288 14246 31340
rect 14274 31288 14280 31340
rect 14332 31328 14338 31340
rect 14415 31331 14473 31337
rect 14415 31328 14427 31331
rect 14332 31300 14427 31328
rect 14332 31288 14338 31300
rect 14415 31297 14427 31300
rect 14461 31297 14473 31331
rect 14826 31328 14832 31340
rect 14787 31300 14832 31328
rect 14415 31291 14473 31297
rect 14826 31288 14832 31300
rect 14884 31288 14890 31340
rect 14918 31288 14924 31340
rect 14976 31288 14982 31340
rect 15212 31337 15240 31368
rect 15562 31356 15568 31368
rect 15620 31396 15626 31408
rect 16301 31399 16359 31405
rect 16301 31396 16313 31399
rect 15620 31368 16313 31396
rect 15620 31356 15626 31368
rect 16301 31365 16313 31368
rect 16347 31365 16359 31399
rect 20073 31399 20131 31405
rect 16301 31359 16359 31365
rect 18892 31368 19932 31396
rect 15197 31331 15255 31337
rect 15197 31297 15209 31331
rect 15243 31297 15255 31331
rect 15197 31291 15255 31297
rect 15286 31288 15292 31340
rect 15344 31288 15350 31340
rect 15746 31288 15752 31340
rect 15804 31288 15810 31340
rect 15838 31288 15844 31340
rect 15896 31288 15902 31340
rect 16117 31331 16175 31337
rect 16117 31297 16129 31331
rect 16163 31328 16175 31331
rect 16393 31331 16451 31337
rect 16163 31300 16344 31328
rect 16163 31297 16175 31300
rect 16117 31291 16175 31297
rect 14292 31260 14320 31288
rect 15565 31263 15623 31269
rect 15565 31260 15577 31263
rect 13924 31232 14320 31260
rect 15396 31232 15577 31260
rect 8496 31164 9352 31192
rect 9646 31164 14596 31192
rect 5994 31084 6000 31136
rect 6052 31084 6058 31136
rect 6825 31127 6883 31133
rect 6825 31093 6837 31127
rect 6871 31124 6883 31127
rect 6914 31124 6920 31136
rect 6871 31096 6920 31124
rect 6871 31093 6883 31096
rect 6825 31087 6883 31093
rect 6914 31084 6920 31096
rect 6972 31084 6978 31136
rect 7742 31084 7748 31136
rect 7800 31124 7806 31136
rect 9646 31124 9674 31164
rect 14568 31136 14596 31164
rect 15396 31136 15424 31232
rect 15565 31229 15577 31232
rect 15611 31229 15623 31263
rect 15565 31223 15623 31229
rect 15654 31220 15660 31272
rect 15712 31220 15718 31272
rect 15856 31260 15884 31288
rect 15933 31263 15991 31269
rect 15933 31260 15945 31263
rect 15856 31232 15945 31260
rect 15933 31229 15945 31232
rect 15979 31229 15991 31263
rect 15933 31223 15991 31229
rect 16022 31220 16028 31272
rect 16080 31220 16086 31272
rect 15470 31152 15476 31204
rect 15528 31152 15534 31204
rect 16316 31192 16344 31300
rect 16393 31297 16405 31331
rect 16439 31297 16451 31331
rect 16393 31291 16451 31297
rect 16408 31260 16436 31291
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 18892 31337 18920 31368
rect 18877 31331 18935 31337
rect 18877 31328 18889 31331
rect 16540 31300 18889 31328
rect 16540 31288 16546 31300
rect 18877 31297 18889 31300
rect 18923 31297 18935 31331
rect 18877 31291 18935 31297
rect 19061 31331 19119 31337
rect 19061 31297 19073 31331
rect 19107 31328 19119 31331
rect 19242 31328 19248 31340
rect 19107 31300 19248 31328
rect 19107 31297 19119 31300
rect 19061 31291 19119 31297
rect 19242 31288 19248 31300
rect 19300 31328 19306 31340
rect 19797 31331 19855 31337
rect 19797 31328 19809 31331
rect 19300 31300 19809 31328
rect 19300 31288 19306 31300
rect 19797 31297 19809 31300
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 19705 31263 19763 31269
rect 16408 31232 19656 31260
rect 18969 31195 19027 31201
rect 16316 31164 18460 31192
rect 7800 31096 9674 31124
rect 7800 31084 7806 31096
rect 13814 31084 13820 31136
rect 13872 31084 13878 31136
rect 14274 31084 14280 31136
rect 14332 31084 14338 31136
rect 14550 31084 14556 31136
rect 14608 31084 14614 31136
rect 15010 31084 15016 31136
rect 15068 31084 15074 31136
rect 15378 31084 15384 31136
rect 15436 31084 15442 31136
rect 15488 31124 15516 31152
rect 18432 31136 18460 31164
rect 18969 31161 18981 31195
rect 19015 31192 19027 31195
rect 19426 31192 19432 31204
rect 19015 31164 19432 31192
rect 19015 31161 19027 31164
rect 18969 31155 19027 31161
rect 19426 31152 19432 31164
rect 19484 31152 19490 31204
rect 15933 31127 15991 31133
rect 15933 31124 15945 31127
rect 15488 31096 15945 31124
rect 15933 31093 15945 31096
rect 15979 31093 15991 31127
rect 15933 31087 15991 31093
rect 18414 31084 18420 31136
rect 18472 31084 18478 31136
rect 19334 31084 19340 31136
rect 19392 31124 19398 31136
rect 19521 31127 19579 31133
rect 19521 31124 19533 31127
rect 19392 31096 19533 31124
rect 19392 31084 19398 31096
rect 19521 31093 19533 31096
rect 19567 31093 19579 31127
rect 19628 31124 19656 31232
rect 19705 31229 19717 31263
rect 19751 31260 19763 31263
rect 19904 31260 19932 31368
rect 20073 31365 20085 31399
rect 20119 31396 20131 31399
rect 20622 31396 20628 31408
rect 20119 31368 20628 31396
rect 20119 31365 20131 31368
rect 20073 31359 20131 31365
rect 20622 31356 20628 31368
rect 20680 31356 20686 31408
rect 20806 31356 20812 31408
rect 20864 31356 20870 31408
rect 21542 31396 21548 31408
rect 21008 31368 21548 31396
rect 21008 31328 21036 31368
rect 21542 31356 21548 31368
rect 21600 31356 21606 31408
rect 23566 31356 23572 31408
rect 23624 31356 23630 31408
rect 24872 31396 24900 31424
rect 25317 31399 25375 31405
rect 25317 31396 25329 31399
rect 24872 31368 25329 31396
rect 25317 31365 25329 31368
rect 25363 31396 25375 31399
rect 26329 31399 26387 31405
rect 26329 31396 26341 31399
rect 25363 31368 26341 31396
rect 25363 31365 25375 31368
rect 25317 31359 25375 31365
rect 26329 31365 26341 31368
rect 26375 31365 26387 31399
rect 26329 31359 26387 31365
rect 26418 31356 26424 31408
rect 26476 31356 26482 31408
rect 27522 31396 27528 31408
rect 26528 31368 27528 31396
rect 20180 31300 21036 31328
rect 20180 31269 20208 31300
rect 21082 31288 21088 31340
rect 21140 31288 21146 31340
rect 21358 31288 21364 31340
rect 21416 31288 21422 31340
rect 26232 31331 26290 31337
rect 26232 31297 26244 31331
rect 26278 31328 26290 31331
rect 26278 31300 26372 31328
rect 26278 31297 26290 31300
rect 26232 31291 26290 31297
rect 20165 31263 20223 31269
rect 20165 31260 20177 31263
rect 19751 31232 19932 31260
rect 19996 31232 20177 31260
rect 19751 31229 19763 31232
rect 19705 31223 19763 31229
rect 19794 31152 19800 31204
rect 19852 31192 19858 31204
rect 19996 31192 20024 31232
rect 20165 31229 20177 31232
rect 20211 31229 20223 31263
rect 20165 31223 20223 31229
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 21376 31260 21404 31288
rect 20864 31232 21404 31260
rect 20864 31220 20870 31232
rect 21542 31220 21548 31272
rect 21600 31220 21606 31272
rect 22554 31220 22560 31272
rect 22612 31220 22618 31272
rect 22830 31220 22836 31272
rect 22888 31220 22894 31272
rect 25866 31220 25872 31272
rect 25924 31220 25930 31272
rect 26344 31260 26372 31300
rect 26528 31260 26556 31368
rect 27522 31356 27528 31368
rect 27580 31356 27586 31408
rect 28626 31396 28632 31408
rect 28276 31368 28632 31396
rect 28276 31340 28304 31368
rect 28626 31356 28632 31368
rect 28684 31356 28690 31408
rect 30006 31396 30012 31408
rect 29762 31368 30012 31396
rect 30006 31356 30012 31368
rect 30064 31356 30070 31408
rect 31110 31396 31116 31408
rect 30668 31368 31116 31396
rect 26604 31331 26662 31337
rect 26604 31297 26616 31331
rect 26650 31297 26662 31331
rect 26604 31291 26662 31297
rect 26697 31331 26755 31337
rect 26697 31297 26709 31331
rect 26743 31328 26755 31331
rect 26786 31328 26792 31340
rect 26743 31300 26792 31328
rect 26743 31297 26755 31300
rect 26697 31291 26755 31297
rect 26344 31232 26556 31260
rect 26620 31260 26648 31291
rect 26786 31288 26792 31300
rect 26844 31288 26850 31340
rect 28258 31288 28264 31340
rect 28316 31288 28322 31340
rect 30374 31288 30380 31340
rect 30432 31288 30438 31340
rect 30466 31288 30472 31340
rect 30524 31288 30530 31340
rect 30668 31337 30696 31368
rect 31110 31356 31116 31368
rect 31168 31396 31174 31408
rect 31570 31396 31576 31408
rect 31168 31368 31576 31396
rect 31168 31356 31174 31368
rect 31570 31356 31576 31368
rect 31628 31356 31634 31408
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 30837 31331 30895 31337
rect 30837 31297 30849 31331
rect 30883 31328 30895 31331
rect 31386 31328 31392 31340
rect 30883 31300 31392 31328
rect 30883 31297 30895 31300
rect 30837 31291 30895 31297
rect 31386 31288 31392 31300
rect 31444 31288 31450 31340
rect 32953 31331 33011 31337
rect 32953 31297 32965 31331
rect 32999 31297 33011 31331
rect 33060 31328 33088 31436
rect 33429 31350 33457 31436
rect 35253 31433 35265 31467
rect 35299 31464 35311 31467
rect 35342 31464 35348 31476
rect 35299 31436 35348 31464
rect 35299 31433 35311 31436
rect 35253 31427 35311 31433
rect 35342 31424 35348 31436
rect 35400 31464 35406 31476
rect 35802 31464 35808 31476
rect 35400 31436 35808 31464
rect 35400 31424 35406 31436
rect 35802 31424 35808 31436
rect 35860 31424 35866 31476
rect 42061 31467 42119 31473
rect 38488 31436 40356 31464
rect 33781 31399 33839 31405
rect 33781 31365 33793 31399
rect 33827 31365 33839 31399
rect 33781 31359 33839 31365
rect 33428 31347 33457 31350
rect 33413 31341 33471 31347
rect 33118 31331 33176 31337
rect 33118 31328 33130 31331
rect 33060 31300 33130 31328
rect 32953 31291 33011 31297
rect 33118 31297 33130 31300
rect 33164 31297 33176 31331
rect 33118 31291 33176 31297
rect 27430 31260 27436 31272
rect 26620 31232 27436 31260
rect 27430 31220 27436 31232
rect 27488 31260 27494 31272
rect 27525 31263 27583 31269
rect 27525 31260 27537 31263
rect 27488 31232 27537 31260
rect 27488 31220 27494 31232
rect 27525 31229 27537 31232
rect 27571 31229 27583 31263
rect 27525 31223 27583 31229
rect 28169 31263 28227 31269
rect 28169 31229 28181 31263
rect 28215 31229 28227 31263
rect 28169 31223 28227 31229
rect 28537 31263 28595 31269
rect 28537 31229 28549 31263
rect 28583 31260 28595 31263
rect 29546 31260 29552 31272
rect 28583 31232 29552 31260
rect 28583 31229 28595 31232
rect 28537 31223 28595 31229
rect 19852 31164 20024 31192
rect 19852 31152 19858 31164
rect 20070 31152 20076 31204
rect 20128 31192 20134 31204
rect 21637 31195 21695 31201
rect 21637 31192 21649 31195
rect 20128 31164 21649 31192
rect 20128 31152 20134 31164
rect 21637 31161 21649 31164
rect 21683 31161 21695 31195
rect 21637 31155 21695 31161
rect 20898 31124 20904 31136
rect 19628 31096 20904 31124
rect 19521 31087 19579 31093
rect 20898 31084 20904 31096
rect 20956 31124 20962 31136
rect 23842 31124 23848 31136
rect 20956 31096 23848 31124
rect 20956 31084 20962 31096
rect 23842 31084 23848 31096
rect 23900 31124 23906 31136
rect 24305 31127 24363 31133
rect 24305 31124 24317 31127
rect 23900 31096 24317 31124
rect 23900 31084 23906 31096
rect 24305 31093 24317 31096
rect 24351 31093 24363 31127
rect 24305 31087 24363 31093
rect 26050 31084 26056 31136
rect 26108 31084 26114 31136
rect 28184 31124 28212 31223
rect 29546 31220 29552 31232
rect 29604 31220 29610 31272
rect 30009 31263 30067 31269
rect 30009 31229 30021 31263
rect 30055 31260 30067 31263
rect 30484 31260 30512 31288
rect 30055 31232 30512 31260
rect 32968 31260 32996 31291
rect 33226 31288 33232 31340
rect 33284 31288 33290 31340
rect 33413 31307 33425 31341
rect 33459 31328 33471 31341
rect 33459 31307 33548 31328
rect 33413 31301 33548 31307
rect 33428 31300 33548 31301
rect 33244 31260 33272 31288
rect 33520 31272 33548 31300
rect 32968 31232 33272 31260
rect 30055 31229 30067 31232
rect 30009 31223 30067 31229
rect 33502 31220 33508 31272
rect 33560 31220 33566 31272
rect 29638 31152 29644 31204
rect 29696 31192 29702 31204
rect 30561 31195 30619 31201
rect 30561 31192 30573 31195
rect 29696 31164 30573 31192
rect 29696 31152 29702 31164
rect 30561 31161 30573 31164
rect 30607 31161 30619 31195
rect 30561 31155 30619 31161
rect 31938 31152 31944 31204
rect 31996 31152 32002 31204
rect 32674 31152 32680 31204
rect 32732 31192 32738 31204
rect 33321 31195 33379 31201
rect 33321 31192 33333 31195
rect 32732 31164 33333 31192
rect 32732 31152 32738 31164
rect 33321 31161 33333 31164
rect 33367 31161 33379 31195
rect 33321 31155 33379 31161
rect 29270 31124 29276 31136
rect 28184 31096 29276 31124
rect 29270 31084 29276 31096
rect 29328 31084 29334 31136
rect 30193 31127 30251 31133
rect 30193 31093 30205 31127
rect 30239 31124 30251 31127
rect 31956 31124 31984 31152
rect 30239 31096 31984 31124
rect 30239 31093 30251 31096
rect 30193 31087 30251 31093
rect 32766 31084 32772 31136
rect 32824 31084 32830 31136
rect 32858 31084 32864 31136
rect 32916 31124 32922 31136
rect 33796 31124 33824 31359
rect 38488 31340 38516 31436
rect 38746 31356 38752 31408
rect 38804 31356 38810 31408
rect 39206 31356 39212 31408
rect 39264 31356 39270 31408
rect 38010 31288 38016 31340
rect 38068 31328 38074 31340
rect 38470 31328 38476 31340
rect 38068 31300 38476 31328
rect 38068 31288 38074 31300
rect 38470 31288 38476 31300
rect 38528 31288 38534 31340
rect 40328 31337 40356 31436
rect 42061 31433 42073 31467
rect 42107 31464 42119 31467
rect 42150 31464 42156 31476
rect 42107 31436 42156 31464
rect 42107 31433 42119 31436
rect 42061 31427 42119 31433
rect 42150 31424 42156 31436
rect 42208 31424 42214 31476
rect 42426 31424 42432 31476
rect 42484 31424 42490 31476
rect 42886 31424 42892 31476
rect 42944 31424 42950 31476
rect 40678 31356 40684 31408
rect 40736 31396 40742 31408
rect 40736 31368 41078 31396
rect 40736 31356 40742 31368
rect 40313 31331 40371 31337
rect 40313 31297 40325 31331
rect 40359 31297 40371 31331
rect 40313 31291 40371 31297
rect 42794 31288 42800 31340
rect 42852 31288 42858 31340
rect 38378 31220 38384 31272
rect 38436 31260 38442 31272
rect 38436 31232 40356 31260
rect 38436 31220 38442 31232
rect 39758 31152 39764 31204
rect 39816 31192 39822 31204
rect 40221 31195 40279 31201
rect 40221 31192 40233 31195
rect 39816 31164 40233 31192
rect 39816 31152 39822 31164
rect 40221 31161 40233 31164
rect 40267 31161 40279 31195
rect 40221 31155 40279 31161
rect 32916 31096 33824 31124
rect 32916 31084 32922 31096
rect 37918 31084 37924 31136
rect 37976 31124 37982 31136
rect 40034 31124 40040 31136
rect 37976 31096 40040 31124
rect 37976 31084 37982 31096
rect 40034 31084 40040 31096
rect 40092 31084 40098 31136
rect 40328 31124 40356 31232
rect 40586 31220 40592 31272
rect 40644 31220 40650 31272
rect 43073 31263 43131 31269
rect 43073 31229 43085 31263
rect 43119 31260 43131 31263
rect 43162 31260 43168 31272
rect 43119 31232 43168 31260
rect 43119 31229 43131 31232
rect 43073 31223 43131 31229
rect 43162 31220 43168 31232
rect 43220 31220 43226 31272
rect 40770 31124 40776 31136
rect 40328 31096 40776 31124
rect 40770 31084 40776 31096
rect 40828 31084 40834 31136
rect 1104 31034 44620 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 44620 31034
rect 1104 30960 44620 30982
rect 3878 30880 3884 30932
rect 3936 30880 3942 30932
rect 5994 30880 6000 30932
rect 6052 30920 6058 30932
rect 7469 30923 7527 30929
rect 7469 30920 7481 30923
rect 6052 30892 7481 30920
rect 6052 30880 6058 30892
rect 7469 30889 7481 30892
rect 7515 30889 7527 30923
rect 7469 30883 7527 30889
rect 8021 30923 8079 30929
rect 8021 30889 8033 30923
rect 8067 30920 8079 30923
rect 8294 30920 8300 30932
rect 8067 30892 8300 30920
rect 8067 30889 8079 30892
rect 8021 30883 8079 30889
rect 8294 30880 8300 30892
rect 8352 30880 8358 30932
rect 12805 30923 12863 30929
rect 12805 30889 12817 30923
rect 12851 30920 12863 30923
rect 13814 30920 13820 30932
rect 12851 30892 13820 30920
rect 12851 30889 12863 30892
rect 12805 30883 12863 30889
rect 13814 30880 13820 30892
rect 13872 30880 13878 30932
rect 14274 30929 14280 30932
rect 14258 30923 14280 30929
rect 14258 30889 14270 30923
rect 14258 30883 14280 30889
rect 14274 30880 14280 30883
rect 14332 30880 14338 30932
rect 14366 30880 14372 30932
rect 14424 30880 14430 30932
rect 14550 30880 14556 30932
rect 14608 30880 14614 30932
rect 15010 30880 15016 30932
rect 15068 30880 15074 30932
rect 17310 30880 17316 30932
rect 17368 30920 17374 30932
rect 19242 30920 19248 30932
rect 17368 30892 19248 30920
rect 17368 30880 17374 30892
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 19518 30880 19524 30932
rect 19576 30880 19582 30932
rect 19702 30880 19708 30932
rect 19760 30920 19766 30932
rect 20165 30923 20223 30929
rect 20165 30920 20177 30923
rect 19760 30892 20177 30920
rect 19760 30880 19766 30892
rect 20165 30889 20177 30892
rect 20211 30889 20223 30923
rect 20165 30883 20223 30889
rect 20441 30923 20499 30929
rect 20441 30889 20453 30923
rect 20487 30889 20499 30923
rect 20441 30883 20499 30889
rect 3789 30787 3847 30793
rect 3789 30753 3801 30787
rect 3835 30784 3847 30787
rect 3896 30784 3924 30880
rect 7009 30855 7067 30861
rect 7009 30821 7021 30855
rect 7055 30852 7067 30855
rect 7055 30824 7604 30852
rect 7055 30821 7067 30824
rect 7009 30815 7067 30821
rect 3835 30756 3924 30784
rect 4065 30787 4123 30793
rect 3835 30753 3847 30756
rect 3789 30747 3847 30753
rect 4065 30753 4077 30787
rect 4111 30784 4123 30787
rect 5997 30787 6055 30793
rect 5997 30784 6009 30787
rect 4111 30756 6009 30784
rect 4111 30753 4123 30756
rect 4065 30747 4123 30753
rect 5997 30753 6009 30756
rect 6043 30753 6055 30787
rect 5997 30747 6055 30753
rect 6641 30787 6699 30793
rect 6641 30753 6653 30787
rect 6687 30784 6699 30787
rect 7190 30784 7196 30796
rect 6687 30756 7196 30784
rect 6687 30753 6699 30756
rect 6641 30747 6699 30753
rect 7190 30744 7196 30756
rect 7248 30784 7254 30796
rect 7248 30756 7328 30784
rect 7248 30744 7254 30756
rect 5166 30676 5172 30728
rect 5224 30676 5230 30728
rect 5626 30676 5632 30728
rect 5684 30716 5690 30728
rect 5905 30719 5963 30725
rect 5905 30716 5917 30719
rect 5684 30688 5917 30716
rect 5684 30676 5690 30688
rect 5905 30685 5917 30688
rect 5951 30685 5963 30719
rect 5905 30679 5963 30685
rect 6086 30676 6092 30728
rect 6144 30676 6150 30728
rect 6825 30719 6883 30725
rect 6825 30685 6837 30719
rect 6871 30685 6883 30719
rect 6825 30679 6883 30685
rect 5810 30608 5816 30660
rect 5868 30608 5874 30660
rect 6104 30648 6132 30676
rect 6840 30648 6868 30679
rect 7300 30657 7328 30756
rect 7576 30728 7604 30824
rect 13078 30812 13084 30864
rect 13136 30812 13142 30864
rect 13170 30812 13176 30864
rect 13228 30852 13234 30864
rect 13228 30824 13308 30852
rect 13228 30812 13234 30824
rect 10413 30787 10471 30793
rect 10413 30753 10425 30787
rect 10459 30753 10471 30787
rect 10413 30747 10471 30753
rect 10873 30787 10931 30793
rect 10873 30753 10885 30787
rect 10919 30753 10931 30787
rect 13096 30784 13124 30812
rect 10873 30747 10931 30753
rect 11992 30756 13124 30784
rect 7558 30676 7564 30728
rect 7616 30676 7622 30728
rect 8021 30719 8079 30725
rect 8021 30716 8033 30719
rect 7668 30688 8033 30716
rect 7101 30651 7159 30657
rect 7101 30648 7113 30651
rect 6104 30620 7113 30648
rect 7101 30617 7113 30620
rect 7147 30617 7159 30651
rect 7101 30611 7159 30617
rect 7285 30651 7343 30657
rect 7285 30617 7297 30651
rect 7331 30617 7343 30651
rect 7285 30611 7343 30617
rect 7300 30580 7328 30611
rect 7374 30608 7380 30660
rect 7432 30648 7438 30660
rect 7668 30648 7696 30688
rect 8021 30685 8033 30688
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 8202 30676 8208 30728
rect 8260 30676 8266 30728
rect 7432 30620 7696 30648
rect 7432 30608 7438 30620
rect 7742 30608 7748 30660
rect 7800 30608 7806 30660
rect 10428 30648 10456 30747
rect 10502 30676 10508 30728
rect 10560 30676 10566 30728
rect 10888 30716 10916 30747
rect 11609 30719 11667 30725
rect 11609 30716 11621 30719
rect 10888 30688 11621 30716
rect 11609 30685 11621 30688
rect 11655 30685 11667 30719
rect 11609 30679 11667 30685
rect 11698 30676 11704 30728
rect 11756 30676 11762 30728
rect 11992 30725 12020 30756
rect 11977 30719 12035 30725
rect 11977 30685 11989 30719
rect 12023 30685 12035 30719
rect 11977 30679 12035 30685
rect 12066 30676 12072 30728
rect 12124 30725 12130 30728
rect 12124 30679 12132 30725
rect 12529 30719 12587 30725
rect 12529 30716 12541 30719
rect 12268 30688 12541 30716
rect 12124 30676 12130 30679
rect 7852 30620 10456 30648
rect 11885 30651 11943 30657
rect 7852 30580 7880 30620
rect 11885 30617 11897 30651
rect 11931 30648 11943 30651
rect 11931 30620 12020 30648
rect 11931 30617 11943 30620
rect 11885 30611 11943 30617
rect 11992 30592 12020 30620
rect 7300 30552 7880 30580
rect 7926 30540 7932 30592
rect 7984 30540 7990 30592
rect 11974 30540 11980 30592
rect 12032 30540 12038 30592
rect 12268 30589 12296 30688
rect 12529 30685 12541 30688
rect 12575 30685 12587 30719
rect 12529 30679 12587 30685
rect 12621 30719 12679 30725
rect 12621 30685 12633 30719
rect 12667 30685 12679 30719
rect 12621 30679 12679 30685
rect 12434 30608 12440 30660
rect 12492 30648 12498 30660
rect 12636 30648 12664 30679
rect 12894 30676 12900 30728
rect 12952 30716 12958 30728
rect 13056 30719 13114 30725
rect 13056 30716 13068 30719
rect 12952 30688 13068 30716
rect 12952 30676 12958 30688
rect 13056 30685 13068 30688
rect 13102 30685 13114 30719
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 13056 30679 13114 30685
rect 13152 30685 13185 30716
rect 13219 30685 13231 30719
rect 13280 30716 13308 30824
rect 13538 30812 13544 30864
rect 13596 30852 13602 30864
rect 15028 30852 15056 30880
rect 13596 30824 15056 30852
rect 13596 30812 13602 30824
rect 15746 30812 15752 30864
rect 15804 30852 15810 30864
rect 19610 30852 19616 30864
rect 15804 30824 19616 30852
rect 15804 30812 15810 30824
rect 19610 30812 19616 30824
rect 19668 30812 19674 30864
rect 19886 30852 19892 30864
rect 19812 30824 19892 30852
rect 13725 30787 13783 30793
rect 13725 30753 13737 30787
rect 13771 30784 13783 30787
rect 13771 30756 14044 30784
rect 13771 30753 13783 30756
rect 13725 30747 13783 30753
rect 13393 30719 13451 30725
rect 13393 30716 13405 30719
rect 13280 30688 13405 30716
rect 13152 30679 13231 30685
rect 13393 30685 13405 30688
rect 13439 30685 13451 30719
rect 13393 30679 13451 30685
rect 12492 30620 12664 30648
rect 12805 30651 12863 30657
rect 12492 30608 12498 30620
rect 12805 30617 12817 30651
rect 12851 30648 12863 30651
rect 13152 30648 13180 30679
rect 13538 30676 13544 30728
rect 13596 30676 13602 30728
rect 13641 30713 13699 30719
rect 13814 30718 13820 30728
rect 13641 30679 13653 30713
rect 13687 30710 13699 30713
rect 13740 30710 13820 30718
rect 13687 30690 13820 30710
rect 13687 30682 13768 30690
rect 13687 30679 13699 30682
rect 13641 30673 13699 30679
rect 13814 30676 13820 30690
rect 13872 30676 13878 30728
rect 12851 30620 12940 30648
rect 12851 30617 12863 30620
rect 12805 30611 12863 30617
rect 12253 30583 12311 30589
rect 12253 30549 12265 30583
rect 12299 30549 12311 30583
rect 12253 30543 12311 30549
rect 12342 30540 12348 30592
rect 12400 30540 12406 30592
rect 12912 30589 12940 30620
rect 13004 30620 13180 30648
rect 13265 30651 13323 30657
rect 13004 30592 13032 30620
rect 13265 30617 13277 30651
rect 13311 30648 13323 30651
rect 13311 30620 13400 30648
rect 13311 30617 13323 30620
rect 13265 30611 13323 30617
rect 13372 30592 13400 30620
rect 12897 30583 12955 30589
rect 12897 30549 12909 30583
rect 12943 30549 12955 30583
rect 12897 30543 12955 30549
rect 12986 30540 12992 30592
rect 13044 30540 13050 30592
rect 13354 30540 13360 30592
rect 13412 30540 13418 30592
rect 13906 30540 13912 30592
rect 13964 30580 13970 30592
rect 14016 30580 14044 30756
rect 14182 30744 14188 30796
rect 14240 30744 14246 30796
rect 14274 30744 14280 30796
rect 14332 30784 14338 30796
rect 14461 30787 14519 30793
rect 14461 30784 14473 30787
rect 14332 30756 14473 30784
rect 14332 30744 14338 30756
rect 14461 30753 14473 30756
rect 14507 30753 14519 30787
rect 14461 30747 14519 30753
rect 14826 30744 14832 30796
rect 14884 30784 14890 30796
rect 14884 30756 15240 30784
rect 14884 30744 14890 30756
rect 14200 30716 14228 30744
rect 15212 30725 15240 30756
rect 15378 30744 15384 30796
rect 15436 30784 15442 30796
rect 17126 30784 17132 30796
rect 15436 30756 17132 30784
rect 15436 30744 15442 30756
rect 17126 30744 17132 30756
rect 17184 30744 17190 30796
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30784 18751 30787
rect 19812 30784 19840 30824
rect 19886 30812 19892 30824
rect 19944 30812 19950 30864
rect 20070 30812 20076 30864
rect 20128 30812 20134 30864
rect 20456 30852 20484 30883
rect 20530 30880 20536 30932
rect 20588 30920 20594 30932
rect 20901 30923 20959 30929
rect 20901 30920 20913 30923
rect 20588 30892 20913 30920
rect 20588 30880 20594 30892
rect 20901 30889 20913 30892
rect 20947 30889 20959 30923
rect 20901 30883 20959 30889
rect 21082 30880 21088 30932
rect 21140 30880 21146 30932
rect 21174 30880 21180 30932
rect 21232 30920 21238 30932
rect 21361 30923 21419 30929
rect 21361 30920 21373 30923
rect 21232 30892 21373 30920
rect 21232 30880 21238 30892
rect 21361 30889 21373 30892
rect 21407 30889 21419 30923
rect 21361 30883 21419 30889
rect 22557 30923 22615 30929
rect 22557 30889 22569 30923
rect 22603 30920 22615 30923
rect 22830 30920 22836 30932
rect 22603 30892 22836 30920
rect 22603 30889 22615 30892
rect 22557 30883 22615 30889
rect 22830 30880 22836 30892
rect 22888 30880 22894 30932
rect 25685 30923 25743 30929
rect 25685 30889 25697 30923
rect 25731 30920 25743 30923
rect 25866 30920 25872 30932
rect 25731 30892 25872 30920
rect 25731 30889 25743 30892
rect 25685 30883 25743 30889
rect 25866 30880 25872 30892
rect 25924 30880 25930 30932
rect 26050 30880 26056 30932
rect 26108 30880 26114 30932
rect 28994 30880 29000 30932
rect 29052 30920 29058 30932
rect 30006 30920 30012 30932
rect 29052 30892 30012 30920
rect 29052 30880 29058 30892
rect 30006 30880 30012 30892
rect 30064 30920 30070 30932
rect 32030 30920 32036 30932
rect 30064 30892 30512 30920
rect 30064 30880 30070 30892
rect 21100 30852 21128 30880
rect 20456 30824 21128 30852
rect 22649 30855 22707 30861
rect 22649 30821 22661 30855
rect 22695 30821 22707 30855
rect 23477 30855 23535 30861
rect 23477 30852 23489 30855
rect 22649 30815 22707 30821
rect 22756 30824 23489 30852
rect 22664 30784 22692 30815
rect 18739 30756 19840 30784
rect 22112 30756 22692 30784
rect 18739 30753 18751 30756
rect 18693 30747 18751 30753
rect 14921 30719 14979 30725
rect 14921 30716 14933 30719
rect 14200 30688 14933 30716
rect 14921 30685 14933 30688
rect 14967 30685 14979 30719
rect 14921 30679 14979 30685
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30685 15163 30719
rect 15105 30679 15163 30685
rect 15197 30719 15255 30725
rect 15197 30685 15209 30719
rect 15243 30685 15255 30719
rect 15197 30679 15255 30685
rect 15473 30719 15531 30725
rect 15473 30685 15485 30719
rect 15519 30716 15531 30719
rect 15654 30716 15660 30728
rect 15519 30688 15660 30716
rect 15519 30685 15531 30688
rect 15473 30679 15531 30685
rect 14090 30608 14096 30660
rect 14148 30608 14154 30660
rect 14642 30608 14648 30660
rect 14700 30648 14706 30660
rect 15120 30648 15148 30679
rect 15654 30676 15660 30688
rect 15712 30716 15718 30728
rect 15712 30688 17632 30716
rect 15712 30676 15718 30688
rect 14700 30620 15148 30648
rect 14700 30608 14706 30620
rect 16482 30608 16488 30660
rect 16540 30608 16546 30660
rect 17604 30648 17632 30688
rect 18322 30676 18328 30728
rect 18380 30676 18386 30728
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 18509 30719 18567 30725
rect 18509 30716 18521 30719
rect 18472 30688 18521 30716
rect 18472 30676 18478 30688
rect 18509 30685 18521 30688
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 18782 30676 18788 30728
rect 18840 30676 18846 30728
rect 18966 30676 18972 30728
rect 19024 30676 19030 30728
rect 19702 30676 19708 30728
rect 19760 30676 19766 30728
rect 20070 30726 20076 30728
rect 19904 30725 20076 30726
rect 19889 30719 20076 30725
rect 19889 30685 19901 30719
rect 19935 30698 20076 30719
rect 19935 30685 19947 30698
rect 19889 30679 19947 30685
rect 20070 30676 20076 30698
rect 20128 30676 20134 30728
rect 20254 30676 20260 30728
rect 20312 30676 20318 30728
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 18984 30648 19012 30676
rect 17604 30620 19012 30648
rect 19429 30651 19487 30657
rect 19429 30617 19441 30651
rect 19475 30648 19487 30651
rect 20272 30648 20300 30676
rect 19475 30620 20300 30648
rect 19475 30617 19487 30620
rect 19429 30611 19487 30617
rect 16500 30580 16528 30608
rect 13964 30552 16528 30580
rect 13964 30540 13970 30552
rect 20254 30540 20260 30592
rect 20312 30580 20318 30592
rect 20364 30580 20392 30679
rect 20530 30676 20536 30728
rect 20588 30676 20594 30728
rect 20806 30676 20812 30728
rect 20864 30676 20870 30728
rect 21085 30719 21143 30725
rect 21085 30685 21097 30719
rect 21131 30685 21143 30719
rect 21085 30679 21143 30685
rect 21100 30648 21128 30679
rect 21174 30676 21180 30728
rect 21232 30676 21238 30728
rect 21266 30676 21272 30728
rect 21324 30716 21330 30728
rect 21453 30719 21511 30725
rect 21453 30716 21465 30719
rect 21324 30688 21465 30716
rect 21324 30676 21330 30688
rect 21453 30685 21465 30688
rect 21499 30716 21511 30719
rect 21913 30719 21971 30725
rect 21913 30716 21925 30719
rect 21499 30688 21925 30716
rect 21499 30685 21511 30688
rect 21453 30679 21511 30685
rect 21913 30685 21925 30688
rect 21959 30685 21971 30719
rect 21913 30679 21971 30685
rect 22002 30676 22008 30728
rect 22060 30676 22066 30728
rect 22112 30725 22140 30756
rect 22097 30719 22155 30725
rect 22097 30685 22109 30719
rect 22143 30685 22155 30719
rect 22097 30679 22155 30685
rect 22373 30719 22431 30725
rect 22373 30685 22385 30719
rect 22419 30716 22431 30719
rect 22756 30716 22784 30824
rect 23477 30821 23489 30824
rect 23523 30821 23535 30855
rect 23477 30815 23535 30821
rect 23584 30824 24164 30852
rect 23293 30787 23351 30793
rect 23293 30753 23305 30787
rect 23339 30784 23351 30787
rect 23584 30784 23612 30824
rect 24136 30796 24164 30824
rect 23339 30756 23612 30784
rect 23339 30753 23351 30756
rect 23293 30747 23351 30753
rect 23308 30716 23336 30747
rect 23750 30744 23756 30796
rect 23808 30744 23814 30796
rect 24118 30744 24124 30796
rect 24176 30744 24182 30796
rect 26068 30784 26096 30880
rect 29270 30812 29276 30864
rect 29328 30812 29334 30864
rect 30484 30852 30512 30892
rect 30852 30892 32036 30920
rect 30852 30852 30880 30892
rect 32030 30880 32036 30892
rect 32088 30880 32094 30932
rect 34333 30923 34391 30929
rect 34333 30889 34345 30923
rect 34379 30920 34391 30923
rect 34422 30920 34428 30932
rect 34379 30892 34428 30920
rect 34379 30889 34391 30892
rect 34333 30883 34391 30889
rect 34422 30880 34428 30892
rect 34480 30880 34486 30932
rect 35986 30880 35992 30932
rect 36044 30920 36050 30932
rect 37277 30923 37335 30929
rect 37277 30920 37289 30923
rect 36044 30892 37289 30920
rect 36044 30880 36050 30892
rect 37277 30889 37289 30892
rect 37323 30889 37335 30923
rect 37277 30883 37335 30889
rect 38105 30923 38163 30929
rect 38105 30889 38117 30923
rect 38151 30920 38163 30923
rect 38378 30920 38384 30932
rect 38151 30892 38384 30920
rect 38151 30889 38163 30892
rect 38105 30883 38163 30889
rect 38378 30880 38384 30892
rect 38436 30880 38442 30932
rect 38746 30880 38752 30932
rect 38804 30920 38810 30932
rect 38933 30923 38991 30929
rect 38933 30920 38945 30923
rect 38804 30892 38945 30920
rect 38804 30880 38810 30892
rect 38933 30889 38945 30892
rect 38979 30889 38991 30923
rect 38933 30883 38991 30889
rect 40586 30880 40592 30932
rect 40644 30880 40650 30932
rect 41046 30880 41052 30932
rect 41104 30920 41110 30932
rect 41322 30920 41328 30932
rect 41104 30892 41328 30920
rect 41104 30880 41110 30892
rect 41322 30880 41328 30892
rect 41380 30920 41386 30932
rect 41785 30923 41843 30929
rect 41785 30920 41797 30923
rect 41380 30892 41797 30920
rect 41380 30880 41386 30892
rect 41785 30889 41797 30892
rect 41831 30889 41843 30923
rect 41785 30883 41843 30889
rect 42150 30880 42156 30932
rect 42208 30880 42214 30932
rect 30484 30824 30880 30852
rect 32968 30824 34376 30852
rect 27157 30787 27215 30793
rect 27157 30784 27169 30787
rect 26068 30756 27169 30784
rect 27157 30753 27169 30756
rect 27203 30753 27215 30787
rect 27157 30747 27215 30753
rect 27433 30787 27491 30793
rect 27433 30753 27445 30787
rect 27479 30784 27491 30787
rect 27525 30787 27583 30793
rect 27525 30784 27537 30787
rect 27479 30756 27537 30784
rect 27479 30753 27491 30756
rect 27433 30747 27491 30753
rect 27525 30753 27537 30756
rect 27571 30784 27583 30787
rect 28258 30784 28264 30796
rect 27571 30756 28264 30784
rect 27571 30753 27583 30756
rect 27525 30747 27583 30753
rect 28258 30744 28264 30756
rect 28316 30744 28322 30796
rect 29288 30784 29316 30812
rect 32968 30784 32996 30824
rect 29288 30756 32996 30784
rect 33045 30787 33103 30793
rect 33045 30753 33057 30787
rect 33091 30784 33103 30787
rect 33686 30784 33692 30796
rect 33091 30756 33692 30784
rect 33091 30753 33103 30756
rect 33045 30747 33103 30753
rect 33686 30744 33692 30756
rect 33744 30744 33750 30796
rect 33965 30787 34023 30793
rect 33965 30753 33977 30787
rect 34011 30784 34023 30787
rect 34238 30784 34244 30796
rect 34011 30756 34244 30784
rect 34011 30753 34023 30756
rect 33965 30747 34023 30753
rect 22419 30688 22784 30716
rect 22940 30688 23336 30716
rect 23768 30716 23796 30744
rect 23845 30719 23903 30725
rect 23845 30716 23857 30719
rect 23768 30688 23857 30716
rect 22419 30685 22431 30688
rect 22373 30679 22431 30685
rect 22940 30648 22968 30688
rect 23845 30685 23857 30688
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 23934 30676 23940 30728
rect 23992 30716 23998 30728
rect 24949 30719 25007 30725
rect 24949 30716 24961 30719
rect 23992 30688 24961 30716
rect 23992 30676 23998 30688
rect 24949 30685 24961 30688
rect 24995 30685 25007 30719
rect 24949 30679 25007 30685
rect 29454 30676 29460 30728
rect 29512 30716 29518 30728
rect 30193 30719 30251 30725
rect 30193 30716 30205 30719
rect 29512 30688 30205 30716
rect 29512 30676 29518 30688
rect 30193 30685 30205 30688
rect 30239 30685 30251 30719
rect 30193 30679 30251 30685
rect 30374 30676 30380 30728
rect 30432 30676 30438 30728
rect 31294 30676 31300 30728
rect 31352 30676 31358 30728
rect 33980 30716 34008 30747
rect 34238 30744 34244 30756
rect 34296 30744 34302 30796
rect 33244 30688 34008 30716
rect 34057 30719 34115 30725
rect 20824 30620 21128 30648
rect 22066 30620 22968 30648
rect 23017 30651 23075 30657
rect 20824 30592 20852 30620
rect 20312 30552 20392 30580
rect 20312 30540 20318 30552
rect 20806 30540 20812 30592
rect 20864 30540 20870 30592
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 22066 30580 22094 30620
rect 23017 30617 23029 30651
rect 23063 30648 23075 30651
rect 24397 30651 24455 30657
rect 24397 30648 24409 30651
rect 23063 30620 24409 30648
rect 23063 30617 23075 30620
rect 23017 30611 23075 30617
rect 24397 30617 24409 30620
rect 24443 30617 24455 30651
rect 24397 30611 24455 30617
rect 26694 30608 26700 30660
rect 26752 30648 26758 30660
rect 26752 30620 26832 30648
rect 26752 30608 26758 30620
rect 20956 30552 22094 30580
rect 22281 30583 22339 30589
rect 20956 30540 20962 30552
rect 22281 30549 22293 30583
rect 22327 30580 22339 30583
rect 22462 30580 22468 30592
rect 22327 30552 22468 30580
rect 22327 30549 22339 30552
rect 22281 30543 22339 30549
rect 22462 30540 22468 30552
rect 22520 30540 22526 30592
rect 23109 30583 23167 30589
rect 23109 30549 23121 30583
rect 23155 30580 23167 30583
rect 23382 30580 23388 30592
rect 23155 30552 23388 30580
rect 23155 30549 23167 30552
rect 23109 30543 23167 30549
rect 23382 30540 23388 30552
rect 23440 30540 23446 30592
rect 23937 30583 23995 30589
rect 23937 30549 23949 30583
rect 23983 30580 23995 30583
rect 26234 30580 26240 30592
rect 23983 30552 26240 30580
rect 23983 30549 23995 30552
rect 23937 30543 23995 30549
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 26804 30580 26832 30620
rect 27798 30608 27804 30660
rect 27856 30608 27862 30660
rect 30392 30648 30420 30676
rect 33244 30660 33272 30688
rect 34057 30685 34069 30719
rect 34103 30716 34115 30719
rect 34146 30716 34152 30728
rect 34103 30688 34152 30716
rect 34103 30685 34115 30688
rect 34057 30679 34115 30685
rect 34146 30676 34152 30688
rect 34204 30676 34210 30728
rect 27908 30620 28290 30648
rect 29104 30620 30420 30648
rect 31573 30651 31631 30657
rect 27908 30580 27936 30620
rect 29104 30592 29132 30620
rect 31573 30617 31585 30651
rect 31619 30648 31631 30651
rect 31846 30648 31852 30660
rect 31619 30620 31852 30648
rect 31619 30617 31631 30620
rect 31573 30611 31631 30617
rect 31846 30608 31852 30620
rect 31904 30608 31910 30660
rect 32030 30608 32036 30660
rect 32088 30608 32094 30660
rect 33226 30648 33232 30660
rect 33060 30620 33232 30648
rect 26804 30552 27936 30580
rect 29086 30540 29092 30592
rect 29144 30540 29150 30592
rect 31205 30583 31263 30589
rect 31205 30549 31217 30583
rect 31251 30580 31263 30583
rect 33060 30580 33088 30620
rect 33226 30608 33232 30620
rect 33284 30608 33290 30660
rect 34348 30648 34376 30824
rect 34440 30716 34468 30880
rect 36814 30812 36820 30864
rect 36872 30852 36878 30864
rect 36872 30824 40540 30852
rect 36872 30812 36878 30824
rect 34790 30744 34796 30796
rect 34848 30744 34854 30796
rect 38304 30756 39252 30784
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34440 30688 34897 30716
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35342 30676 35348 30728
rect 35400 30716 35406 30728
rect 35529 30719 35587 30725
rect 35529 30716 35541 30719
rect 35400 30688 35541 30716
rect 35400 30676 35406 30688
rect 35529 30685 35541 30688
rect 35575 30685 35587 30719
rect 35529 30679 35587 30685
rect 37918 30676 37924 30728
rect 37976 30676 37982 30728
rect 38194 30676 38200 30728
rect 38252 30676 38258 30728
rect 38304 30725 38332 30756
rect 38289 30719 38347 30725
rect 38289 30685 38301 30719
rect 38335 30685 38347 30719
rect 38289 30679 38347 30685
rect 38657 30719 38715 30725
rect 38657 30685 38669 30719
rect 38703 30716 38715 30719
rect 38746 30716 38752 30728
rect 38703 30688 38752 30716
rect 38703 30685 38715 30688
rect 38657 30679 38715 30685
rect 38746 30676 38752 30688
rect 38804 30716 38810 30728
rect 39117 30719 39175 30725
rect 39117 30716 39129 30719
rect 38804 30688 39129 30716
rect 38804 30676 38810 30688
rect 39117 30685 39129 30688
rect 39163 30685 39175 30719
rect 39117 30679 39175 30685
rect 34348 30620 35388 30648
rect 31251 30552 33088 30580
rect 31251 30549 31263 30552
rect 31205 30543 31263 30549
rect 33134 30540 33140 30592
rect 33192 30540 33198 30592
rect 35250 30540 35256 30592
rect 35308 30540 35314 30592
rect 35360 30580 35388 30620
rect 35710 30608 35716 30660
rect 35768 30648 35774 30660
rect 35805 30651 35863 30657
rect 35805 30648 35817 30651
rect 35768 30620 35817 30648
rect 35768 30608 35774 30620
rect 35805 30617 35817 30620
rect 35851 30617 35863 30651
rect 37030 30620 37780 30648
rect 35805 30611 35863 30617
rect 36446 30580 36452 30592
rect 35360 30552 36452 30580
rect 36446 30540 36452 30552
rect 36504 30540 36510 30592
rect 37752 30580 37780 30620
rect 38010 30608 38016 30660
rect 38068 30648 38074 30660
rect 38473 30651 38531 30657
rect 38473 30648 38485 30651
rect 38068 30620 38485 30648
rect 38068 30608 38074 30620
rect 38473 30617 38485 30620
rect 38519 30617 38531 30651
rect 38473 30611 38531 30617
rect 38562 30608 38568 30660
rect 38620 30608 38626 30660
rect 39224 30657 39252 30756
rect 40512 30728 40540 30824
rect 41138 30744 41144 30796
rect 41196 30744 41202 30796
rect 42168 30784 42196 30880
rect 42337 30787 42395 30793
rect 42337 30784 42349 30787
rect 42168 30756 42349 30784
rect 42337 30753 42349 30756
rect 42383 30753 42395 30787
rect 42337 30747 42395 30753
rect 42794 30744 42800 30796
rect 42852 30784 42858 30796
rect 43346 30784 43352 30796
rect 42852 30756 43352 30784
rect 42852 30744 42858 30756
rect 43346 30744 43352 30756
rect 43404 30784 43410 30796
rect 44085 30787 44143 30793
rect 44085 30784 44097 30787
rect 43404 30756 44097 30784
rect 43404 30744 43410 30756
rect 44085 30753 44097 30756
rect 44131 30753 44143 30787
rect 44085 30747 44143 30753
rect 39482 30676 39488 30728
rect 39540 30676 39546 30728
rect 39758 30676 39764 30728
rect 39816 30716 39822 30728
rect 40405 30719 40463 30725
rect 40405 30716 40417 30719
rect 39816 30688 40417 30716
rect 39816 30676 39822 30688
rect 40405 30685 40417 30688
rect 40451 30685 40463 30719
rect 40405 30679 40463 30685
rect 39209 30651 39267 30657
rect 38764 30620 39160 30648
rect 38764 30580 38792 30620
rect 39132 30592 39160 30620
rect 39209 30617 39221 30651
rect 39255 30617 39267 30651
rect 39209 30611 39267 30617
rect 37752 30552 38792 30580
rect 38838 30540 38844 30592
rect 38896 30540 38902 30592
rect 39114 30540 39120 30592
rect 39172 30540 39178 30592
rect 39224 30580 39252 30611
rect 39298 30608 39304 30660
rect 39356 30608 39362 30660
rect 40420 30648 40448 30679
rect 40494 30676 40500 30728
rect 40552 30676 40558 30728
rect 40770 30676 40776 30728
rect 40828 30716 40834 30728
rect 41509 30719 41567 30725
rect 41509 30716 41521 30719
rect 40828 30688 41521 30716
rect 40828 30676 40834 30688
rect 41509 30685 41521 30688
rect 41555 30685 41567 30719
rect 41509 30679 41567 30685
rect 41601 30719 41659 30725
rect 41601 30685 41613 30719
rect 41647 30685 41659 30719
rect 41601 30679 41659 30685
rect 41877 30719 41935 30725
rect 41877 30685 41889 30719
rect 41923 30685 41935 30719
rect 41877 30679 41935 30685
rect 41616 30648 41644 30679
rect 40420 30620 41644 30648
rect 41892 30648 41920 30679
rect 41966 30676 41972 30728
rect 42024 30716 42030 30728
rect 42061 30719 42119 30725
rect 42061 30716 42073 30719
rect 42024 30688 42073 30716
rect 42024 30676 42030 30688
rect 42061 30685 42073 30688
rect 42107 30685 42119 30719
rect 42061 30679 42119 30685
rect 43438 30676 43444 30728
rect 43496 30676 43502 30728
rect 41892 30620 42748 30648
rect 39853 30583 39911 30589
rect 39853 30580 39865 30583
rect 39224 30552 39865 30580
rect 39853 30549 39865 30552
rect 39899 30549 39911 30583
rect 39853 30543 39911 30549
rect 41325 30583 41383 30589
rect 41325 30549 41337 30583
rect 41371 30580 41383 30583
rect 41874 30580 41880 30592
rect 41371 30552 41880 30580
rect 41371 30549 41383 30552
rect 41325 30543 41383 30549
rect 41874 30540 41880 30552
rect 41932 30540 41938 30592
rect 42720 30580 42748 30620
rect 43070 30580 43076 30592
rect 42720 30552 43076 30580
rect 43070 30540 43076 30552
rect 43128 30540 43134 30592
rect 1104 30490 44620 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 44620 30490
rect 1104 30416 44620 30438
rect 5626 30336 5632 30388
rect 5684 30336 5690 30388
rect 6086 30336 6092 30388
rect 6144 30336 6150 30388
rect 7374 30336 7380 30388
rect 7432 30336 7438 30388
rect 7558 30336 7564 30388
rect 7616 30336 7622 30388
rect 7834 30336 7840 30388
rect 7892 30376 7898 30388
rect 9493 30379 9551 30385
rect 9493 30376 9505 30379
rect 7892 30348 9505 30376
rect 7892 30336 7898 30348
rect 9493 30345 9505 30348
rect 9539 30345 9551 30379
rect 9493 30339 9551 30345
rect 11977 30379 12035 30385
rect 11977 30345 11989 30379
rect 12023 30376 12035 30379
rect 12066 30376 12072 30388
rect 12023 30348 12072 30376
rect 12023 30345 12035 30348
rect 11977 30339 12035 30345
rect 5721 30311 5779 30317
rect 5721 30277 5733 30311
rect 5767 30277 5779 30311
rect 5721 30271 5779 30277
rect 5951 30277 6009 30283
rect 5951 30274 5963 30277
rect 5353 30243 5411 30249
rect 5353 30209 5365 30243
rect 5399 30240 5411 30243
rect 5399 30212 5580 30240
rect 5399 30209 5411 30212
rect 5353 30203 5411 30209
rect 5442 29996 5448 30048
rect 5500 29996 5506 30048
rect 5552 30036 5580 30212
rect 5736 30184 5764 30271
rect 5936 30243 5963 30274
rect 5997 30243 6009 30277
rect 5936 30240 6009 30243
rect 7469 30243 7527 30249
rect 5936 30212 6040 30240
rect 6012 30184 6040 30212
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 7576 30240 7604 30336
rect 9508 30308 9536 30339
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 12894 30376 12900 30388
rect 12268 30348 12900 30376
rect 12158 30308 12164 30320
rect 9508 30280 12164 30308
rect 9306 30240 9312 30252
rect 7515 30212 7604 30240
rect 9154 30212 9312 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 9306 30200 9312 30212
rect 9364 30240 9370 30252
rect 9490 30240 9496 30252
rect 9364 30212 9496 30240
rect 9364 30200 9370 30212
rect 9490 30200 9496 30212
rect 9548 30200 9554 30252
rect 10796 30249 10824 30280
rect 12158 30268 12164 30280
rect 12216 30268 12222 30320
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30209 10839 30243
rect 10781 30203 10839 30209
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 12268 30240 12296 30348
rect 12894 30336 12900 30348
rect 12952 30376 12958 30388
rect 13630 30376 13636 30388
rect 12952 30348 13636 30376
rect 12952 30336 12958 30348
rect 13630 30336 13636 30348
rect 13688 30336 13694 30388
rect 13722 30336 13728 30388
rect 13780 30376 13786 30388
rect 13780 30348 13952 30376
rect 13780 30336 13786 30348
rect 12437 30311 12495 30317
rect 12437 30277 12449 30311
rect 12483 30308 12495 30311
rect 13170 30308 13176 30320
rect 12483 30280 13032 30308
rect 12483 30277 12495 30280
rect 12437 30271 12495 30277
rect 11931 30212 12296 30240
rect 12529 30243 12587 30249
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 12529 30209 12541 30243
rect 12575 30240 12587 30243
rect 12710 30241 12716 30252
rect 12636 30240 12716 30241
rect 12575 30213 12716 30240
rect 12575 30212 12664 30213
rect 12575 30209 12587 30212
rect 12529 30203 12587 30209
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30141 5687 30175
rect 5629 30135 5687 30141
rect 5644 30104 5672 30135
rect 5718 30132 5724 30184
rect 5776 30132 5782 30184
rect 5994 30132 6000 30184
rect 6052 30132 6058 30184
rect 6914 30132 6920 30184
rect 6972 30172 6978 30184
rect 7745 30175 7803 30181
rect 7745 30172 7757 30175
rect 6972 30144 7757 30172
rect 6972 30132 6978 30144
rect 7745 30141 7757 30144
rect 7791 30141 7803 30175
rect 7745 30135 7803 30141
rect 8018 30132 8024 30184
rect 8076 30132 8082 30184
rect 7558 30104 7564 30116
rect 5644 30076 7564 30104
rect 7558 30064 7564 30076
rect 7616 30064 7622 30116
rect 11900 30104 11928 30203
rect 12710 30200 12716 30213
rect 12768 30200 12774 30252
rect 12820 30249 12848 30280
rect 13004 30252 13032 30280
rect 13096 30280 13176 30308
rect 12805 30243 12863 30249
rect 12805 30209 12817 30243
rect 12851 30209 12863 30243
rect 12805 30203 12863 30209
rect 12897 30243 12955 30249
rect 12897 30209 12909 30243
rect 12943 30209 12955 30243
rect 12897 30203 12955 30209
rect 12250 30132 12256 30184
rect 12308 30132 12314 30184
rect 12912 30172 12940 30203
rect 12986 30200 12992 30252
rect 13044 30200 13050 30252
rect 13096 30172 13124 30280
rect 13170 30268 13176 30280
rect 13228 30268 13234 30320
rect 13924 30317 13952 30348
rect 18782 30336 18788 30388
rect 18840 30336 18846 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19484 30348 20300 30376
rect 19484 30336 19490 30348
rect 13909 30311 13967 30317
rect 13909 30277 13921 30311
rect 13955 30277 13967 30311
rect 13909 30271 13967 30277
rect 15194 30268 15200 30320
rect 15252 30268 15258 30320
rect 18414 30268 18420 30320
rect 18472 30308 18478 30320
rect 18800 30308 18828 30336
rect 18472 30280 18736 30308
rect 18800 30280 19196 30308
rect 18472 30268 18478 30280
rect 13633 30243 13691 30249
rect 13633 30240 13645 30243
rect 13188 30212 13645 30240
rect 13188 30181 13216 30212
rect 13633 30209 13645 30212
rect 13679 30209 13691 30243
rect 15105 30243 15163 30249
rect 15105 30240 15117 30243
rect 13633 30203 13691 30209
rect 13924 30212 15117 30240
rect 12544 30144 12848 30172
rect 12912 30144 13124 30172
rect 13173 30175 13231 30181
rect 9048 30076 11928 30104
rect 12268 30104 12296 30132
rect 12544 30104 12572 30144
rect 12268 30076 12572 30104
rect 5810 30036 5816 30048
rect 5552 30008 5816 30036
rect 5810 29996 5816 30008
rect 5868 30036 5874 30048
rect 5905 30039 5963 30045
rect 5905 30036 5917 30039
rect 5868 30008 5917 30036
rect 5868 29996 5874 30008
rect 5905 30005 5917 30008
rect 5951 30036 5963 30039
rect 9048 30036 9076 30076
rect 12618 30064 12624 30116
rect 12676 30064 12682 30116
rect 12820 30104 12848 30144
rect 13173 30141 13185 30175
rect 13219 30141 13231 30175
rect 13173 30135 13231 30141
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30172 13323 30175
rect 13541 30175 13599 30181
rect 13541 30172 13553 30175
rect 13311 30144 13553 30172
rect 13311 30141 13323 30144
rect 13265 30135 13323 30141
rect 13541 30141 13553 30144
rect 13587 30172 13599 30175
rect 13814 30172 13820 30184
rect 13587 30144 13820 30172
rect 13587 30141 13599 30144
rect 13541 30135 13599 30141
rect 13188 30104 13216 30135
rect 13814 30132 13820 30144
rect 13872 30132 13878 30184
rect 13924 30104 13952 30212
rect 15105 30209 15117 30212
rect 15151 30240 15163 30243
rect 15151 30212 15700 30240
rect 15151 30209 15163 30212
rect 15105 30203 15163 30209
rect 13998 30132 14004 30184
rect 14056 30172 14062 30184
rect 15562 30172 15568 30184
rect 14056 30144 15568 30172
rect 14056 30132 14062 30144
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 12820 30076 13216 30104
rect 13280 30076 13952 30104
rect 5951 30008 9076 30036
rect 10689 30039 10747 30045
rect 5951 30005 5963 30008
rect 5905 29999 5963 30005
rect 10689 30005 10701 30039
rect 10735 30036 10747 30039
rect 11606 30036 11612 30048
rect 10735 30008 11612 30036
rect 10735 30005 10747 30008
rect 10689 29999 10747 30005
rect 11606 29996 11612 30008
rect 11664 29996 11670 30048
rect 11882 29996 11888 30048
rect 11940 30036 11946 30048
rect 13280 30036 13308 30076
rect 11940 30008 13308 30036
rect 11940 29996 11946 30008
rect 13354 29996 13360 30048
rect 13412 29996 13418 30048
rect 15672 30036 15700 30212
rect 18046 30200 18052 30252
rect 18104 30200 18110 30252
rect 18322 30200 18328 30252
rect 18380 30240 18386 30252
rect 18708 30249 18736 30280
rect 18966 30249 18972 30252
rect 18509 30243 18567 30249
rect 18509 30240 18521 30243
rect 18380 30212 18521 30240
rect 18380 30200 18386 30212
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 16669 30175 16727 30181
rect 16669 30172 16681 30175
rect 16632 30144 16681 30172
rect 16632 30132 16638 30144
rect 16669 30141 16681 30144
rect 16715 30141 16727 30175
rect 16669 30135 16727 30141
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30172 17003 30175
rect 16991 30144 18092 30172
rect 16991 30141 17003 30144
rect 16945 30135 17003 30141
rect 18064 30116 18092 30144
rect 18046 30064 18052 30116
rect 18104 30064 18110 30116
rect 17310 30036 17316 30048
rect 15672 30008 17316 30036
rect 17310 29996 17316 30008
rect 17368 29996 17374 30048
rect 17954 29996 17960 30048
rect 18012 30036 18018 30048
rect 18432 30045 18460 30212
rect 18509 30209 18521 30212
rect 18555 30209 18567 30243
rect 18509 30203 18567 30209
rect 18693 30243 18751 30249
rect 18693 30209 18705 30243
rect 18739 30209 18751 30243
rect 18961 30240 18972 30249
rect 18927 30212 18972 30240
rect 18693 30203 18751 30209
rect 18961 30203 18972 30212
rect 18966 30200 18972 30203
rect 19024 30200 19030 30252
rect 19168 30249 19196 30280
rect 19153 30243 19211 30249
rect 19153 30209 19165 30243
rect 19199 30209 19211 30243
rect 19153 30203 19211 30209
rect 19334 30200 19340 30252
rect 19392 30200 19398 30252
rect 19444 30240 19472 30336
rect 20162 30308 20168 30320
rect 19904 30280 20168 30308
rect 19613 30243 19671 30249
rect 19613 30240 19625 30243
rect 19444 30212 19625 30240
rect 19613 30209 19625 30212
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 19794 30200 19800 30252
rect 19852 30200 19858 30252
rect 19904 30249 19932 30280
rect 20162 30268 20168 30280
rect 20220 30268 20226 30320
rect 20272 30317 20300 30348
rect 20438 30336 20444 30388
rect 20496 30376 20502 30388
rect 20533 30379 20591 30385
rect 20533 30376 20545 30379
rect 20496 30348 20545 30376
rect 20496 30336 20502 30348
rect 20533 30345 20545 30348
rect 20579 30345 20591 30379
rect 20533 30339 20591 30345
rect 22002 30336 22008 30388
rect 22060 30376 22066 30388
rect 23934 30376 23940 30388
rect 22060 30348 22232 30376
rect 22060 30336 22066 30348
rect 20257 30311 20315 30317
rect 20257 30277 20269 30311
rect 20303 30277 20315 30311
rect 22204 30308 22232 30348
rect 22572 30348 23940 30376
rect 22572 30308 22600 30348
rect 23934 30336 23940 30348
rect 23992 30336 23998 30388
rect 26694 30376 26700 30388
rect 26160 30348 26700 30376
rect 26160 30308 26188 30348
rect 26694 30336 26700 30348
rect 26752 30336 26758 30388
rect 27430 30336 27436 30388
rect 27488 30336 27494 30388
rect 27617 30379 27675 30385
rect 27617 30345 27629 30379
rect 27663 30376 27675 30379
rect 27798 30376 27804 30388
rect 27663 30348 27804 30376
rect 27663 30345 27675 30348
rect 27617 30339 27675 30345
rect 27798 30336 27804 30348
rect 27856 30336 27862 30388
rect 30098 30376 30104 30388
rect 28966 30348 30104 30376
rect 22204 30280 22600 30308
rect 25622 30280 26188 30308
rect 20257 30271 20315 30277
rect 26418 30268 26424 30320
rect 26476 30308 26482 30320
rect 27249 30311 27307 30317
rect 27249 30308 27261 30311
rect 26476 30280 27261 30308
rect 26476 30268 26482 30280
rect 27249 30277 27261 30280
rect 27295 30277 27307 30311
rect 27249 30271 27307 30277
rect 27341 30311 27399 30317
rect 27341 30277 27353 30311
rect 27387 30308 27399 30311
rect 27448 30308 27476 30336
rect 27387 30280 27476 30308
rect 27387 30277 27399 30280
rect 27341 30271 27399 30277
rect 27522 30268 27528 30320
rect 27580 30308 27586 30320
rect 28966 30308 28994 30348
rect 30098 30336 30104 30348
rect 30156 30376 30162 30388
rect 30156 30348 30696 30376
rect 30156 30336 30162 30348
rect 27580 30280 28994 30308
rect 27580 30268 27586 30280
rect 29086 30268 29092 30320
rect 29144 30308 29150 30320
rect 29144 30280 29408 30308
rect 29144 30268 29150 30280
rect 19889 30243 19947 30249
rect 19889 30209 19901 30243
rect 19935 30209 19947 30243
rect 19889 30203 19947 30209
rect 20346 30200 20352 30252
rect 20404 30249 20410 30252
rect 20404 30243 20432 30249
rect 20420 30209 20432 30243
rect 20898 30240 20904 30252
rect 20404 30203 20432 30209
rect 20548 30212 20904 30240
rect 20404 30200 20410 30203
rect 19426 30132 19432 30184
rect 19484 30132 19490 30184
rect 19521 30175 19579 30181
rect 19521 30141 19533 30175
rect 19567 30172 19579 30175
rect 19812 30172 19840 30200
rect 19567 30144 19840 30172
rect 20165 30175 20223 30181
rect 19567 30141 19579 30144
rect 19521 30135 19579 30141
rect 19061 30107 19119 30113
rect 19061 30073 19073 30107
rect 19107 30104 19119 30107
rect 19628 30104 19656 30144
rect 20165 30141 20177 30175
rect 20211 30141 20223 30175
rect 20165 30135 20223 30141
rect 19107 30076 19656 30104
rect 19797 30107 19855 30113
rect 19107 30073 19119 30076
rect 19061 30067 19119 30073
rect 19797 30073 19809 30107
rect 19843 30104 19855 30107
rect 19978 30104 19984 30116
rect 19843 30076 19984 30104
rect 19843 30073 19855 30076
rect 19797 30067 19855 30073
rect 19978 30064 19984 30076
rect 20036 30064 20042 30116
rect 20180 30104 20208 30135
rect 20548 30104 20576 30212
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 21082 30200 21088 30252
rect 21140 30200 21146 30252
rect 23566 30200 23572 30252
rect 23624 30200 23630 30252
rect 26973 30243 27031 30249
rect 26973 30209 26985 30243
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27121 30243 27179 30249
rect 27121 30209 27133 30243
rect 27167 30240 27179 30243
rect 27438 30243 27496 30249
rect 27167 30212 27384 30240
rect 27167 30209 27179 30212
rect 27121 30203 27179 30209
rect 20622 30132 20628 30184
rect 20680 30172 20686 30184
rect 20806 30172 20812 30184
rect 20680 30144 20812 30172
rect 20680 30132 20686 30144
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 20990 30132 20996 30184
rect 21048 30132 21054 30184
rect 22189 30175 22247 30181
rect 22189 30141 22201 30175
rect 22235 30141 22247 30175
rect 22189 30135 22247 30141
rect 20180 30076 20576 30104
rect 18417 30039 18475 30045
rect 18417 30036 18429 30039
rect 18012 30008 18429 30036
rect 18012 29996 18018 30008
rect 18417 30005 18429 30008
rect 18463 30005 18475 30039
rect 18417 29999 18475 30005
rect 18598 29996 18604 30048
rect 18656 29996 18662 30048
rect 19426 29996 19432 30048
rect 19484 30036 19490 30048
rect 20625 30039 20683 30045
rect 20625 30036 20637 30039
rect 19484 30008 20637 30036
rect 19484 29996 19490 30008
rect 20625 30005 20637 30008
rect 20671 30005 20683 30039
rect 22204 30036 22232 30135
rect 22462 30132 22468 30184
rect 22520 30132 22526 30184
rect 24121 30175 24179 30181
rect 24121 30172 24133 30175
rect 23584 30144 24133 30172
rect 23584 30116 23612 30144
rect 24121 30141 24133 30144
rect 24167 30141 24179 30175
rect 24121 30135 24179 30141
rect 24394 30132 24400 30184
rect 24452 30132 24458 30184
rect 24486 30132 24492 30184
rect 24544 30172 24550 30184
rect 25869 30175 25927 30181
rect 25869 30172 25881 30175
rect 24544 30144 25881 30172
rect 24544 30132 24550 30144
rect 25869 30141 25881 30144
rect 25915 30141 25927 30175
rect 25869 30135 25927 30141
rect 26418 30132 26424 30184
rect 26476 30172 26482 30184
rect 26988 30172 27016 30203
rect 26476 30144 27016 30172
rect 27356 30172 27384 30212
rect 27438 30209 27450 30243
rect 27484 30240 27496 30243
rect 27540 30240 27568 30268
rect 27484 30212 27568 30240
rect 27484 30209 27496 30212
rect 27438 30203 27496 30209
rect 27890 30200 27896 30252
rect 27948 30240 27954 30252
rect 29273 30243 29331 30249
rect 27948 30212 29132 30240
rect 27948 30200 27954 30212
rect 28994 30172 29000 30184
rect 27356 30144 29000 30172
rect 26476 30132 26482 30144
rect 28994 30132 29000 30144
rect 29052 30132 29058 30184
rect 29104 30181 29132 30212
rect 29273 30209 29285 30243
rect 29319 30209 29331 30243
rect 29380 30240 29408 30280
rect 29454 30268 29460 30320
rect 29512 30268 29518 30320
rect 29549 30243 29607 30249
rect 29380 30238 29500 30240
rect 29549 30238 29561 30243
rect 29380 30212 29561 30238
rect 29472 30210 29561 30212
rect 29273 30203 29331 30209
rect 29549 30209 29561 30210
rect 29595 30209 29607 30243
rect 29549 30203 29607 30209
rect 29089 30175 29147 30181
rect 29089 30141 29101 30175
rect 29135 30172 29147 30175
rect 29178 30172 29184 30184
rect 29135 30144 29184 30172
rect 29135 30141 29147 30144
rect 29089 30135 29147 30141
rect 29178 30132 29184 30144
rect 29236 30132 29242 30184
rect 29288 30172 29316 30203
rect 29638 30200 29644 30252
rect 29696 30200 29702 30252
rect 30009 30243 30067 30249
rect 30009 30209 30021 30243
rect 30055 30240 30067 30243
rect 30190 30240 30196 30252
rect 30055 30212 30196 30240
rect 30055 30209 30067 30212
rect 30009 30203 30067 30209
rect 30190 30200 30196 30212
rect 30248 30200 30254 30252
rect 29656 30172 29684 30200
rect 29288 30144 29684 30172
rect 23566 30064 23572 30116
rect 23624 30064 23630 30116
rect 29288 30104 29316 30144
rect 29730 30132 29736 30184
rect 29788 30172 29794 30184
rect 29825 30175 29883 30181
rect 29825 30172 29837 30175
rect 29788 30144 29837 30172
rect 29788 30132 29794 30144
rect 29825 30141 29837 30144
rect 29871 30141 29883 30175
rect 30668 30172 30696 30348
rect 31846 30336 31852 30388
rect 31904 30376 31910 30388
rect 32674 30376 32680 30388
rect 31904 30348 32260 30376
rect 31904 30336 31910 30348
rect 32232 30317 32260 30348
rect 32416 30348 32680 30376
rect 32217 30311 32275 30317
rect 32217 30277 32229 30311
rect 32263 30277 32275 30311
rect 32217 30271 32275 30277
rect 32416 30249 32444 30348
rect 32674 30336 32680 30348
rect 32732 30336 32738 30388
rect 32766 30336 32772 30388
rect 32824 30336 32830 30388
rect 33134 30336 33140 30388
rect 33192 30336 33198 30388
rect 33318 30385 33324 30388
rect 33314 30339 33324 30385
rect 33318 30336 33324 30339
rect 33376 30336 33382 30388
rect 34701 30379 34759 30385
rect 34072 30348 34560 30376
rect 32493 30311 32551 30317
rect 32493 30277 32505 30311
rect 32539 30308 32551 30311
rect 32784 30308 32812 30336
rect 33152 30308 33180 30336
rect 32539 30280 32812 30308
rect 32876 30280 33180 30308
rect 33413 30311 33471 30317
rect 32539 30277 32551 30280
rect 32493 30271 32551 30277
rect 32401 30243 32459 30249
rect 32401 30209 32413 30243
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 32582 30200 32588 30252
rect 32640 30200 32646 30252
rect 32876 30249 32904 30280
rect 33413 30277 33425 30311
rect 33459 30308 33471 30311
rect 33873 30311 33931 30317
rect 33873 30308 33885 30311
rect 33459 30280 33885 30308
rect 33459 30277 33471 30280
rect 33413 30271 33471 30277
rect 33873 30277 33885 30280
rect 33919 30277 33931 30311
rect 33873 30271 33931 30277
rect 34072 30252 34100 30348
rect 34532 30308 34560 30348
rect 34701 30345 34713 30379
rect 34747 30376 34759 30379
rect 34790 30376 34796 30388
rect 34747 30348 34796 30376
rect 34747 30345 34759 30348
rect 34701 30339 34759 30345
rect 34790 30336 34796 30348
rect 34848 30336 34854 30388
rect 35250 30336 35256 30388
rect 35308 30336 35314 30388
rect 35621 30379 35679 30385
rect 35621 30345 35633 30379
rect 35667 30376 35679 30379
rect 35710 30376 35716 30388
rect 35667 30348 35716 30376
rect 35667 30345 35679 30348
rect 35621 30339 35679 30345
rect 35710 30336 35716 30348
rect 35768 30336 35774 30388
rect 36722 30336 36728 30388
rect 36780 30336 36786 30388
rect 38194 30336 38200 30388
rect 38252 30376 38258 30388
rect 38289 30379 38347 30385
rect 38289 30376 38301 30379
rect 38252 30348 38301 30376
rect 38252 30336 38258 30348
rect 38289 30345 38301 30348
rect 38335 30345 38347 30379
rect 38289 30339 38347 30345
rect 38470 30336 38476 30388
rect 38528 30376 38534 30388
rect 38528 30348 38792 30376
rect 38528 30336 38534 30348
rect 35268 30308 35296 30336
rect 36740 30308 36768 30336
rect 34532 30280 34744 30308
rect 32723 30243 32781 30249
rect 32723 30240 32735 30243
rect 32718 30209 32735 30240
rect 32769 30209 32781 30243
rect 32718 30203 32781 30209
rect 32861 30243 32919 30249
rect 32861 30209 32873 30243
rect 32907 30209 32919 30243
rect 32861 30203 32919 30209
rect 32718 30172 32746 30203
rect 33134 30200 33140 30252
rect 33192 30200 33198 30252
rect 33229 30243 33287 30249
rect 33229 30209 33241 30243
rect 33275 30240 33287 30243
rect 33275 30212 33640 30240
rect 33275 30209 33287 30212
rect 33229 30203 33287 30209
rect 33612 30181 33640 30212
rect 33686 30200 33692 30252
rect 33744 30200 33750 30252
rect 34054 30200 34060 30252
rect 34112 30200 34118 30252
rect 34238 30200 34244 30252
rect 34296 30200 34302 30252
rect 34422 30200 34428 30252
rect 34480 30200 34486 30252
rect 30668 30144 32746 30172
rect 33597 30175 33655 30181
rect 29825 30135 29883 30141
rect 33597 30141 33609 30175
rect 33643 30172 33655 30175
rect 34146 30172 34152 30184
rect 33643 30144 34152 30172
rect 33643 30141 33655 30144
rect 33597 30135 33655 30141
rect 34146 30132 34152 30144
rect 34204 30172 34210 30184
rect 34716 30181 34744 30280
rect 35084 30280 35296 30308
rect 35452 30280 36768 30308
rect 35084 30249 35112 30280
rect 35452 30252 35480 30280
rect 35069 30243 35127 30249
rect 35069 30209 35081 30243
rect 35115 30209 35127 30243
rect 35069 30203 35127 30209
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30209 35311 30243
rect 35253 30203 35311 30209
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30209 35403 30243
rect 35345 30203 35403 30209
rect 34333 30175 34391 30181
rect 34333 30172 34345 30175
rect 34204 30144 34345 30172
rect 34204 30132 34210 30144
rect 34333 30141 34345 30144
rect 34379 30141 34391 30175
rect 34333 30135 34391 30141
rect 34701 30175 34759 30181
rect 34701 30141 34713 30175
rect 34747 30141 34759 30175
rect 34701 30135 34759 30141
rect 35268 30104 35296 30203
rect 35360 30172 35388 30203
rect 35434 30200 35440 30252
rect 35492 30200 35498 30252
rect 35986 30200 35992 30252
rect 36044 30240 36050 30252
rect 36265 30243 36323 30249
rect 36265 30240 36277 30243
rect 36044 30212 36277 30240
rect 36044 30200 36050 30212
rect 36265 30209 36277 30212
rect 36311 30209 36323 30243
rect 36265 30203 36323 30209
rect 36446 30200 36452 30252
rect 36504 30200 36510 30252
rect 36538 30200 36544 30252
rect 36596 30200 36602 30252
rect 37826 30200 37832 30252
rect 37884 30200 37890 30252
rect 38764 30249 38792 30348
rect 38838 30336 38844 30388
rect 38896 30376 38902 30388
rect 38896 30348 39068 30376
rect 38896 30336 38902 30348
rect 39040 30317 39068 30348
rect 40494 30336 40500 30388
rect 40552 30376 40558 30388
rect 40552 30348 42748 30376
rect 40552 30336 40558 30348
rect 39025 30311 39083 30317
rect 39025 30277 39037 30311
rect 39071 30277 39083 30311
rect 39025 30271 39083 30277
rect 39114 30268 39120 30320
rect 39172 30308 39178 30320
rect 39172 30280 39514 30308
rect 39172 30268 39178 30280
rect 38105 30243 38163 30249
rect 38105 30209 38117 30243
rect 38151 30209 38163 30243
rect 38105 30203 38163 30209
rect 38749 30243 38807 30249
rect 38749 30209 38761 30243
rect 38795 30209 38807 30243
rect 38749 30203 38807 30209
rect 35713 30175 35771 30181
rect 35713 30172 35725 30175
rect 35360 30144 35725 30172
rect 35713 30141 35725 30144
rect 35759 30141 35771 30175
rect 35713 30135 35771 30141
rect 36556 30104 36584 30200
rect 36722 30132 36728 30184
rect 36780 30132 36786 30184
rect 37921 30175 37979 30181
rect 37921 30172 37933 30175
rect 37016 30144 37933 30172
rect 37016 30113 37044 30144
rect 37921 30141 37933 30144
rect 37967 30141 37979 30175
rect 38120 30172 38148 30203
rect 41874 30200 41880 30252
rect 41932 30200 41938 30252
rect 42720 30240 42748 30348
rect 43070 30336 43076 30388
rect 43128 30336 43134 30388
rect 43162 30240 43168 30252
rect 42720 30212 43168 30240
rect 43162 30200 43168 30212
rect 43220 30200 43226 30252
rect 39758 30172 39764 30184
rect 38120 30144 39764 30172
rect 37921 30135 37979 30141
rect 39758 30132 39764 30144
rect 39816 30132 39822 30184
rect 41138 30132 41144 30184
rect 41196 30132 41202 30184
rect 42518 30132 42524 30184
rect 42576 30132 42582 30184
rect 27632 30076 29316 30104
rect 33428 30076 36584 30104
rect 37001 30107 37059 30113
rect 22554 30036 22560 30048
rect 22204 30008 22560 30036
rect 20625 29999 20683 30005
rect 22554 29996 22560 30008
rect 22612 30036 22618 30048
rect 23198 30036 23204 30048
rect 22612 30008 23204 30036
rect 22612 29996 22618 30008
rect 23198 29996 23204 30008
rect 23256 30036 23262 30048
rect 23584 30036 23612 30064
rect 27632 30048 27660 30076
rect 23256 30008 23612 30036
rect 23256 29996 23262 30008
rect 27614 29996 27620 30048
rect 27672 29996 27678 30048
rect 32858 29996 32864 30048
rect 32916 30036 32922 30048
rect 33428 30036 33456 30076
rect 37001 30073 37013 30107
rect 37047 30073 37059 30107
rect 37001 30067 37059 30073
rect 38010 30064 38016 30116
rect 38068 30104 38074 30116
rect 40497 30107 40555 30113
rect 38068 30076 38608 30104
rect 38068 30064 38074 30076
rect 32916 30008 33456 30036
rect 32916 29996 32922 30008
rect 33502 29996 33508 30048
rect 33560 30036 33566 30048
rect 34517 30039 34575 30045
rect 34517 30036 34529 30039
rect 33560 30008 34529 30036
rect 33560 29996 33566 30008
rect 34517 30005 34529 30008
rect 34563 30005 34575 30039
rect 34517 29999 34575 30005
rect 36817 30039 36875 30045
rect 36817 30005 36829 30039
rect 36863 30036 36875 30039
rect 36906 30036 36912 30048
rect 36863 30008 36912 30036
rect 36863 30005 36875 30008
rect 36817 29999 36875 30005
rect 36906 29996 36912 30008
rect 36964 29996 36970 30048
rect 38102 29996 38108 30048
rect 38160 29996 38166 30048
rect 38580 30036 38608 30076
rect 40497 30073 40509 30107
rect 40543 30104 40555 30107
rect 40543 30076 41092 30104
rect 40543 30073 40555 30076
rect 40497 30067 40555 30073
rect 41064 30048 41092 30076
rect 39206 30036 39212 30048
rect 38580 30008 39212 30036
rect 39206 29996 39212 30008
rect 39264 29996 39270 30048
rect 40586 29996 40592 30048
rect 40644 29996 40650 30048
rect 41046 29996 41052 30048
rect 41104 29996 41110 30048
rect 41230 29996 41236 30048
rect 41288 30036 41294 30048
rect 41325 30039 41383 30045
rect 41325 30036 41337 30039
rect 41288 30008 41337 30036
rect 41288 29996 41294 30008
rect 41325 30005 41337 30008
rect 41371 30005 41383 30039
rect 41325 29999 41383 30005
rect 1104 29946 44620 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 44620 29946
rect 1104 29872 44620 29894
rect 3878 29792 3884 29844
rect 3936 29792 3942 29844
rect 5442 29792 5448 29844
rect 5500 29832 5506 29844
rect 5721 29835 5779 29841
rect 5721 29832 5733 29835
rect 5500 29804 5733 29832
rect 5500 29792 5506 29804
rect 5721 29801 5733 29804
rect 5767 29801 5779 29835
rect 5721 29795 5779 29801
rect 7926 29792 7932 29844
rect 7984 29792 7990 29844
rect 8018 29792 8024 29844
rect 8076 29832 8082 29844
rect 8205 29835 8263 29841
rect 8205 29832 8217 29835
rect 8076 29804 8217 29832
rect 8076 29792 8082 29804
rect 8205 29801 8217 29804
rect 8251 29801 8263 29835
rect 8205 29795 8263 29801
rect 12526 29792 12532 29844
rect 12584 29832 12590 29844
rect 12621 29835 12679 29841
rect 12621 29832 12633 29835
rect 12584 29804 12633 29832
rect 12584 29792 12590 29804
rect 12621 29801 12633 29804
rect 12667 29801 12679 29835
rect 12621 29795 12679 29801
rect 13354 29792 13360 29844
rect 13412 29792 13418 29844
rect 13814 29792 13820 29844
rect 13872 29832 13878 29844
rect 13872 29804 17080 29832
rect 13872 29792 13878 29804
rect 3789 29699 3847 29705
rect 3789 29665 3801 29699
rect 3835 29696 3847 29699
rect 3896 29696 3924 29792
rect 3835 29668 3924 29696
rect 3835 29665 3847 29668
rect 3789 29659 3847 29665
rect 5994 29656 6000 29708
rect 6052 29696 6058 29708
rect 7944 29696 7972 29792
rect 10410 29724 10416 29776
rect 10468 29764 10474 29776
rect 11333 29767 11391 29773
rect 11333 29764 11345 29767
rect 10468 29736 11345 29764
rect 10468 29724 10474 29736
rect 11333 29733 11345 29736
rect 11379 29764 11391 29767
rect 12161 29767 12219 29773
rect 11379 29736 12020 29764
rect 11379 29733 11391 29736
rect 11333 29727 11391 29733
rect 6052 29668 6592 29696
rect 6052 29656 6058 29668
rect 5166 29588 5172 29640
rect 5224 29588 5230 29640
rect 5905 29631 5963 29637
rect 5905 29597 5917 29631
rect 5951 29628 5963 29631
rect 6012 29628 6040 29656
rect 5951 29600 6040 29628
rect 6089 29631 6147 29637
rect 5951 29597 5964 29600
rect 6089 29597 6101 29631
rect 6135 29597 6147 29631
rect 5905 29591 5963 29597
rect 6089 29591 6147 29597
rect 4062 29520 4068 29572
rect 4120 29520 4126 29572
rect 5718 29560 5724 29572
rect 5552 29532 5724 29560
rect 5552 29501 5580 29532
rect 5718 29520 5724 29532
rect 5776 29560 5782 29572
rect 6104 29560 6132 29591
rect 6564 29572 6592 29668
rect 7760 29668 7972 29696
rect 7374 29588 7380 29640
rect 7432 29588 7438 29640
rect 7561 29631 7619 29637
rect 7561 29597 7573 29631
rect 7607 29628 7619 29631
rect 7650 29628 7656 29640
rect 7607 29600 7656 29628
rect 7607 29597 7619 29600
rect 7561 29591 7619 29597
rect 7650 29588 7656 29600
rect 7708 29588 7714 29640
rect 7760 29637 7788 29668
rect 8938 29656 8944 29708
rect 8996 29656 9002 29708
rect 9600 29668 11652 29696
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 7837 29631 7895 29637
rect 7837 29597 7849 29631
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29628 7987 29631
rect 8202 29628 8208 29640
rect 7975 29600 8208 29628
rect 7975 29597 7987 29600
rect 7929 29591 7987 29597
rect 6365 29563 6423 29569
rect 6365 29560 6377 29563
rect 5776 29532 6377 29560
rect 5776 29520 5782 29532
rect 6365 29529 6377 29532
rect 6411 29529 6423 29563
rect 6365 29523 6423 29529
rect 5537 29495 5595 29501
rect 5537 29461 5549 29495
rect 5583 29461 5595 29495
rect 5537 29455 5595 29461
rect 6178 29452 6184 29504
rect 6236 29452 6242 29504
rect 6380 29492 6408 29523
rect 6546 29520 6552 29572
rect 6604 29520 6610 29572
rect 7392 29560 7420 29588
rect 7852 29560 7880 29591
rect 8202 29588 8208 29600
rect 8260 29628 8266 29640
rect 9600 29628 9628 29668
rect 11624 29640 11652 29668
rect 8260 29600 9628 29628
rect 8260 29588 8266 29600
rect 11054 29588 11060 29640
rect 11112 29628 11118 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 11112 29600 11437 29628
rect 11112 29588 11118 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 11514 29588 11520 29640
rect 11572 29588 11578 29640
rect 11606 29588 11612 29640
rect 11664 29588 11670 29640
rect 11790 29588 11796 29640
rect 11848 29588 11854 29640
rect 11882 29588 11888 29640
rect 11940 29588 11946 29640
rect 11992 29637 12020 29736
rect 12161 29733 12173 29767
rect 12207 29764 12219 29767
rect 12207 29736 12434 29764
rect 12207 29733 12219 29736
rect 12161 29727 12219 29733
rect 12406 29696 12434 29736
rect 12713 29699 12771 29705
rect 12713 29696 12725 29699
rect 12406 29668 12725 29696
rect 12713 29665 12725 29668
rect 12759 29665 12771 29699
rect 12713 29659 12771 29665
rect 11982 29631 12040 29637
rect 11982 29597 11994 29631
rect 12028 29597 12040 29631
rect 11982 29591 12040 29597
rect 12618 29588 12624 29640
rect 12676 29588 12682 29640
rect 12897 29631 12955 29637
rect 12897 29597 12909 29631
rect 12943 29628 12955 29631
rect 13372 29628 13400 29792
rect 17052 29764 17080 29804
rect 18598 29792 18604 29844
rect 18656 29832 18662 29844
rect 20806 29832 20812 29844
rect 18656 29804 20812 29832
rect 18656 29792 18662 29804
rect 20806 29792 20812 29804
rect 20864 29792 20870 29844
rect 21174 29792 21180 29844
rect 21232 29792 21238 29844
rect 24213 29835 24271 29841
rect 24213 29801 24225 29835
rect 24259 29832 24271 29835
rect 24394 29832 24400 29844
rect 24259 29804 24400 29832
rect 24259 29801 24271 29804
rect 24213 29795 24271 29801
rect 24394 29792 24400 29804
rect 24452 29792 24458 29844
rect 26234 29792 26240 29844
rect 26292 29832 26298 29844
rect 27249 29835 27307 29841
rect 27249 29832 27261 29835
rect 26292 29804 27261 29832
rect 26292 29792 26298 29804
rect 27249 29801 27261 29804
rect 27295 29801 27307 29835
rect 27249 29795 27307 29801
rect 27614 29792 27620 29844
rect 27672 29792 27678 29844
rect 33873 29835 33931 29841
rect 33873 29801 33885 29835
rect 33919 29832 33931 29835
rect 34054 29832 34060 29844
rect 33919 29804 34060 29832
rect 33919 29801 33931 29804
rect 33873 29795 33931 29801
rect 34054 29792 34060 29804
rect 34112 29792 34118 29844
rect 35434 29792 35440 29844
rect 35492 29832 35498 29844
rect 35529 29835 35587 29841
rect 35529 29832 35541 29835
rect 35492 29804 35541 29832
rect 35492 29792 35498 29804
rect 35529 29801 35541 29804
rect 35575 29832 35587 29835
rect 35894 29832 35900 29844
rect 35575 29804 35900 29832
rect 35575 29801 35587 29804
rect 35529 29795 35587 29801
rect 35894 29792 35900 29804
rect 35952 29792 35958 29844
rect 38562 29792 38568 29844
rect 38620 29792 38626 29844
rect 38933 29835 38991 29841
rect 38933 29801 38945 29835
rect 38979 29832 38991 29835
rect 41138 29832 41144 29844
rect 38979 29804 41144 29832
rect 38979 29801 38991 29804
rect 38933 29795 38991 29801
rect 41138 29792 41144 29804
rect 41196 29792 41202 29844
rect 42518 29792 42524 29844
rect 42576 29832 42582 29844
rect 42613 29835 42671 29841
rect 42613 29832 42625 29835
rect 42576 29804 42625 29832
rect 42576 29792 42582 29804
rect 42613 29801 42625 29804
rect 42659 29801 42671 29835
rect 42613 29795 42671 29801
rect 21192 29764 21220 29792
rect 17052 29736 21220 29764
rect 15378 29696 15384 29708
rect 12943 29600 13400 29628
rect 14384 29668 15384 29696
rect 12943 29597 12955 29600
rect 12897 29591 12955 29597
rect 14384 29560 14412 29668
rect 15378 29656 15384 29668
rect 15436 29656 15442 29708
rect 15749 29699 15807 29705
rect 15749 29665 15761 29699
rect 15795 29696 15807 29699
rect 16574 29696 16580 29708
rect 15795 29668 16580 29696
rect 15795 29665 15807 29668
rect 15749 29659 15807 29665
rect 16574 29656 16580 29668
rect 16632 29656 16638 29708
rect 17218 29696 17224 29708
rect 17144 29668 17224 29696
rect 17144 29614 17172 29668
rect 17218 29656 17224 29668
rect 17276 29656 17282 29708
rect 17773 29699 17831 29705
rect 17773 29665 17785 29699
rect 17819 29696 17831 29699
rect 18230 29696 18236 29708
rect 17819 29668 18236 29696
rect 17819 29665 17831 29668
rect 17773 29659 17831 29665
rect 18230 29656 18236 29668
rect 18288 29696 18294 29708
rect 19058 29696 19064 29708
rect 18288 29668 19064 29696
rect 18288 29656 18294 29668
rect 19058 29656 19064 29668
rect 19116 29656 19122 29708
rect 20254 29656 20260 29708
rect 20312 29696 20318 29708
rect 20990 29696 20996 29708
rect 20312 29668 20996 29696
rect 20312 29656 20318 29668
rect 20990 29656 20996 29668
rect 21048 29656 21054 29708
rect 24118 29656 24124 29708
rect 24176 29696 24182 29708
rect 24949 29699 25007 29705
rect 24949 29696 24961 29699
rect 24176 29668 24961 29696
rect 24176 29656 24182 29668
rect 24949 29665 24961 29668
rect 24995 29665 25007 29699
rect 24949 29659 25007 29665
rect 17954 29588 17960 29640
rect 18012 29588 18018 29640
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29628 24087 29631
rect 24075 29600 24440 29628
rect 24075 29597 24087 29600
rect 24029 29591 24087 29597
rect 7392 29532 7880 29560
rect 7944 29532 14412 29560
rect 7944 29492 7972 29532
rect 16022 29520 16028 29572
rect 16080 29520 16086 29572
rect 17310 29520 17316 29572
rect 17368 29560 17374 29572
rect 17368 29532 20392 29560
rect 17368 29520 17374 29532
rect 20364 29504 20392 29532
rect 6380 29464 7972 29492
rect 8846 29452 8852 29504
rect 8904 29492 8910 29504
rect 9585 29495 9643 29501
rect 9585 29492 9597 29495
rect 8904 29464 9597 29492
rect 8904 29452 8910 29464
rect 9585 29461 9597 29464
rect 9631 29461 9643 29495
rect 9585 29455 9643 29461
rect 11238 29452 11244 29504
rect 11296 29492 11302 29504
rect 12986 29492 12992 29504
rect 11296 29464 12992 29492
rect 11296 29452 11302 29464
rect 12986 29452 12992 29464
rect 13044 29452 13050 29504
rect 13081 29495 13139 29501
rect 13081 29461 13093 29495
rect 13127 29492 13139 29495
rect 14274 29492 14280 29504
rect 13127 29464 14280 29492
rect 13127 29461 13139 29464
rect 13081 29455 13139 29461
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 17494 29452 17500 29504
rect 17552 29452 17558 29504
rect 17862 29452 17868 29504
rect 17920 29452 17926 29504
rect 18322 29452 18328 29504
rect 18380 29452 18386 29504
rect 20346 29452 20352 29504
rect 20404 29452 20410 29504
rect 24412 29501 24440 29600
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24544 29600 24777 29628
rect 24544 29588 24550 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 27249 29631 27307 29637
rect 27249 29597 27261 29631
rect 27295 29597 27307 29631
rect 27249 29591 27307 29597
rect 27264 29560 27292 29591
rect 27430 29588 27436 29640
rect 27488 29588 27494 29640
rect 33962 29588 33968 29640
rect 34020 29588 34026 29640
rect 34072 29628 34100 29792
rect 38580 29764 38608 29792
rect 39025 29767 39083 29773
rect 39025 29764 39037 29767
rect 38580 29736 39037 29764
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 34072 29600 34161 29628
rect 34149 29597 34161 29600
rect 34195 29597 34207 29631
rect 34149 29591 34207 29597
rect 34698 29588 34704 29640
rect 34756 29628 34762 29640
rect 35253 29631 35311 29637
rect 35253 29628 35265 29631
rect 34756 29600 35265 29628
rect 34756 29588 34762 29600
rect 35253 29597 35265 29600
rect 35299 29597 35311 29631
rect 35253 29591 35311 29597
rect 38381 29631 38439 29637
rect 38381 29597 38393 29631
rect 38427 29628 38439 29631
rect 38580 29628 38608 29736
rect 39025 29733 39037 29736
rect 39071 29733 39083 29767
rect 39025 29727 39083 29733
rect 41141 29699 41199 29705
rect 41141 29665 41153 29699
rect 41187 29696 41199 29699
rect 41230 29696 41236 29708
rect 41187 29668 41236 29696
rect 41187 29665 41199 29668
rect 41141 29659 41199 29665
rect 41230 29656 41236 29668
rect 41288 29656 41294 29708
rect 43070 29656 43076 29708
rect 43128 29696 43134 29708
rect 43165 29699 43223 29705
rect 43165 29696 43177 29699
rect 43128 29668 43177 29696
rect 43128 29656 43134 29668
rect 43165 29665 43177 29668
rect 43211 29665 43223 29699
rect 43165 29659 43223 29665
rect 43257 29699 43315 29705
rect 43257 29665 43269 29699
rect 43303 29665 43315 29699
rect 43257 29659 43315 29665
rect 38427 29600 38608 29628
rect 38427 29597 38439 29600
rect 38381 29591 38439 29597
rect 38746 29588 38752 29640
rect 38804 29628 38810 29640
rect 39114 29628 39120 29640
rect 38804 29600 39120 29628
rect 38804 29588 38810 29600
rect 39114 29588 39120 29600
rect 39172 29588 39178 29640
rect 39669 29631 39727 29637
rect 39669 29597 39681 29631
rect 39715 29597 39727 29631
rect 39669 29591 39727 29597
rect 33505 29563 33563 29569
rect 33505 29560 33517 29563
rect 27264 29532 27660 29560
rect 27632 29504 27660 29532
rect 33428 29532 33517 29560
rect 33428 29504 33456 29532
rect 33505 29529 33517 29532
rect 33551 29529 33563 29563
rect 33505 29523 33563 29529
rect 33686 29520 33692 29572
rect 33744 29520 33750 29572
rect 38010 29520 38016 29572
rect 38068 29560 38074 29572
rect 38470 29560 38476 29572
rect 38068 29532 38476 29560
rect 38068 29520 38074 29532
rect 38470 29520 38476 29532
rect 38528 29560 38534 29572
rect 38565 29563 38623 29569
rect 38565 29560 38577 29563
rect 38528 29532 38577 29560
rect 38528 29520 38534 29532
rect 38565 29529 38577 29532
rect 38611 29529 38623 29563
rect 38565 29523 38623 29529
rect 38657 29563 38715 29569
rect 38657 29529 38669 29563
rect 38703 29529 38715 29563
rect 38657 29523 38715 29529
rect 24397 29495 24455 29501
rect 24397 29461 24409 29495
rect 24443 29461 24455 29495
rect 24397 29455 24455 29461
rect 24857 29495 24915 29501
rect 24857 29461 24869 29495
rect 24903 29492 24915 29495
rect 26326 29492 26332 29504
rect 24903 29464 26332 29492
rect 24903 29461 24915 29464
rect 24857 29455 24915 29461
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 27614 29452 27620 29504
rect 27672 29452 27678 29504
rect 33410 29452 33416 29504
rect 33468 29452 33474 29504
rect 34149 29495 34207 29501
rect 34149 29461 34161 29495
rect 34195 29492 34207 29495
rect 34422 29492 34428 29504
rect 34195 29464 34428 29492
rect 34195 29461 34207 29464
rect 34149 29455 34207 29461
rect 34422 29452 34428 29464
rect 34480 29452 34486 29504
rect 38672 29492 38700 29523
rect 38838 29520 38844 29572
rect 38896 29560 38902 29572
rect 39684 29560 39712 29591
rect 39850 29588 39856 29640
rect 39908 29588 39914 29640
rect 40770 29588 40776 29640
rect 40828 29628 40834 29640
rect 40865 29631 40923 29637
rect 40865 29628 40877 29631
rect 40828 29600 40877 29628
rect 40828 29588 40834 29600
rect 40865 29597 40877 29600
rect 40911 29597 40923 29631
rect 43272 29628 43300 29659
rect 40865 29591 40923 29597
rect 43180 29600 43300 29628
rect 41046 29560 41052 29572
rect 38896 29532 41052 29560
rect 38896 29520 38902 29532
rect 41046 29520 41052 29532
rect 41104 29520 41110 29572
rect 42978 29560 42984 29572
rect 41248 29532 41630 29560
rect 42628 29532 42984 29560
rect 38930 29492 38936 29504
rect 38672 29464 38936 29492
rect 38930 29452 38936 29464
rect 38988 29452 38994 29504
rect 40494 29452 40500 29504
rect 40552 29452 40558 29504
rect 40678 29452 40684 29504
rect 40736 29492 40742 29504
rect 41248 29492 41276 29532
rect 40736 29464 41276 29492
rect 41524 29492 41552 29532
rect 42628 29492 42656 29532
rect 42978 29520 42984 29532
rect 43036 29520 43042 29572
rect 43180 29504 43208 29600
rect 41524 29464 42656 29492
rect 40736 29452 40742 29464
rect 42702 29452 42708 29504
rect 42760 29452 42766 29504
rect 43070 29452 43076 29504
rect 43128 29452 43134 29504
rect 43162 29452 43168 29504
rect 43220 29452 43226 29504
rect 1104 29402 44620 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 44620 29402
rect 1104 29328 44620 29350
rect 4062 29248 4068 29300
rect 4120 29288 4126 29300
rect 4157 29291 4215 29297
rect 4157 29288 4169 29291
rect 4120 29260 4169 29288
rect 4120 29248 4126 29260
rect 4157 29257 4169 29260
rect 4203 29257 4215 29291
rect 4157 29251 4215 29257
rect 5337 29291 5395 29297
rect 5337 29257 5349 29291
rect 5383 29288 5395 29291
rect 5721 29291 5779 29297
rect 5721 29288 5733 29291
rect 5383 29260 5733 29288
rect 5383 29257 5395 29260
rect 5337 29251 5395 29257
rect 5721 29257 5733 29260
rect 5767 29257 5779 29291
rect 5721 29251 5779 29257
rect 7742 29248 7748 29300
rect 7800 29288 7806 29300
rect 8662 29288 8668 29300
rect 7800 29260 8668 29288
rect 7800 29248 7806 29260
rect 8662 29248 8668 29260
rect 8720 29248 8726 29300
rect 9217 29291 9275 29297
rect 9217 29257 9229 29291
rect 9263 29257 9275 29291
rect 9217 29251 9275 29257
rect 5442 29180 5448 29232
rect 5500 29180 5506 29232
rect 5534 29180 5540 29232
rect 5592 29220 5598 29232
rect 7190 29220 7196 29232
rect 5592 29192 7196 29220
rect 5592 29180 5598 29192
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 9232 29220 9260 29251
rect 9490 29248 9496 29300
rect 9548 29288 9554 29300
rect 9548 29260 9720 29288
rect 9548 29248 9554 29260
rect 9585 29223 9643 29229
rect 9585 29220 9597 29223
rect 9232 29192 9597 29220
rect 9585 29189 9597 29192
rect 9631 29189 9643 29223
rect 9692 29220 9720 29260
rect 11054 29248 11060 29300
rect 11112 29288 11118 29300
rect 15102 29288 15108 29300
rect 11112 29260 15108 29288
rect 11112 29248 11118 29260
rect 15102 29248 15108 29260
rect 15160 29248 15166 29300
rect 16022 29248 16028 29300
rect 16080 29288 16086 29300
rect 16669 29291 16727 29297
rect 16669 29288 16681 29291
rect 16080 29260 16681 29288
rect 16080 29248 16086 29260
rect 16669 29257 16681 29260
rect 16715 29257 16727 29291
rect 16669 29251 16727 29257
rect 16942 29248 16948 29300
rect 17000 29248 17006 29300
rect 17494 29248 17500 29300
rect 17552 29248 17558 29300
rect 17862 29248 17868 29300
rect 17920 29288 17926 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17920 29260 17969 29288
rect 17920 29248 17926 29260
rect 17957 29257 17969 29260
rect 18003 29257 18015 29291
rect 17957 29251 18015 29257
rect 18046 29248 18052 29300
rect 18104 29248 18110 29300
rect 18322 29248 18328 29300
rect 18380 29248 18386 29300
rect 20349 29291 20407 29297
rect 20349 29288 20361 29291
rect 20088 29260 20361 29288
rect 9692 29192 10074 29220
rect 9585 29183 9643 29189
rect 13078 29180 13084 29232
rect 13136 29220 13142 29232
rect 13446 29220 13452 29232
rect 13136 29192 13452 29220
rect 13136 29180 13142 29192
rect 13446 29180 13452 29192
rect 13504 29220 13510 29232
rect 13722 29220 13728 29232
rect 13504 29192 13728 29220
rect 13504 29180 13510 29192
rect 13722 29180 13728 29192
rect 13780 29180 13786 29232
rect 16960 29220 16988 29248
rect 16960 29192 17172 29220
rect 4341 29155 4399 29161
rect 4341 29121 4353 29155
rect 4387 29152 4399 29155
rect 5460 29152 5488 29180
rect 17144 29164 17172 29192
rect 5813 29155 5871 29161
rect 5813 29152 5825 29155
rect 4387 29124 5212 29152
rect 5460 29124 5825 29152
rect 4387 29121 4399 29124
rect 4341 29115 4399 29121
rect 5184 29025 5212 29124
rect 5813 29121 5825 29124
rect 5859 29121 5871 29155
rect 5813 29115 5871 29121
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29152 9091 29155
rect 9214 29152 9220 29164
rect 9079 29124 9220 29152
rect 9079 29121 9091 29124
rect 9033 29115 9091 29121
rect 9214 29112 9220 29124
rect 9272 29112 9278 29164
rect 16853 29155 16911 29161
rect 16853 29121 16865 29155
rect 16899 29152 16911 29155
rect 17037 29155 17095 29161
rect 16899 29124 16988 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 9306 29044 9312 29096
rect 9364 29044 9370 29096
rect 16960 29028 16988 29124
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17052 29084 17080 29115
rect 17126 29112 17132 29164
rect 17184 29112 17190 29164
rect 17405 29155 17463 29161
rect 17405 29121 17417 29155
rect 17451 29152 17463 29155
rect 17512 29152 17540 29248
rect 17451 29124 17540 29152
rect 17451 29121 17463 29124
rect 17405 29115 17463 29121
rect 17880 29084 17908 29248
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29152 18291 29155
rect 18340 29152 18368 29248
rect 20088 29229 20116 29260
rect 20349 29257 20361 29260
rect 20395 29288 20407 29291
rect 20530 29288 20536 29300
rect 20395 29260 20536 29288
rect 20395 29257 20407 29260
rect 20349 29251 20407 29257
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 20993 29291 21051 29297
rect 20993 29288 21005 29291
rect 20956 29260 21005 29288
rect 20956 29248 20962 29260
rect 20993 29257 21005 29260
rect 21039 29257 21051 29291
rect 20993 29251 21051 29257
rect 27525 29291 27583 29297
rect 27525 29257 27537 29291
rect 27571 29257 27583 29291
rect 27525 29251 27583 29257
rect 20073 29223 20131 29229
rect 20073 29189 20085 29223
rect 20119 29189 20131 29223
rect 20073 29183 20131 29189
rect 20254 29180 20260 29232
rect 20312 29180 20318 29232
rect 20438 29220 20444 29232
rect 20364 29192 20444 29220
rect 18279 29124 18368 29152
rect 18279 29121 18291 29124
rect 18233 29115 18291 29121
rect 18690 29112 18696 29164
rect 18748 29112 18754 29164
rect 19334 29112 19340 29164
rect 19392 29112 19398 29164
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 19978 29152 19984 29164
rect 19935 29124 19984 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20364 29152 20392 29192
rect 20438 29180 20444 29192
rect 20496 29220 20502 29232
rect 20625 29223 20683 29229
rect 20625 29220 20637 29223
rect 20496 29192 20637 29220
rect 20496 29180 20502 29192
rect 20625 29189 20637 29192
rect 20671 29220 20683 29223
rect 21177 29223 21235 29229
rect 21177 29220 21189 29223
rect 20671 29192 21189 29220
rect 20671 29189 20683 29192
rect 20625 29183 20683 29189
rect 21177 29189 21189 29192
rect 21223 29189 21235 29223
rect 21177 29183 21235 29189
rect 21361 29223 21419 29229
rect 21361 29189 21373 29223
rect 21407 29220 21419 29223
rect 22186 29220 22192 29232
rect 21407 29192 22192 29220
rect 21407 29189 21419 29192
rect 21361 29183 21419 29189
rect 20806 29161 20812 29164
rect 20088 29124 20392 29152
rect 20533 29155 20591 29161
rect 17052 29056 17908 29084
rect 5169 29019 5227 29025
rect 5169 28985 5181 29019
rect 5215 28985 5227 29019
rect 5169 28979 5227 28985
rect 16942 28976 16948 29028
rect 17000 29016 17006 29028
rect 18708 29016 18736 29112
rect 19352 29084 19380 29112
rect 20088 29084 20116 29124
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20763 29155 20812 29161
rect 20763 29121 20775 29155
rect 20809 29121 20812 29155
rect 20763 29115 20812 29121
rect 19352 29056 20116 29084
rect 20548 29084 20576 29115
rect 20806 29112 20812 29115
rect 20864 29112 20870 29164
rect 20901 29155 20959 29161
rect 20901 29121 20913 29155
rect 20947 29152 20959 29155
rect 20990 29152 20996 29164
rect 20947 29124 20996 29152
rect 20947 29121 20959 29124
rect 20901 29115 20959 29121
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 21376 29084 21404 29183
rect 22186 29180 22192 29192
rect 22244 29180 22250 29232
rect 23014 29180 23020 29232
rect 23072 29180 23078 29232
rect 27540 29220 27568 29251
rect 28994 29248 29000 29300
rect 29052 29288 29058 29300
rect 32125 29291 32183 29297
rect 32125 29288 32137 29291
rect 29052 29260 32137 29288
rect 29052 29248 29058 29260
rect 32125 29257 32137 29260
rect 32171 29257 32183 29291
rect 32125 29251 32183 29257
rect 33597 29291 33655 29297
rect 33597 29257 33609 29291
rect 33643 29288 33655 29291
rect 33962 29288 33968 29300
rect 33643 29260 33968 29288
rect 33643 29257 33655 29260
rect 33597 29251 33655 29257
rect 33962 29248 33968 29260
rect 34020 29248 34026 29300
rect 37461 29291 37519 29297
rect 37461 29257 37473 29291
rect 37507 29288 37519 29291
rect 37826 29288 37832 29300
rect 37507 29260 37832 29288
rect 37507 29257 37519 29260
rect 37461 29251 37519 29257
rect 37826 29248 37832 29260
rect 37884 29248 37890 29300
rect 40586 29288 40592 29300
rect 40420 29260 40592 29288
rect 34606 29220 34612 29232
rect 27540 29192 31754 29220
rect 26326 29112 26332 29164
rect 26384 29152 26390 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 26384 29124 27169 29152
rect 26384 29112 26390 29124
rect 27157 29121 27169 29124
rect 27203 29152 27215 29155
rect 27430 29152 27436 29164
rect 27203 29124 27436 29152
rect 27203 29121 27215 29124
rect 27157 29115 27215 29121
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 27890 29112 27896 29164
rect 27948 29112 27954 29164
rect 29086 29112 29092 29164
rect 29144 29152 29150 29164
rect 30285 29155 30343 29161
rect 30285 29152 30297 29155
rect 29144 29124 30297 29152
rect 29144 29112 29150 29124
rect 30285 29121 30297 29124
rect 30331 29121 30343 29155
rect 30285 29115 30343 29121
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29121 30527 29155
rect 30469 29115 30527 29121
rect 30653 29155 30711 29161
rect 30653 29121 30665 29155
rect 30699 29152 30711 29155
rect 31202 29152 31208 29164
rect 30699 29124 31208 29152
rect 30699 29121 30711 29124
rect 30653 29115 30711 29121
rect 20548 29056 21404 29084
rect 27249 29087 27307 29093
rect 27249 29053 27261 29087
rect 27295 29053 27307 29087
rect 27249 29047 27307 29053
rect 27264 29016 27292 29047
rect 27522 29044 27528 29096
rect 27580 29084 27586 29096
rect 27617 29087 27675 29093
rect 27617 29084 27629 29087
rect 27580 29056 27629 29084
rect 27580 29044 27586 29056
rect 27617 29053 27629 29056
rect 27663 29053 27675 29087
rect 27617 29047 27675 29053
rect 28077 29019 28135 29025
rect 28077 29016 28089 29019
rect 17000 28988 18736 29016
rect 24412 28988 24808 29016
rect 27264 28988 28089 29016
rect 17000 28976 17006 28988
rect 5353 28951 5411 28957
rect 5353 28917 5365 28951
rect 5399 28948 5411 28951
rect 6178 28948 6184 28960
rect 5399 28920 6184 28948
rect 5399 28917 5411 28920
rect 5353 28911 5411 28917
rect 6178 28908 6184 28920
rect 6236 28908 6242 28960
rect 17494 28908 17500 28960
rect 17552 28948 17558 28960
rect 24412 28948 24440 28988
rect 17552 28920 24440 28948
rect 24489 28951 24547 28957
rect 17552 28908 17558 28920
rect 24489 28917 24501 28951
rect 24535 28948 24547 28951
rect 24670 28948 24676 28960
rect 24535 28920 24676 28948
rect 24535 28917 24547 28920
rect 24489 28911 24547 28917
rect 24670 28908 24676 28920
rect 24728 28908 24734 28960
rect 24780 28948 24808 28988
rect 28077 28985 28089 28988
rect 28123 28985 28135 29019
rect 28077 28979 28135 28985
rect 26786 28948 26792 28960
rect 24780 28920 26792 28948
rect 26786 28908 26792 28920
rect 26844 28908 26850 28960
rect 27614 28908 27620 28960
rect 27672 28948 27678 28960
rect 27709 28951 27767 28957
rect 27709 28948 27721 28951
rect 27672 28920 27721 28948
rect 27672 28908 27678 28920
rect 27709 28917 27721 28920
rect 27755 28917 27767 28951
rect 30300 28948 30328 29115
rect 30484 29084 30512 29115
rect 31202 29112 31208 29124
rect 31260 29152 31266 29164
rect 31297 29155 31355 29161
rect 31297 29152 31309 29155
rect 31260 29124 31309 29152
rect 31260 29112 31266 29124
rect 31297 29121 31309 29124
rect 31343 29121 31355 29155
rect 31297 29115 31355 29121
rect 31481 29155 31539 29161
rect 31481 29121 31493 29155
rect 31527 29152 31539 29155
rect 31570 29152 31576 29164
rect 31527 29124 31576 29152
rect 31527 29121 31539 29124
rect 31481 29115 31539 29121
rect 31570 29112 31576 29124
rect 31628 29112 31634 29164
rect 31726 29084 31754 29192
rect 33520 29192 34612 29220
rect 33410 29152 33416 29164
rect 32692 29124 33416 29152
rect 32692 29084 32720 29124
rect 33410 29112 33416 29124
rect 33468 29112 33474 29164
rect 30484 29056 31064 29084
rect 31726 29056 32720 29084
rect 32769 29087 32827 29093
rect 31036 29028 31064 29056
rect 32769 29053 32781 29087
rect 32815 29084 32827 29087
rect 33520 29084 33548 29192
rect 34606 29180 34612 29192
rect 34664 29180 34670 29232
rect 34698 29180 34704 29232
rect 34756 29220 34762 29232
rect 34885 29223 34943 29229
rect 34885 29220 34897 29223
rect 34756 29192 34897 29220
rect 34756 29180 34762 29192
rect 34885 29189 34897 29192
rect 34931 29189 34943 29223
rect 38930 29220 38936 29232
rect 34885 29183 34943 29189
rect 37660 29192 38936 29220
rect 33597 29155 33655 29161
rect 33597 29121 33609 29155
rect 33643 29152 33655 29155
rect 33686 29152 33692 29164
rect 33643 29124 33692 29152
rect 33643 29121 33655 29124
rect 33597 29115 33655 29121
rect 33686 29112 33692 29124
rect 33744 29152 33750 29164
rect 37660 29161 37688 29192
rect 38930 29180 38936 29192
rect 38988 29180 38994 29232
rect 40420 29229 40448 29260
rect 40586 29248 40592 29260
rect 40644 29248 40650 29300
rect 42702 29248 42708 29300
rect 42760 29248 42766 29300
rect 40405 29223 40463 29229
rect 40405 29189 40417 29223
rect 40451 29189 40463 29223
rect 40405 29183 40463 29189
rect 37645 29155 37703 29161
rect 33744 29124 34008 29152
rect 33744 29112 33750 29124
rect 32815 29056 33548 29084
rect 32815 29053 32827 29056
rect 32769 29047 32827 29053
rect 33980 29028 34008 29124
rect 37645 29121 37657 29155
rect 37691 29121 37703 29155
rect 37645 29115 37703 29121
rect 37921 29155 37979 29161
rect 37921 29121 37933 29155
rect 37967 29152 37979 29155
rect 37967 29124 38516 29152
rect 37967 29121 37979 29124
rect 37921 29115 37979 29121
rect 36538 29044 36544 29096
rect 36596 29044 36602 29096
rect 37826 29044 37832 29096
rect 37884 29044 37890 29096
rect 31018 28976 31024 29028
rect 31076 28976 31082 29028
rect 31389 29019 31447 29025
rect 31389 28985 31401 29019
rect 31435 29016 31447 29019
rect 32122 29016 32128 29028
rect 31435 28988 32128 29016
rect 31435 28985 31447 28988
rect 31389 28979 31447 28985
rect 32122 28976 32128 28988
rect 32180 28976 32186 29028
rect 33962 28976 33968 29028
rect 34020 28976 34026 29028
rect 34514 28976 34520 29028
rect 34572 29016 34578 29028
rect 34609 29019 34667 29025
rect 34609 29016 34621 29019
rect 34572 28988 34621 29016
rect 34572 28976 34578 28988
rect 34609 28985 34621 28988
rect 34655 28985 34667 29019
rect 34609 28979 34667 28985
rect 38013 29019 38071 29025
rect 38013 28985 38025 29019
rect 38059 29016 38071 29019
rect 38194 29016 38200 29028
rect 38059 28988 38200 29016
rect 38059 28985 38071 28988
rect 38013 28979 38071 28985
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 38488 29016 38516 29124
rect 38654 29112 38660 29164
rect 38712 29112 38718 29164
rect 39298 29112 39304 29164
rect 39356 29112 39362 29164
rect 42061 29155 42119 29161
rect 42061 29121 42073 29155
rect 42107 29152 42119 29155
rect 42720 29152 42748 29248
rect 42794 29180 42800 29232
rect 42852 29220 42858 29232
rect 42889 29223 42947 29229
rect 42889 29220 42901 29223
rect 42852 29192 42901 29220
rect 42852 29180 42858 29192
rect 42889 29189 42901 29192
rect 42935 29189 42947 29223
rect 42889 29183 42947 29189
rect 42107 29124 42748 29152
rect 42107 29121 42119 29124
rect 42061 29115 42119 29121
rect 40681 29087 40739 29093
rect 40681 29053 40693 29087
rect 40727 29084 40739 29087
rect 40862 29084 40868 29096
rect 40727 29056 40868 29084
rect 40727 29053 40739 29056
rect 40681 29047 40739 29053
rect 40862 29044 40868 29056
rect 40920 29044 40926 29096
rect 42886 29044 42892 29096
rect 42944 29084 42950 29096
rect 43441 29087 43499 29093
rect 43441 29084 43453 29087
rect 42944 29056 43453 29084
rect 42944 29044 42950 29056
rect 43441 29053 43453 29056
rect 43487 29053 43499 29087
rect 43441 29047 43499 29053
rect 39206 29016 39212 29028
rect 38488 28988 39212 29016
rect 39206 28976 39212 28988
rect 39264 28976 39270 29028
rect 31938 28948 31944 28960
rect 30300 28920 31944 28948
rect 27709 28911 27767 28917
rect 31938 28908 31944 28920
rect 31996 28908 32002 28960
rect 35986 28908 35992 28960
rect 36044 28908 36050 28960
rect 37921 28951 37979 28957
rect 37921 28917 37933 28951
rect 37967 28948 37979 28951
rect 38838 28948 38844 28960
rect 37967 28920 38844 28948
rect 37967 28917 37979 28920
rect 37921 28911 37979 28917
rect 38838 28908 38844 28920
rect 38896 28908 38902 28960
rect 38930 28908 38936 28960
rect 38988 28948 38994 28960
rect 39942 28948 39948 28960
rect 38988 28920 39948 28948
rect 38988 28908 38994 28920
rect 39942 28908 39948 28920
rect 40000 28908 40006 28960
rect 42245 28951 42303 28957
rect 42245 28917 42257 28951
rect 42291 28948 42303 28951
rect 42426 28948 42432 28960
rect 42291 28920 42432 28948
rect 42291 28917 42303 28920
rect 42245 28911 42303 28917
rect 42426 28908 42432 28920
rect 42484 28908 42490 28960
rect 1104 28858 44620 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 44620 28858
rect 1104 28784 44620 28806
rect 7098 28704 7104 28756
rect 7156 28704 7162 28756
rect 8389 28747 8447 28753
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 9125 28747 9183 28753
rect 9125 28744 9137 28747
rect 8435 28716 9137 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 9125 28713 9137 28716
rect 9171 28713 9183 28747
rect 9125 28707 9183 28713
rect 9214 28704 9220 28756
rect 9272 28744 9278 28756
rect 9309 28747 9367 28753
rect 9309 28744 9321 28747
rect 9272 28716 9321 28744
rect 9272 28704 9278 28716
rect 9309 28713 9321 28716
rect 9355 28713 9367 28747
rect 9309 28707 9367 28713
rect 10410 28704 10416 28756
rect 10468 28704 10474 28756
rect 11514 28704 11520 28756
rect 11572 28704 11578 28756
rect 14737 28747 14795 28753
rect 14737 28713 14749 28747
rect 14783 28744 14795 28747
rect 14918 28744 14924 28756
rect 14783 28716 14924 28744
rect 14783 28713 14795 28716
rect 14737 28707 14795 28713
rect 14918 28704 14924 28716
rect 14976 28704 14982 28756
rect 16942 28704 16948 28756
rect 17000 28704 17006 28756
rect 19978 28704 19984 28756
rect 20036 28744 20042 28756
rect 20073 28747 20131 28753
rect 20073 28744 20085 28747
rect 20036 28716 20085 28744
rect 20036 28704 20042 28716
rect 20073 28713 20085 28716
rect 20119 28713 20131 28747
rect 20073 28707 20131 28713
rect 20809 28747 20867 28753
rect 20809 28713 20821 28747
rect 20855 28744 20867 28747
rect 21174 28744 21180 28756
rect 20855 28716 21180 28744
rect 20855 28713 20867 28716
rect 20809 28707 20867 28713
rect 21174 28704 21180 28716
rect 21232 28704 21238 28756
rect 29086 28704 29092 28756
rect 29144 28704 29150 28756
rect 32582 28744 32588 28756
rect 30116 28716 32588 28744
rect 6917 28679 6975 28685
rect 6917 28645 6929 28679
rect 6963 28645 6975 28679
rect 8573 28679 8631 28685
rect 8573 28676 8585 28679
rect 6917 28639 6975 28645
rect 8312 28648 8585 28676
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 6546 28608 6552 28620
rect 5592 28580 6552 28608
rect 5592 28568 5598 28580
rect 6546 28568 6552 28580
rect 6604 28608 6610 28620
rect 6932 28608 6960 28639
rect 6604 28580 6960 28608
rect 6604 28568 6610 28580
rect 7190 28568 7196 28620
rect 7248 28608 7254 28620
rect 7248 28580 7420 28608
rect 7248 28568 7254 28580
rect 7392 28549 7420 28580
rect 7466 28568 7472 28620
rect 7524 28608 7530 28620
rect 8312 28608 8340 28648
rect 8573 28645 8585 28648
rect 8619 28645 8631 28679
rect 8573 28639 8631 28645
rect 9030 28608 9036 28620
rect 7524 28580 8340 28608
rect 7524 28568 7530 28580
rect 8312 28549 8340 28580
rect 8588 28580 9036 28608
rect 8588 28549 8616 28580
rect 9030 28568 9036 28580
rect 9088 28568 9094 28620
rect 10428 28608 10456 28704
rect 13541 28679 13599 28685
rect 13541 28645 13553 28679
rect 13587 28676 13599 28679
rect 16960 28676 16988 28704
rect 13587 28648 16988 28676
rect 13587 28645 13599 28648
rect 13541 28639 13599 28645
rect 20346 28636 20352 28688
rect 20404 28676 20410 28688
rect 27985 28679 28043 28685
rect 27985 28676 27997 28679
rect 20404 28648 20484 28676
rect 20404 28636 20410 28648
rect 9416 28580 10456 28608
rect 11241 28611 11299 28617
rect 9416 28549 9444 28580
rect 11241 28577 11253 28611
rect 11287 28577 11299 28611
rect 11241 28571 11299 28577
rect 14461 28611 14519 28617
rect 14461 28577 14473 28611
rect 14507 28608 14519 28611
rect 14918 28608 14924 28620
rect 14507 28580 14924 28608
rect 14507 28577 14519 28580
rect 14461 28571 14519 28577
rect 6641 28543 6699 28549
rect 6641 28509 6653 28543
rect 6687 28509 6699 28543
rect 6641 28503 6699 28509
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28540 6883 28543
rect 7377 28543 7435 28549
rect 6871 28512 7236 28540
rect 6871 28509 6883 28512
rect 6825 28503 6883 28509
rect 6656 28472 6684 28503
rect 7208 28484 7236 28512
rect 7377 28509 7389 28543
rect 7423 28509 7435 28543
rect 7377 28503 7435 28509
rect 8297 28543 8355 28549
rect 8297 28509 8309 28543
rect 8343 28509 8355 28543
rect 8297 28503 8355 28509
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28509 8631 28543
rect 8573 28503 8631 28509
rect 8757 28543 8815 28549
rect 8757 28509 8769 28543
rect 8803 28540 8815 28543
rect 9401 28543 9459 28549
rect 9401 28540 9413 28543
rect 8803 28512 9413 28540
rect 8803 28509 8815 28512
rect 8757 28503 8815 28509
rect 9401 28509 9413 28512
rect 9447 28509 9459 28543
rect 9401 28503 9459 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28509 11207 28543
rect 11256 28540 11284 28571
rect 14918 28568 14924 28580
rect 14976 28568 14982 28620
rect 18046 28608 18052 28620
rect 16316 28580 18052 28608
rect 11606 28540 11612 28552
rect 11256 28512 11612 28540
rect 11149 28503 11207 28509
rect 6656 28444 7128 28472
rect 6086 28364 6092 28416
rect 6144 28404 6150 28416
rect 7100 28413 7128 28444
rect 7190 28432 7196 28484
rect 7248 28472 7254 28484
rect 7285 28475 7343 28481
rect 7285 28472 7297 28475
rect 7248 28444 7297 28472
rect 7248 28432 7254 28444
rect 7285 28441 7297 28444
rect 7331 28441 7343 28475
rect 7392 28472 7420 28503
rect 8967 28475 9025 28481
rect 8967 28472 8979 28475
rect 7392 28444 8156 28472
rect 7285 28435 7343 28441
rect 6457 28407 6515 28413
rect 6457 28404 6469 28407
rect 6144 28376 6469 28404
rect 6144 28364 6150 28376
rect 6457 28373 6469 28376
rect 6503 28373 6515 28407
rect 6457 28367 6515 28373
rect 7085 28407 7143 28413
rect 7085 28373 7097 28407
rect 7131 28404 7143 28407
rect 7466 28404 7472 28416
rect 7131 28376 7472 28404
rect 7131 28373 7143 28376
rect 7085 28367 7143 28373
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 7561 28407 7619 28413
rect 7561 28373 7573 28407
rect 7607 28404 7619 28407
rect 7742 28404 7748 28416
rect 7607 28376 7748 28404
rect 7607 28373 7619 28376
rect 7561 28367 7619 28373
rect 7742 28364 7748 28376
rect 7800 28364 7806 28416
rect 8128 28404 8156 28444
rect 8772 28444 8979 28472
rect 8772 28416 8800 28444
rect 8967 28441 8979 28444
rect 9013 28441 9025 28475
rect 8967 28435 9025 28441
rect 9157 28475 9215 28481
rect 9157 28441 9169 28475
rect 9203 28472 9215 28475
rect 9493 28475 9551 28481
rect 9493 28472 9505 28475
rect 9203 28444 9505 28472
rect 9203 28441 9215 28444
rect 9157 28435 9215 28441
rect 9493 28441 9505 28444
rect 9539 28441 9551 28475
rect 9493 28435 9551 28441
rect 9600 28416 9628 28503
rect 11164 28472 11192 28503
rect 11606 28500 11612 28512
rect 11664 28500 11670 28552
rect 11974 28500 11980 28552
rect 12032 28500 12038 28552
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 13173 28543 13231 28549
rect 13173 28540 13185 28543
rect 12860 28512 13185 28540
rect 12860 28500 12866 28512
rect 13173 28509 13185 28512
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28509 13415 28543
rect 13357 28503 13415 28509
rect 14369 28543 14427 28549
rect 14369 28509 14381 28543
rect 14415 28540 14427 28543
rect 16316 28540 16344 28580
rect 18046 28568 18052 28580
rect 18104 28568 18110 28620
rect 20070 28568 20076 28620
rect 20128 28568 20134 28620
rect 20456 28608 20484 28648
rect 27540 28648 27997 28676
rect 20990 28608 20996 28620
rect 20456 28580 20996 28608
rect 14415 28512 16344 28540
rect 14415 28509 14427 28512
rect 14369 28503 14427 28509
rect 13372 28472 13400 28503
rect 16390 28500 16396 28552
rect 16448 28500 16454 28552
rect 16666 28500 16672 28552
rect 16724 28500 16730 28552
rect 18506 28500 18512 28552
rect 18564 28500 18570 28552
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28540 19855 28543
rect 20088 28540 20116 28568
rect 19843 28512 20116 28540
rect 19843 28509 19855 28512
rect 19797 28503 19855 28509
rect 20162 28500 20168 28552
rect 20220 28500 20226 28552
rect 20355 28543 20413 28549
rect 20355 28509 20367 28543
rect 20401 28540 20413 28543
rect 20456 28540 20484 28580
rect 20990 28568 20996 28580
rect 21048 28568 21054 28620
rect 22738 28568 22744 28620
rect 22796 28568 22802 28620
rect 23842 28568 23848 28620
rect 23900 28608 23906 28620
rect 27540 28617 27568 28648
rect 27985 28645 27997 28648
rect 28031 28645 28043 28679
rect 27985 28639 28043 28645
rect 27525 28611 27583 28617
rect 23900 28580 24256 28608
rect 23900 28568 23906 28580
rect 20401 28512 20484 28540
rect 20533 28543 20591 28549
rect 20401 28509 20413 28512
rect 20355 28503 20413 28509
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20806 28540 20812 28552
rect 20579 28512 20812 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 20806 28500 20812 28512
rect 20864 28500 20870 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 20947 28512 21588 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 16684 28472 16712 28500
rect 19334 28472 19340 28484
rect 11164 28444 12434 28472
rect 13372 28444 16712 28472
rect 16868 28444 19340 28472
rect 8754 28404 8760 28416
rect 8128 28376 8760 28404
rect 8754 28364 8760 28376
rect 8812 28364 8818 28416
rect 9582 28364 9588 28416
rect 9640 28364 9646 28416
rect 12066 28364 12072 28416
rect 12124 28364 12130 28416
rect 12250 28364 12256 28416
rect 12308 28364 12314 28416
rect 12406 28404 12434 28444
rect 16868 28404 16896 28444
rect 19334 28432 19340 28444
rect 19392 28432 19398 28484
rect 20073 28475 20131 28481
rect 20073 28441 20085 28475
rect 20119 28472 20131 28475
rect 20180 28472 20208 28500
rect 20441 28475 20499 28481
rect 20441 28472 20453 28475
rect 20119 28444 20453 28472
rect 20119 28441 20131 28444
rect 20073 28435 20131 28441
rect 20441 28441 20453 28444
rect 20487 28441 20499 28475
rect 20441 28435 20499 28441
rect 21560 28416 21588 28512
rect 23014 28500 23020 28552
rect 23072 28500 23078 28552
rect 23937 28543 23995 28549
rect 23937 28540 23949 28543
rect 23308 28512 23949 28540
rect 21726 28432 21732 28484
rect 21784 28472 21790 28484
rect 23308 28472 23336 28512
rect 23937 28509 23949 28512
rect 23983 28540 23995 28543
rect 24026 28540 24032 28552
rect 23983 28512 24032 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 24026 28500 24032 28512
rect 24084 28500 24090 28552
rect 24228 28549 24256 28580
rect 27525 28577 27537 28611
rect 27571 28577 27583 28611
rect 27525 28571 27583 28577
rect 27801 28611 27859 28617
rect 27801 28577 27813 28611
rect 27847 28608 27859 28611
rect 30116 28608 30144 28716
rect 32582 28704 32588 28716
rect 32640 28704 32646 28756
rect 33962 28704 33968 28756
rect 34020 28704 34026 28756
rect 36906 28704 36912 28756
rect 36964 28744 36970 28756
rect 37369 28747 37427 28753
rect 37369 28744 37381 28747
rect 36964 28716 37381 28744
rect 36964 28704 36970 28716
rect 37369 28713 37381 28716
rect 37415 28744 37427 28747
rect 37918 28744 37924 28756
rect 37415 28716 37924 28744
rect 37415 28713 37427 28716
rect 37369 28707 37427 28713
rect 37918 28704 37924 28716
rect 37976 28704 37982 28756
rect 42153 28747 42211 28753
rect 42153 28713 42165 28747
rect 42199 28744 42211 28747
rect 42886 28744 42892 28756
rect 42199 28716 42892 28744
rect 42199 28713 42211 28716
rect 42153 28707 42211 28713
rect 42886 28704 42892 28716
rect 42944 28704 42950 28756
rect 31570 28636 31576 28688
rect 31628 28676 31634 28688
rect 31628 28648 31708 28676
rect 31628 28636 31634 28648
rect 27847 28580 29040 28608
rect 27847 28577 27859 28580
rect 27801 28571 27859 28577
rect 24213 28543 24271 28549
rect 24213 28509 24225 28543
rect 24259 28509 24271 28543
rect 24213 28503 24271 28509
rect 26234 28500 26240 28552
rect 26292 28540 26298 28552
rect 27430 28540 27436 28552
rect 26292 28512 27436 28540
rect 26292 28500 26298 28512
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 29012 28549 29040 28580
rect 29196 28580 30144 28608
rect 27893 28543 27951 28549
rect 27893 28540 27905 28543
rect 27632 28512 27905 28540
rect 24121 28475 24179 28481
rect 24121 28472 24133 28475
rect 21784 28444 23336 28472
rect 23676 28444 24133 28472
rect 21784 28432 21790 28444
rect 12406 28376 16896 28404
rect 16942 28364 16948 28416
rect 17000 28364 17006 28416
rect 17954 28364 17960 28416
rect 18012 28364 18018 28416
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 19978 28404 19984 28416
rect 19935 28376 19984 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 21542 28364 21548 28416
rect 21600 28364 21606 28416
rect 22094 28364 22100 28416
rect 22152 28404 22158 28416
rect 22189 28407 22247 28413
rect 22189 28404 22201 28407
rect 22152 28376 22201 28404
rect 22152 28364 22158 28376
rect 22189 28373 22201 28376
rect 22235 28373 22247 28407
rect 22189 28367 22247 28373
rect 22554 28364 22560 28416
rect 22612 28364 22618 28416
rect 23676 28413 23704 28444
rect 24121 28441 24133 28444
rect 24167 28441 24179 28475
rect 24121 28435 24179 28441
rect 27632 28416 27660 28512
rect 27893 28509 27905 28512
rect 27939 28509 27951 28543
rect 27893 28503 27951 28509
rect 28077 28543 28135 28549
rect 28077 28509 28089 28543
rect 28123 28509 28135 28543
rect 28077 28503 28135 28509
rect 28997 28543 29055 28549
rect 28997 28509 29009 28543
rect 29043 28509 29055 28543
rect 28997 28503 29055 28509
rect 28092 28472 28120 28503
rect 29196 28484 29224 28580
rect 29914 28500 29920 28552
rect 29972 28500 29978 28552
rect 30116 28549 30144 28580
rect 31202 28568 31208 28620
rect 31260 28568 31266 28620
rect 31680 28617 31708 28648
rect 32122 28636 32128 28688
rect 32180 28676 32186 28688
rect 32180 28648 33088 28676
rect 32180 28636 32186 28648
rect 31665 28611 31723 28617
rect 31665 28577 31677 28611
rect 31711 28577 31723 28611
rect 31665 28571 31723 28577
rect 32950 28568 32956 28620
rect 33008 28568 33014 28620
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 30377 28543 30435 28549
rect 30377 28509 30389 28543
rect 30423 28540 30435 28543
rect 30469 28543 30527 28549
rect 30469 28540 30481 28543
rect 30423 28512 30481 28540
rect 30423 28509 30435 28512
rect 30377 28503 30435 28509
rect 30469 28509 30481 28512
rect 30515 28509 30527 28543
rect 30469 28503 30527 28509
rect 30558 28500 30564 28552
rect 30616 28540 30622 28552
rect 31018 28540 31024 28552
rect 30616 28512 31024 28540
rect 30616 28500 30622 28512
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 31573 28543 31631 28549
rect 31573 28509 31585 28543
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 31849 28543 31907 28549
rect 31849 28509 31861 28543
rect 31895 28540 31907 28543
rect 32033 28543 32091 28549
rect 32033 28540 32045 28543
rect 31895 28512 32045 28540
rect 31895 28509 31907 28512
rect 31849 28503 31907 28509
rect 32033 28509 32045 28512
rect 32079 28509 32091 28543
rect 32033 28503 32091 28509
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 27908 28444 28120 28472
rect 27908 28416 27936 28444
rect 29178 28432 29184 28484
rect 29236 28432 29242 28484
rect 30009 28475 30067 28481
rect 30009 28441 30021 28475
rect 30055 28441 30067 28475
rect 30009 28435 30067 28441
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28404 22707 28407
rect 23661 28407 23719 28413
rect 23661 28404 23673 28407
rect 22695 28376 23673 28404
rect 22695 28373 22707 28376
rect 22649 28367 22707 28373
rect 23661 28373 23673 28376
rect 23707 28373 23719 28407
rect 23661 28367 23719 28373
rect 23750 28364 23756 28416
rect 23808 28364 23814 28416
rect 27614 28364 27620 28416
rect 27672 28364 27678 28416
rect 27890 28364 27896 28416
rect 27948 28364 27954 28416
rect 29730 28364 29736 28416
rect 29788 28364 29794 28416
rect 30024 28404 30052 28435
rect 30190 28432 30196 28484
rect 30248 28481 30254 28484
rect 30248 28475 30297 28481
rect 30248 28441 30251 28475
rect 30285 28472 30297 28475
rect 31386 28472 31392 28484
rect 30285 28444 31392 28472
rect 30285 28441 30297 28444
rect 30248 28435 30297 28441
rect 30248 28432 30254 28435
rect 31386 28432 31392 28444
rect 31444 28432 31450 28484
rect 30466 28404 30472 28416
rect 30024 28376 30472 28404
rect 30466 28364 30472 28376
rect 30524 28364 30530 28416
rect 31588 28404 31616 28503
rect 31754 28432 31760 28484
rect 31812 28472 31818 28484
rect 32232 28472 32260 28503
rect 32306 28500 32312 28552
rect 32364 28500 32370 28552
rect 33060 28549 33088 28648
rect 35897 28611 35955 28617
rect 35897 28577 35909 28611
rect 35943 28608 35955 28611
rect 35986 28608 35992 28620
rect 35943 28580 35992 28608
rect 35943 28577 35955 28580
rect 35897 28571 35955 28577
rect 35986 28568 35992 28580
rect 36044 28568 36050 28620
rect 40405 28611 40463 28617
rect 40405 28577 40417 28611
rect 40451 28608 40463 28611
rect 40770 28608 40776 28620
rect 40451 28580 40776 28608
rect 40451 28577 40463 28580
rect 40405 28571 40463 28577
rect 40770 28568 40776 28580
rect 40828 28608 40834 28620
rect 41966 28608 41972 28620
rect 40828 28580 41972 28608
rect 40828 28568 40834 28580
rect 41966 28568 41972 28580
rect 42024 28608 42030 28620
rect 42024 28580 42288 28608
rect 42024 28568 42030 28580
rect 33045 28543 33103 28549
rect 33045 28509 33057 28543
rect 33091 28509 33103 28543
rect 33045 28503 33103 28509
rect 34057 28543 34115 28549
rect 34057 28509 34069 28543
rect 34103 28540 34115 28543
rect 34103 28512 34376 28540
rect 34103 28509 34115 28512
rect 34057 28503 34115 28509
rect 31812 28444 32260 28472
rect 32493 28475 32551 28481
rect 31812 28432 31818 28444
rect 32493 28441 32505 28475
rect 32539 28472 32551 28475
rect 33502 28472 33508 28484
rect 32539 28444 33508 28472
rect 32539 28441 32551 28444
rect 32493 28435 32551 28441
rect 33502 28432 33508 28444
rect 33560 28432 33566 28484
rect 34348 28416 34376 28512
rect 35342 28500 35348 28552
rect 35400 28540 35406 28552
rect 35621 28543 35679 28549
rect 35621 28540 35633 28543
rect 35400 28512 35633 28540
rect 35400 28500 35406 28512
rect 35621 28509 35633 28512
rect 35667 28509 35679 28543
rect 35621 28503 35679 28509
rect 37826 28500 37832 28552
rect 37884 28540 37890 28552
rect 38473 28543 38531 28549
rect 38473 28540 38485 28543
rect 37884 28512 38485 28540
rect 37884 28500 37890 28512
rect 38473 28509 38485 28512
rect 38519 28540 38531 28543
rect 38562 28540 38568 28552
rect 38519 28512 38568 28540
rect 38519 28509 38531 28512
rect 38473 28503 38531 28509
rect 38562 28500 38568 28512
rect 38620 28500 38626 28552
rect 39669 28543 39727 28549
rect 39669 28509 39681 28543
rect 39715 28540 39727 28543
rect 39942 28540 39948 28552
rect 39715 28512 39948 28540
rect 39715 28509 39727 28512
rect 39669 28503 39727 28509
rect 39942 28500 39948 28512
rect 40000 28500 40006 28552
rect 42260 28549 42288 28580
rect 43070 28568 43076 28620
rect 43128 28608 43134 28620
rect 44269 28611 44327 28617
rect 44269 28608 44281 28611
rect 43128 28580 44281 28608
rect 43128 28568 43134 28580
rect 44269 28577 44281 28580
rect 44315 28577 44327 28611
rect 44269 28571 44327 28577
rect 42245 28543 42303 28549
rect 42245 28509 42257 28543
rect 42291 28509 42303 28543
rect 42245 28503 42303 28509
rect 35986 28432 35992 28484
rect 36044 28472 36050 28484
rect 36044 28444 36386 28472
rect 36044 28432 36050 28444
rect 40678 28432 40684 28484
rect 40736 28432 40742 28484
rect 41138 28432 41144 28484
rect 41196 28432 41202 28484
rect 42260 28472 42288 28503
rect 42260 28444 42380 28472
rect 42352 28416 42380 28444
rect 42426 28432 42432 28484
rect 42484 28472 42490 28484
rect 42521 28475 42579 28481
rect 42521 28472 42533 28475
rect 42484 28444 42533 28472
rect 42484 28432 42490 28444
rect 42521 28441 42533 28444
rect 42567 28441 42579 28475
rect 42521 28435 42579 28441
rect 42978 28432 42984 28484
rect 43036 28432 43042 28484
rect 32030 28404 32036 28416
rect 31588 28376 32036 28404
rect 32030 28364 32036 28376
rect 32088 28364 32094 28416
rect 32674 28364 32680 28416
rect 32732 28364 32738 28416
rect 34330 28364 34336 28416
rect 34388 28364 34394 28416
rect 37829 28407 37887 28413
rect 37829 28373 37841 28407
rect 37875 28404 37887 28407
rect 38194 28404 38200 28416
rect 37875 28376 38200 28404
rect 37875 28373 37887 28376
rect 37829 28367 37887 28373
rect 38194 28364 38200 28376
rect 38252 28364 38258 28416
rect 38838 28364 38844 28416
rect 38896 28404 38902 28416
rect 39025 28407 39083 28413
rect 39025 28404 39037 28407
rect 38896 28376 39037 28404
rect 38896 28364 38902 28376
rect 39025 28373 39037 28376
rect 39071 28373 39083 28407
rect 39025 28367 39083 28373
rect 42334 28364 42340 28416
rect 42392 28364 42398 28416
rect 1104 28314 44620 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 44620 28314
rect 1104 28240 44620 28262
rect 5905 28203 5963 28209
rect 5905 28200 5917 28203
rect 5368 28172 5917 28200
rect 5368 28073 5396 28172
rect 5905 28169 5917 28172
rect 5951 28169 5963 28203
rect 5905 28163 5963 28169
rect 8573 28203 8631 28209
rect 8573 28169 8585 28203
rect 8619 28169 8631 28203
rect 8573 28163 8631 28169
rect 8741 28203 8799 28209
rect 8741 28169 8753 28203
rect 8787 28200 8799 28203
rect 9030 28200 9036 28212
rect 8787 28172 9036 28200
rect 8787 28169 8799 28172
rect 8741 28163 8799 28169
rect 5736 28104 6132 28132
rect 5736 28086 5764 28104
rect 5353 28067 5411 28073
rect 5353 28033 5365 28067
rect 5399 28033 5411 28067
rect 5353 28027 5411 28033
rect 5534 28024 5540 28076
rect 5592 28024 5598 28076
rect 5644 28073 5764 28086
rect 6104 28076 6132 28104
rect 7098 28092 7104 28144
rect 7156 28092 7162 28144
rect 7300 28104 7512 28132
rect 5629 28067 5764 28073
rect 5629 28033 5641 28067
rect 5675 28058 5764 28067
rect 5675 28033 5687 28058
rect 5629 28027 5687 28033
rect 5810 28024 5816 28076
rect 5868 28073 5874 28076
rect 5868 28067 5883 28073
rect 5871 28033 5883 28067
rect 5868 28027 5883 28033
rect 5868 28024 5874 28027
rect 6086 28024 6092 28076
rect 6144 28024 6150 28076
rect 6181 28067 6239 28073
rect 6181 28033 6193 28067
rect 6227 28064 6239 28067
rect 6365 28067 6423 28073
rect 6365 28064 6377 28067
rect 6227 28036 6377 28064
rect 6227 28033 6239 28036
rect 6181 28027 6239 28033
rect 6365 28033 6377 28036
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 7009 28067 7067 28073
rect 7009 28033 7021 28067
rect 7055 28064 7067 28067
rect 7116 28064 7144 28092
rect 7300 28073 7328 28104
rect 7484 28076 7512 28104
rect 7834 28092 7840 28144
rect 7892 28092 7898 28144
rect 7055 28036 7144 28064
rect 7285 28067 7343 28073
rect 7055 28033 7067 28036
rect 7009 28027 7067 28033
rect 7285 28033 7297 28067
rect 7331 28033 7343 28067
rect 7285 28027 7343 28033
rect 7377 28067 7435 28073
rect 7377 28033 7389 28067
rect 7423 28033 7435 28067
rect 7377 28027 7435 28033
rect 5905 27999 5963 28005
rect 5905 27965 5917 27999
rect 5951 27996 5963 27999
rect 7101 27999 7159 28005
rect 7101 27996 7113 27999
rect 5951 27968 7113 27996
rect 5951 27965 5963 27968
rect 5905 27959 5963 27965
rect 7101 27965 7113 27968
rect 7147 27965 7159 27999
rect 7101 27959 7159 27965
rect 5813 27931 5871 27937
rect 5813 27897 5825 27931
rect 5859 27928 5871 27931
rect 6362 27928 6368 27940
rect 5859 27900 6368 27928
rect 5859 27897 5871 27900
rect 5813 27891 5871 27897
rect 6362 27888 6368 27900
rect 6420 27888 6426 27940
rect 7116 27928 7144 27959
rect 7190 27956 7196 28008
rect 7248 27996 7254 28008
rect 7392 27996 7420 28027
rect 7466 28024 7472 28076
rect 7524 28024 7530 28076
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28064 8355 28067
rect 8588 28064 8616 28163
rect 9030 28160 9036 28172
rect 9088 28200 9094 28212
rect 9582 28200 9588 28212
rect 9088 28172 9588 28200
rect 9088 28160 9094 28172
rect 9582 28160 9588 28172
rect 9640 28160 9646 28212
rect 11517 28203 11575 28209
rect 11517 28169 11529 28203
rect 11563 28169 11575 28203
rect 11517 28163 11575 28169
rect 11885 28203 11943 28209
rect 11885 28169 11897 28203
rect 11931 28200 11943 28203
rect 12250 28200 12256 28212
rect 11931 28172 12256 28200
rect 11931 28169 11943 28172
rect 11885 28163 11943 28169
rect 8941 28135 8999 28141
rect 8941 28101 8953 28135
rect 8987 28101 8999 28135
rect 8941 28095 8999 28101
rect 8343 28036 8616 28064
rect 8343 28033 8355 28036
rect 8297 28027 8355 28033
rect 8754 28024 8760 28076
rect 8812 28064 8818 28076
rect 8956 28064 8984 28095
rect 9398 28092 9404 28144
rect 9456 28132 9462 28144
rect 9456 28104 9628 28132
rect 9456 28092 9462 28104
rect 8812 28036 8984 28064
rect 9217 28067 9275 28073
rect 8812 28024 8818 28036
rect 9217 28033 9229 28067
rect 9263 28033 9275 28067
rect 9217 28027 9275 28033
rect 9232 27996 9260 28027
rect 9490 28024 9496 28076
rect 9548 28024 9554 28076
rect 9600 28073 9628 28104
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28033 9643 28067
rect 9585 28027 9643 28033
rect 9674 28024 9680 28076
rect 9732 28024 9738 28076
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28064 9919 28067
rect 10318 28064 10324 28076
rect 9907 28036 10324 28064
rect 9907 28033 9919 28036
rect 9861 28027 9919 28033
rect 9876 27996 9904 28027
rect 10318 28024 10324 28036
rect 10376 28024 10382 28076
rect 11333 28067 11391 28073
rect 11333 28033 11345 28067
rect 11379 28064 11391 28067
rect 11532 28064 11560 28163
rect 12250 28160 12256 28172
rect 12308 28160 12314 28212
rect 12434 28160 12440 28212
rect 12492 28160 12498 28212
rect 13909 28203 13967 28209
rect 13909 28169 13921 28203
rect 13955 28169 13967 28203
rect 13909 28163 13967 28169
rect 15749 28203 15807 28209
rect 15749 28169 15761 28203
rect 15795 28200 15807 28203
rect 16390 28200 16396 28212
rect 15795 28172 16396 28200
rect 15795 28169 15807 28172
rect 15749 28163 15807 28169
rect 11606 28092 11612 28144
rect 11664 28132 11670 28144
rect 11977 28135 12035 28141
rect 11977 28132 11989 28135
rect 11664 28104 11989 28132
rect 11664 28092 11670 28104
rect 11977 28101 11989 28104
rect 12023 28101 12035 28135
rect 11977 28095 12035 28101
rect 12066 28092 12072 28144
rect 12124 28132 12130 28144
rect 12805 28135 12863 28141
rect 12805 28132 12817 28135
rect 12124 28104 12817 28132
rect 12124 28092 12130 28104
rect 12805 28101 12817 28104
rect 12851 28101 12863 28135
rect 13924 28132 13952 28163
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 16942 28200 16948 28212
rect 16776 28172 16948 28200
rect 14277 28135 14335 28141
rect 14277 28132 14289 28135
rect 13924 28104 14289 28132
rect 12805 28095 12863 28101
rect 14277 28101 14289 28104
rect 14323 28101 14335 28135
rect 15654 28132 15660 28144
rect 15502 28104 15660 28132
rect 14277 28095 14335 28101
rect 15654 28092 15660 28104
rect 15712 28092 15718 28144
rect 11379 28036 11560 28064
rect 11379 28033 11391 28036
rect 11333 28027 11391 28033
rect 7248 27968 8432 27996
rect 9232 27968 9904 27996
rect 7248 27956 7254 27968
rect 8404 27940 8432 27968
rect 7834 27928 7840 27940
rect 7116 27900 7840 27928
rect 7834 27888 7840 27900
rect 7892 27888 7898 27940
rect 8386 27888 8392 27940
rect 8444 27928 8450 27940
rect 11624 27928 11652 28092
rect 12618 28073 12624 28076
rect 12616 28027 12624 28073
rect 12618 28024 12624 28027
rect 12676 28024 12682 28076
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 12161 27999 12219 28005
rect 12161 27965 12173 27999
rect 12207 27996 12219 27999
rect 12526 27996 12532 28008
rect 12207 27968 12532 27996
rect 12207 27965 12219 27968
rect 12161 27959 12219 27965
rect 12526 27956 12532 27968
rect 12584 27956 12590 28008
rect 12728 27996 12756 28027
rect 12986 28024 12992 28076
rect 13044 28024 13050 28076
rect 13078 28024 13084 28076
rect 13136 28024 13142 28076
rect 13725 28067 13783 28073
rect 13725 28033 13737 28067
rect 13771 28064 13783 28067
rect 13906 28064 13912 28076
rect 13771 28036 13912 28064
rect 13771 28033 13783 28036
rect 13725 28027 13783 28033
rect 13906 28024 13912 28036
rect 13964 28024 13970 28076
rect 16408 28073 16436 28160
rect 16776 28073 16804 28172
rect 16942 28160 16948 28172
rect 17000 28160 17006 28212
rect 17126 28160 17132 28212
rect 17184 28160 17190 28212
rect 17497 28203 17555 28209
rect 17497 28169 17509 28203
rect 17543 28200 17555 28203
rect 17954 28200 17960 28212
rect 17543 28172 17960 28200
rect 17543 28169 17555 28172
rect 17497 28163 17555 28169
rect 17954 28160 17960 28172
rect 18012 28200 18018 28212
rect 18141 28203 18199 28209
rect 18141 28200 18153 28203
rect 18012 28172 18153 28200
rect 18012 28160 18018 28172
rect 18141 28169 18153 28172
rect 18187 28169 18199 28203
rect 18141 28163 18199 28169
rect 19889 28203 19947 28209
rect 19889 28169 19901 28203
rect 19935 28200 19947 28203
rect 20070 28200 20076 28212
rect 19935 28172 20076 28200
rect 19935 28169 19947 28172
rect 19889 28163 19947 28169
rect 20070 28160 20076 28172
rect 20128 28160 20134 28212
rect 20806 28160 20812 28212
rect 20864 28200 20870 28212
rect 21545 28203 21603 28209
rect 21545 28200 21557 28203
rect 20864 28172 21557 28200
rect 20864 28160 20870 28172
rect 21545 28169 21557 28172
rect 21591 28169 21603 28203
rect 21545 28163 21603 28169
rect 21821 28203 21879 28209
rect 21821 28169 21833 28203
rect 21867 28200 21879 28203
rect 23014 28200 23020 28212
rect 21867 28172 23020 28200
rect 21867 28169 21879 28172
rect 21821 28163 21879 28169
rect 23014 28160 23020 28172
rect 23072 28160 23078 28212
rect 23106 28160 23112 28212
rect 23164 28200 23170 28212
rect 23658 28200 23664 28212
rect 23164 28172 23664 28200
rect 23164 28160 23170 28172
rect 23658 28160 23664 28172
rect 23716 28160 23722 28212
rect 23750 28160 23756 28212
rect 23808 28160 23814 28212
rect 25314 28160 25320 28212
rect 25372 28160 25378 28212
rect 26234 28160 26240 28212
rect 26292 28200 26298 28212
rect 26421 28203 26479 28209
rect 26421 28200 26433 28203
rect 26292 28172 26433 28200
rect 26292 28160 26298 28172
rect 26421 28169 26433 28172
rect 26467 28169 26479 28203
rect 29730 28200 29736 28212
rect 26421 28163 26479 28169
rect 28920 28172 29736 28200
rect 17144 28132 17172 28160
rect 23124 28132 23152 28160
rect 17144 28104 17632 28132
rect 22862 28104 23152 28132
rect 23293 28135 23351 28141
rect 16393 28067 16451 28073
rect 16393 28033 16405 28067
rect 16439 28033 16451 28067
rect 16393 28027 16451 28033
rect 16761 28067 16819 28073
rect 16761 28033 16773 28067
rect 16807 28033 16819 28067
rect 16761 28027 16819 28033
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 12728 27968 13032 27996
rect 8444 27900 11652 27928
rect 8444 27888 8450 27900
rect 13004 27872 13032 27968
rect 13814 27956 13820 28008
rect 13872 27996 13878 28008
rect 14001 27999 14059 28005
rect 14001 27996 14013 27999
rect 13872 27968 14013 27996
rect 13872 27956 13878 27968
rect 14001 27965 14013 27968
rect 14047 27965 14059 27999
rect 14001 27959 14059 27965
rect 16666 27956 16672 28008
rect 16724 27996 16730 28008
rect 16868 27996 16896 28027
rect 17034 28024 17040 28076
rect 17092 28064 17098 28076
rect 17313 28067 17371 28073
rect 17313 28064 17325 28067
rect 17092 28036 17325 28064
rect 17092 28024 17098 28036
rect 17313 28033 17325 28036
rect 17359 28064 17371 28067
rect 17494 28064 17500 28076
rect 17359 28036 17500 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 17494 28024 17500 28036
rect 17552 28024 17558 28076
rect 17604 28073 17632 28104
rect 23293 28101 23305 28135
rect 23339 28132 23351 28135
rect 23768 28132 23796 28160
rect 23339 28104 23796 28132
rect 25332 28132 25360 28160
rect 28920 28141 28948 28172
rect 29730 28160 29736 28172
rect 29788 28160 29794 28212
rect 29914 28160 29920 28212
rect 29972 28200 29978 28212
rect 29972 28172 30420 28200
rect 29972 28160 29978 28172
rect 28905 28135 28963 28141
rect 25332 28104 25438 28132
rect 23339 28101 23351 28104
rect 23293 28095 23351 28101
rect 28905 28101 28917 28135
rect 28951 28101 28963 28135
rect 28905 28095 28963 28101
rect 29362 28092 29368 28144
rect 29420 28092 29426 28144
rect 30392 28132 30420 28172
rect 30466 28160 30472 28212
rect 30524 28160 30530 28212
rect 30929 28203 30987 28209
rect 30929 28200 30941 28203
rect 30576 28172 30941 28200
rect 30576 28132 30604 28172
rect 30929 28169 30941 28172
rect 30975 28169 30987 28203
rect 30929 28163 30987 28169
rect 31662 28160 31668 28212
rect 31720 28200 31726 28212
rect 31757 28203 31815 28209
rect 31757 28200 31769 28203
rect 31720 28172 31769 28200
rect 31720 28160 31726 28172
rect 31757 28169 31769 28172
rect 31803 28169 31815 28203
rect 31757 28163 31815 28169
rect 32217 28203 32275 28209
rect 32217 28169 32229 28203
rect 32263 28200 32275 28203
rect 32306 28200 32312 28212
rect 32263 28172 32312 28200
rect 32263 28169 32275 28172
rect 32217 28163 32275 28169
rect 32306 28160 32312 28172
rect 32364 28160 32370 28212
rect 32950 28160 32956 28212
rect 33008 28160 33014 28212
rect 35713 28203 35771 28209
rect 35713 28169 35725 28203
rect 35759 28200 35771 28203
rect 36538 28200 36544 28212
rect 35759 28172 36544 28200
rect 35759 28169 35771 28172
rect 35713 28163 35771 28169
rect 36538 28160 36544 28172
rect 36596 28160 36602 28212
rect 38194 28200 38200 28212
rect 37200 28172 38200 28200
rect 30834 28141 30840 28144
rect 30392 28104 30604 28132
rect 30653 28135 30711 28141
rect 30653 28101 30665 28135
rect 30699 28101 30711 28135
rect 30653 28095 30711 28101
rect 30818 28135 30840 28141
rect 30818 28101 30830 28135
rect 30818 28095 30840 28101
rect 17589 28067 17647 28073
rect 17589 28033 17601 28067
rect 17635 28033 17647 28067
rect 17589 28027 17647 28033
rect 18049 28067 18107 28073
rect 18049 28033 18061 28067
rect 18095 28064 18107 28067
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 18095 28036 18521 28064
rect 18095 28033 18107 28036
rect 18049 28027 18107 28033
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20070 28064 20076 28076
rect 19935 28036 20076 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 16724 27968 16896 27996
rect 16724 27956 16730 27968
rect 18322 27956 18328 28008
rect 18380 27956 18386 28008
rect 19150 27956 19156 28008
rect 19208 27956 19214 28008
rect 19702 27956 19708 28008
rect 19760 27996 19766 28008
rect 19978 27996 19984 28008
rect 19760 27968 19984 27996
rect 19760 27956 19766 27968
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 20272 27996 20300 28027
rect 20622 28024 20628 28076
rect 20680 28024 20686 28076
rect 21542 28024 21548 28076
rect 21600 28024 21606 28076
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28064 21695 28067
rect 21683 28036 22094 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 21560 27996 21588 28024
rect 20272 27968 21588 27996
rect 21726 27956 21732 28008
rect 21784 27956 21790 28008
rect 22066 27996 22094 28036
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 27338 28024 27344 28076
rect 27396 28024 27402 28076
rect 28074 28024 28080 28076
rect 28132 28024 28138 28076
rect 22554 27996 22560 28008
rect 22066 27968 22560 27996
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 23569 27999 23627 28005
rect 23569 27965 23581 27999
rect 23615 27996 23627 27999
rect 24670 27996 24676 28008
rect 23615 27968 24676 27996
rect 23615 27965 23627 27968
rect 23569 27959 23627 27965
rect 17037 27931 17095 27937
rect 17037 27897 17049 27931
rect 17083 27928 17095 27931
rect 21744 27928 21772 27956
rect 17083 27900 21772 27928
rect 17083 27897 17095 27900
rect 17037 27891 17095 27897
rect 5350 27820 5356 27872
rect 5408 27820 5414 27872
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 7193 27863 7251 27869
rect 7193 27860 7205 27863
rect 5960 27832 7205 27860
rect 5960 27820 5966 27832
rect 7193 27829 7205 27832
rect 7239 27829 7251 27863
rect 7193 27823 7251 27829
rect 7374 27820 7380 27872
rect 7432 27860 7438 27872
rect 7745 27863 7803 27869
rect 7745 27860 7757 27863
rect 7432 27832 7757 27860
rect 7432 27820 7438 27832
rect 7745 27829 7757 27832
rect 7791 27860 7803 27863
rect 8202 27860 8208 27872
rect 7791 27832 8208 27860
rect 7791 27829 7803 27832
rect 7745 27823 7803 27829
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 8478 27820 8484 27872
rect 8536 27820 8542 27872
rect 8757 27863 8815 27869
rect 8757 27829 8769 27863
rect 8803 27860 8815 27863
rect 9033 27863 9091 27869
rect 9033 27860 9045 27863
rect 8803 27832 9045 27860
rect 8803 27829 8815 27832
rect 8757 27823 8815 27829
rect 9033 27829 9045 27832
rect 9079 27829 9091 27863
rect 9033 27823 9091 27829
rect 11146 27820 11152 27872
rect 11204 27820 11210 27872
rect 12986 27820 12992 27872
rect 13044 27820 13050 27872
rect 15838 27820 15844 27872
rect 15896 27820 15902 27872
rect 17126 27820 17132 27872
rect 17184 27820 17190 27872
rect 17218 27820 17224 27872
rect 17276 27860 17282 27872
rect 17681 27863 17739 27869
rect 17681 27860 17693 27863
rect 17276 27832 17693 27860
rect 17276 27820 17282 27832
rect 17681 27829 17693 27832
rect 17727 27829 17739 27863
rect 17681 27823 17739 27829
rect 20165 27863 20223 27869
rect 20165 27829 20177 27863
rect 20211 27860 20223 27863
rect 20533 27863 20591 27869
rect 20533 27860 20545 27863
rect 20211 27832 20545 27860
rect 20211 27829 20223 27832
rect 20165 27823 20223 27829
rect 20533 27829 20545 27832
rect 20579 27829 20591 27863
rect 20533 27823 20591 27829
rect 23290 27820 23296 27872
rect 23348 27860 23354 27872
rect 23584 27860 23612 27959
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 24946 27956 24952 28008
rect 25004 27956 25010 28008
rect 28353 27999 28411 28005
rect 28353 27965 28365 27999
rect 28399 27996 28411 27999
rect 28534 27996 28540 28008
rect 28399 27968 28540 27996
rect 28399 27965 28411 27968
rect 28353 27959 28411 27965
rect 28534 27956 28540 27968
rect 28592 27956 28598 28008
rect 28629 27999 28687 28005
rect 28629 27965 28641 27999
rect 28675 27996 28687 27999
rect 30377 27999 30435 28005
rect 28675 27968 28764 27996
rect 28675 27965 28687 27968
rect 28629 27959 28687 27965
rect 28736 27872 28764 27968
rect 30377 27965 30389 27999
rect 30423 27996 30435 27999
rect 30558 27996 30564 28008
rect 30423 27968 30564 27996
rect 30423 27965 30435 27968
rect 30377 27959 30435 27965
rect 30558 27956 30564 27968
rect 30616 27956 30622 28008
rect 30668 27996 30696 28095
rect 30834 28092 30840 28095
rect 30892 28092 30898 28144
rect 31202 28132 31208 28144
rect 30944 28104 31208 28132
rect 30944 28073 30972 28104
rect 31202 28092 31208 28104
rect 31260 28092 31266 28144
rect 30929 28067 30987 28073
rect 30929 28033 30941 28067
rect 30975 28033 30987 28067
rect 30929 28027 30987 28033
rect 31110 28024 31116 28076
rect 31168 28024 31174 28076
rect 31220 28064 31248 28092
rect 31389 28067 31447 28073
rect 31220 28062 31340 28064
rect 31389 28062 31401 28067
rect 31220 28036 31401 28062
rect 31220 27996 31248 28036
rect 31312 28034 31401 28036
rect 31389 28033 31401 28034
rect 31435 28033 31447 28067
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31389 28027 31447 28033
rect 31588 28036 31769 28064
rect 31588 27996 31616 28036
rect 31757 28033 31769 28036
rect 31803 28033 31815 28067
rect 31757 28027 31815 28033
rect 31938 28024 31944 28076
rect 31996 28024 32002 28076
rect 32030 28024 32036 28076
rect 32088 28064 32094 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 32088 28036 32137 28064
rect 32088 28024 32094 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32306 28024 32312 28076
rect 32364 28024 32370 28076
rect 30668 27968 31248 27996
rect 31496 27968 31616 27996
rect 31665 27999 31723 28005
rect 30576 27928 30604 27956
rect 31496 27928 31524 27968
rect 31665 27965 31677 27999
rect 31711 27996 31723 27999
rect 32048 27996 32076 28024
rect 31711 27968 32076 27996
rect 31711 27965 31723 27968
rect 31665 27959 31723 27965
rect 30576 27900 31524 27928
rect 31573 27931 31631 27937
rect 31573 27897 31585 27931
rect 31619 27928 31631 27931
rect 32968 27928 32996 28160
rect 33870 28132 33876 28144
rect 33336 28104 33876 28132
rect 33336 28073 33364 28104
rect 33870 28092 33876 28104
rect 33928 28092 33934 28144
rect 33321 28067 33379 28073
rect 33321 28033 33333 28067
rect 33367 28033 33379 28067
rect 35529 28067 35587 28073
rect 34730 28036 35388 28064
rect 33321 28027 33379 28033
rect 33594 27956 33600 28008
rect 33652 27956 33658 28008
rect 34330 27956 34336 28008
rect 34388 27996 34394 28008
rect 35069 27999 35127 28005
rect 35069 27996 35081 27999
rect 34388 27968 35081 27996
rect 34388 27956 34394 27968
rect 35069 27965 35081 27968
rect 35115 27965 35127 27999
rect 35069 27959 35127 27965
rect 35360 27937 35388 28036
rect 35529 28033 35541 28067
rect 35575 28064 35587 28067
rect 35575 28036 35756 28064
rect 35575 28033 35587 28036
rect 35529 28027 35587 28033
rect 35728 28008 35756 28036
rect 35894 28024 35900 28076
rect 35952 28024 35958 28076
rect 35989 28067 36047 28073
rect 35989 28033 36001 28067
rect 36035 28033 36047 28067
rect 35989 28027 36047 28033
rect 36081 28067 36139 28073
rect 36081 28033 36093 28067
rect 36127 28064 36139 28067
rect 36170 28064 36176 28076
rect 36127 28036 36176 28064
rect 36127 28033 36139 28036
rect 36081 28027 36139 28033
rect 35710 27956 35716 28008
rect 35768 27956 35774 28008
rect 36004 27996 36032 28027
rect 36170 28024 36176 28036
rect 36228 28024 36234 28076
rect 36265 28067 36323 28073
rect 36265 28033 36277 28067
rect 36311 28064 36323 28067
rect 37200 28064 37228 28172
rect 38194 28160 38200 28172
rect 38252 28160 38258 28212
rect 40678 28160 40684 28212
rect 40736 28200 40742 28212
rect 41141 28203 41199 28209
rect 41141 28200 41153 28203
rect 40736 28172 41153 28200
rect 40736 28160 40742 28172
rect 41141 28169 41153 28172
rect 41187 28169 41199 28203
rect 41141 28163 41199 28169
rect 37274 28092 37280 28144
rect 37332 28132 37338 28144
rect 38010 28132 38016 28144
rect 37332 28104 38016 28132
rect 37332 28092 37338 28104
rect 38010 28092 38016 28104
rect 38068 28092 38074 28144
rect 40494 28092 40500 28144
rect 40552 28132 40558 28144
rect 40589 28135 40647 28141
rect 40589 28132 40601 28135
rect 40552 28104 40601 28132
rect 40552 28092 40558 28104
rect 40589 28101 40601 28104
rect 40635 28101 40647 28135
rect 40589 28095 40647 28101
rect 39298 28064 39304 28076
rect 36311 28036 37228 28064
rect 38580 28036 39304 28064
rect 36311 28033 36323 28036
rect 36265 28027 36323 28033
rect 36906 27996 36912 28008
rect 36004 27968 36912 27996
rect 36906 27956 36912 27968
rect 36964 27956 36970 28008
rect 37277 27999 37335 28005
rect 37277 27965 37289 27999
rect 37323 27965 37335 27999
rect 37277 27959 37335 27965
rect 31619 27900 32996 27928
rect 35345 27931 35403 27937
rect 31619 27897 31631 27900
rect 31573 27891 31631 27897
rect 35345 27897 35357 27931
rect 35391 27928 35403 27931
rect 35986 27928 35992 27940
rect 35391 27900 35992 27928
rect 35391 27897 35403 27900
rect 35345 27891 35403 27897
rect 35986 27888 35992 27900
rect 36044 27928 36050 27940
rect 37182 27928 37188 27940
rect 36044 27900 37188 27928
rect 36044 27888 36050 27900
rect 37182 27888 37188 27900
rect 37240 27888 37246 27940
rect 23348 27832 23612 27860
rect 23348 27820 23354 27832
rect 24578 27820 24584 27872
rect 24636 27820 24642 27872
rect 27890 27820 27896 27872
rect 27948 27820 27954 27872
rect 28718 27820 28724 27872
rect 28776 27820 28782 27872
rect 30834 27820 30840 27872
rect 30892 27860 30898 27872
rect 31110 27860 31116 27872
rect 30892 27832 31116 27860
rect 30892 27820 30898 27832
rect 31110 27820 31116 27832
rect 31168 27860 31174 27872
rect 31481 27863 31539 27869
rect 31481 27860 31493 27863
rect 31168 27832 31493 27860
rect 31168 27820 31174 27832
rect 31481 27829 31493 27832
rect 31527 27860 31539 27863
rect 31754 27860 31760 27872
rect 31527 27832 31760 27860
rect 31527 27829 31539 27832
rect 31481 27823 31539 27829
rect 31754 27820 31760 27832
rect 31812 27820 31818 27872
rect 34698 27820 34704 27872
rect 34756 27860 34762 27872
rect 36357 27863 36415 27869
rect 36357 27860 36369 27863
rect 34756 27832 36369 27860
rect 34756 27820 34762 27832
rect 36357 27829 36369 27832
rect 36403 27829 36415 27863
rect 37292 27860 37320 27959
rect 37550 27956 37556 28008
rect 37608 27956 37614 28008
rect 38010 27956 38016 28008
rect 38068 27996 38074 28008
rect 38580 27996 38608 28036
rect 39298 28024 39304 28036
rect 39356 28064 39362 28076
rect 39356 28036 39514 28064
rect 39356 28024 39362 28036
rect 42518 28024 42524 28076
rect 42576 28024 42582 28076
rect 38068 27968 38608 27996
rect 39025 27999 39083 28005
rect 38068 27956 38074 27968
rect 39025 27965 39037 27999
rect 39071 27996 39083 27999
rect 40218 27996 40224 28008
rect 39071 27968 40224 27996
rect 39071 27965 39083 27968
rect 39025 27959 39083 27965
rect 38562 27888 38568 27940
rect 38620 27928 38626 27940
rect 39040 27928 39068 27959
rect 40218 27956 40224 27968
rect 40276 27956 40282 28008
rect 40862 27956 40868 28008
rect 40920 27956 40926 28008
rect 41690 27956 41696 28008
rect 41748 27956 41754 28008
rect 38620 27900 39068 27928
rect 38620 27888 38626 27900
rect 38102 27860 38108 27872
rect 37292 27832 38108 27860
rect 36357 27823 36415 27829
rect 38102 27820 38108 27832
rect 38160 27820 38166 27872
rect 39117 27863 39175 27869
rect 39117 27829 39129 27863
rect 39163 27860 39175 27863
rect 39206 27860 39212 27872
rect 39163 27832 39212 27860
rect 39163 27829 39175 27832
rect 39117 27823 39175 27829
rect 39206 27820 39212 27832
rect 39264 27820 39270 27872
rect 40034 27820 40040 27872
rect 40092 27860 40098 27872
rect 40880 27860 40908 27956
rect 40092 27832 40908 27860
rect 43993 27863 44051 27869
rect 40092 27820 40098 27832
rect 43993 27829 44005 27863
rect 44039 27860 44051 27863
rect 44266 27860 44272 27872
rect 44039 27832 44272 27860
rect 44039 27829 44051 27832
rect 43993 27823 44051 27829
rect 44266 27820 44272 27832
rect 44324 27820 44330 27872
rect 1104 27770 44620 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 44620 27770
rect 1104 27696 44620 27718
rect 4972 27659 5030 27665
rect 4972 27625 4984 27659
rect 5018 27656 5030 27659
rect 5350 27656 5356 27668
rect 5018 27628 5356 27656
rect 5018 27625 5030 27628
rect 4972 27619 5030 27625
rect 5350 27616 5356 27628
rect 5408 27616 5414 27668
rect 6362 27616 6368 27668
rect 6420 27656 6426 27668
rect 6898 27659 6956 27665
rect 6898 27656 6910 27659
rect 6420 27628 6910 27656
rect 6420 27616 6426 27628
rect 6898 27625 6910 27628
rect 6944 27625 6956 27659
rect 6898 27619 6956 27625
rect 8386 27616 8392 27668
rect 8444 27616 8450 27668
rect 10952 27659 11010 27665
rect 10952 27625 10964 27659
rect 10998 27656 11010 27659
rect 11146 27656 11152 27668
rect 10998 27628 11152 27656
rect 10998 27625 11010 27628
rect 10952 27619 11010 27625
rect 11146 27616 11152 27628
rect 11204 27616 11210 27668
rect 12437 27659 12495 27665
rect 12437 27625 12449 27659
rect 12483 27656 12495 27659
rect 12802 27656 12808 27668
rect 12483 27628 12808 27656
rect 12483 27625 12495 27628
rect 12437 27619 12495 27625
rect 12802 27616 12808 27628
rect 12860 27616 12866 27668
rect 12897 27659 12955 27665
rect 12897 27625 12909 27659
rect 12943 27656 12955 27659
rect 13078 27656 13084 27668
rect 12943 27628 13084 27656
rect 12943 27625 12955 27628
rect 12897 27619 12955 27625
rect 13078 27616 13084 27628
rect 13136 27616 13142 27668
rect 13906 27616 13912 27668
rect 13964 27656 13970 27668
rect 13964 27628 14504 27656
rect 13964 27616 13970 27628
rect 14476 27597 14504 27628
rect 15654 27616 15660 27668
rect 15712 27616 15718 27668
rect 16761 27659 16819 27665
rect 16761 27625 16773 27659
rect 16807 27656 16819 27659
rect 17034 27656 17040 27668
rect 16807 27628 17040 27656
rect 16807 27625 16819 27628
rect 16761 27619 16819 27625
rect 17034 27616 17040 27628
rect 17092 27616 17098 27668
rect 17218 27616 17224 27668
rect 17276 27616 17282 27668
rect 19521 27659 19579 27665
rect 19521 27625 19533 27659
rect 19567 27625 19579 27659
rect 19521 27619 19579 27625
rect 14461 27591 14519 27597
rect 14461 27557 14473 27591
rect 14507 27557 14519 27591
rect 15672 27588 15700 27616
rect 15933 27591 15991 27597
rect 15933 27588 15945 27591
rect 15672 27560 15945 27588
rect 14461 27551 14519 27557
rect 15933 27557 15945 27560
rect 15979 27557 15991 27591
rect 16942 27588 16948 27600
rect 15933 27551 15991 27557
rect 16224 27560 16948 27588
rect 4709 27523 4767 27529
rect 4709 27489 4721 27523
rect 4755 27520 4767 27523
rect 6914 27520 6920 27532
rect 4755 27492 6920 27520
rect 4755 27489 4767 27492
rect 4709 27483 4767 27489
rect 6914 27480 6920 27492
rect 6972 27480 6978 27532
rect 12618 27480 12624 27532
rect 12676 27520 12682 27532
rect 13541 27523 13599 27529
rect 12676 27492 13216 27520
rect 12676 27480 12682 27492
rect 934 27412 940 27464
rect 992 27452 998 27464
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 992 27424 1409 27452
rect 992 27412 998 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 6638 27412 6644 27464
rect 6696 27412 6702 27464
rect 9306 27412 9312 27464
rect 9364 27452 9370 27464
rect 9674 27452 9680 27464
rect 9364 27424 9680 27452
rect 9364 27412 9370 27424
rect 9674 27412 9680 27424
rect 9732 27452 9738 27464
rect 10689 27455 10747 27461
rect 10689 27452 10701 27455
rect 9732 27424 10701 27452
rect 9732 27412 9738 27424
rect 10689 27421 10701 27424
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 13078 27412 13084 27464
rect 13136 27412 13142 27464
rect 13188 27461 13216 27492
rect 13541 27489 13553 27523
rect 13587 27520 13599 27523
rect 13587 27492 14688 27520
rect 13587 27489 13599 27492
rect 13541 27483 13599 27489
rect 14660 27464 14688 27492
rect 15102 27480 15108 27532
rect 15160 27480 15166 27532
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 13495 27424 14504 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 7374 27384 7380 27396
rect 6210 27356 7380 27384
rect 7374 27344 7380 27356
rect 7432 27344 7438 27396
rect 8202 27384 8208 27396
rect 8142 27356 8208 27384
rect 8202 27344 8208 27356
rect 8260 27384 8266 27396
rect 9582 27384 9588 27396
rect 8260 27356 9588 27384
rect 8260 27344 8266 27356
rect 9582 27344 9588 27356
rect 9640 27344 9646 27396
rect 12434 27384 12440 27396
rect 12190 27356 12440 27384
rect 12434 27344 12440 27356
rect 12492 27344 12498 27396
rect 1578 27276 1584 27328
rect 1636 27276 1642 27328
rect 6457 27319 6515 27325
rect 6457 27285 6469 27319
rect 6503 27316 6515 27319
rect 7098 27316 7104 27328
rect 6503 27288 7104 27316
rect 6503 27285 6515 27288
rect 6457 27279 6515 27285
rect 7098 27276 7104 27288
rect 7156 27316 7162 27328
rect 13464 27316 13492 27415
rect 14476 27384 14504 27424
rect 14642 27412 14648 27464
rect 14700 27412 14706 27464
rect 14829 27455 14887 27461
rect 14829 27421 14841 27455
rect 14875 27452 14887 27455
rect 15838 27452 15844 27464
rect 14875 27424 15844 27452
rect 14875 27421 14887 27424
rect 14829 27415 14887 27421
rect 15838 27412 15844 27424
rect 15896 27412 15902 27464
rect 15930 27412 15936 27464
rect 15988 27412 15994 27464
rect 16224 27461 16252 27560
rect 16942 27548 16948 27560
rect 17000 27548 17006 27600
rect 17236 27520 17264 27616
rect 18877 27591 18935 27597
rect 18877 27557 18889 27591
rect 18923 27588 18935 27591
rect 19150 27588 19156 27600
rect 18923 27560 19156 27588
rect 18923 27557 18935 27560
rect 18877 27551 18935 27557
rect 19150 27548 19156 27560
rect 19208 27588 19214 27600
rect 19536 27588 19564 27619
rect 19702 27616 19708 27668
rect 19760 27616 19766 27668
rect 19889 27659 19947 27665
rect 19889 27625 19901 27659
rect 19935 27625 19947 27659
rect 19889 27619 19947 27625
rect 19208 27560 19840 27588
rect 19208 27548 19214 27560
rect 16868 27492 17264 27520
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 16577 27455 16635 27461
rect 16577 27421 16589 27455
rect 16623 27452 16635 27455
rect 16666 27452 16672 27464
rect 16623 27424 16672 27452
rect 16623 27421 16635 27424
rect 16577 27415 16635 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 16868 27461 16896 27492
rect 18046 27480 18052 27532
rect 18104 27520 18110 27532
rect 18104 27492 19288 27520
rect 18104 27480 18110 27492
rect 19260 27461 19288 27492
rect 19812 27461 19840 27560
rect 16853 27455 16911 27461
rect 16853 27421 16865 27455
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 17129 27455 17187 27461
rect 17129 27421 17141 27455
rect 17175 27421 17187 27455
rect 17129 27415 17187 27421
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 15948 27384 15976 27412
rect 17144 27384 17172 27415
rect 14476 27356 15976 27384
rect 16592 27356 17172 27384
rect 17405 27387 17463 27393
rect 16592 27328 16620 27356
rect 17405 27353 17417 27387
rect 17451 27353 17463 27387
rect 17405 27347 17463 27353
rect 7156 27288 13492 27316
rect 7156 27276 7162 27288
rect 14918 27276 14924 27328
rect 14976 27276 14982 27328
rect 16574 27276 16580 27328
rect 16632 27276 16638 27328
rect 17037 27319 17095 27325
rect 17037 27285 17049 27319
rect 17083 27316 17095 27319
rect 17420 27316 17448 27347
rect 18046 27344 18052 27396
rect 18104 27344 18110 27396
rect 19150 27344 19156 27396
rect 19208 27384 19214 27396
rect 19260 27384 19288 27415
rect 19904 27384 19932 27619
rect 20070 27616 20076 27668
rect 20128 27656 20134 27668
rect 20257 27659 20315 27665
rect 20257 27656 20269 27659
rect 20128 27628 20269 27656
rect 20128 27616 20134 27628
rect 20257 27625 20269 27628
rect 20303 27625 20315 27659
rect 20257 27619 20315 27625
rect 22554 27616 22560 27668
rect 22612 27656 22618 27668
rect 23385 27659 23443 27665
rect 23385 27656 23397 27659
rect 22612 27628 23397 27656
rect 22612 27616 22618 27628
rect 23385 27625 23397 27628
rect 23431 27625 23443 27659
rect 23385 27619 23443 27625
rect 24213 27659 24271 27665
rect 24213 27625 24225 27659
rect 24259 27656 24271 27659
rect 24394 27656 24400 27668
rect 24259 27628 24400 27656
rect 24259 27625 24271 27628
rect 24213 27619 24271 27625
rect 24394 27616 24400 27628
rect 24452 27616 24458 27668
rect 24578 27616 24584 27668
rect 24636 27656 24642 27668
rect 25298 27659 25356 27665
rect 25298 27656 25310 27659
rect 24636 27628 25310 27656
rect 24636 27616 24642 27628
rect 25298 27625 25310 27628
rect 25344 27625 25356 27659
rect 25298 27619 25356 27625
rect 33321 27659 33379 27665
rect 33321 27625 33333 27659
rect 33367 27656 33379 27659
rect 33594 27656 33600 27668
rect 33367 27628 33600 27656
rect 33367 27625 33379 27628
rect 33321 27619 33379 27625
rect 33594 27616 33600 27628
rect 33652 27616 33658 27668
rect 35710 27616 35716 27668
rect 35768 27656 35774 27668
rect 37642 27656 37648 27668
rect 35768 27628 37648 27656
rect 35768 27616 35774 27628
rect 37642 27616 37648 27628
rect 37700 27656 37706 27668
rect 39574 27656 39580 27668
rect 37700 27628 39580 27656
rect 37700 27616 37706 27628
rect 39574 27616 39580 27628
rect 39632 27616 39638 27668
rect 23106 27548 23112 27600
rect 23164 27548 23170 27600
rect 23860 27560 25181 27588
rect 21634 27412 21640 27464
rect 21692 27412 21698 27464
rect 23124 27452 23152 27548
rect 23474 27480 23480 27532
rect 23532 27520 23538 27532
rect 23569 27523 23627 27529
rect 23569 27520 23581 27523
rect 23532 27492 23581 27520
rect 23532 27480 23538 27492
rect 23569 27489 23581 27492
rect 23615 27489 23627 27523
rect 23569 27483 23627 27489
rect 23860 27461 23888 27560
rect 24670 27480 24676 27532
rect 24728 27520 24734 27532
rect 25041 27523 25099 27529
rect 25041 27520 25053 27523
rect 24728 27492 25053 27520
rect 24728 27480 24734 27492
rect 25041 27489 25053 27492
rect 25087 27489 25099 27523
rect 25153 27520 25181 27560
rect 36170 27548 36176 27600
rect 36228 27588 36234 27600
rect 37734 27588 37740 27600
rect 36228 27560 37740 27588
rect 36228 27548 36234 27560
rect 37734 27548 37740 27560
rect 37792 27548 37798 27600
rect 38378 27548 38384 27600
rect 38436 27548 38442 27600
rect 39301 27591 39359 27597
rect 39301 27557 39313 27591
rect 39347 27588 39359 27591
rect 39850 27588 39856 27600
rect 39347 27560 39856 27588
rect 39347 27557 39359 27560
rect 39301 27551 39359 27557
rect 39850 27548 39856 27560
rect 39908 27548 39914 27600
rect 40957 27591 41015 27597
rect 40957 27557 40969 27591
rect 41003 27588 41015 27591
rect 41690 27588 41696 27600
rect 41003 27560 41696 27588
rect 41003 27557 41015 27560
rect 40957 27551 41015 27557
rect 41690 27548 41696 27560
rect 41748 27548 41754 27600
rect 43165 27591 43223 27597
rect 42628 27560 42932 27588
rect 26326 27520 26332 27532
rect 25153 27492 26332 27520
rect 25041 27483 25099 27489
rect 26326 27480 26332 27492
rect 26384 27520 26390 27532
rect 26789 27523 26847 27529
rect 26789 27520 26801 27523
rect 26384 27492 26801 27520
rect 26384 27480 26390 27492
rect 26789 27489 26801 27492
rect 26835 27489 26847 27523
rect 26789 27483 26847 27489
rect 34057 27523 34115 27529
rect 34057 27489 34069 27523
rect 34103 27520 34115 27523
rect 34330 27520 34336 27532
rect 34103 27492 34336 27520
rect 34103 27489 34115 27492
rect 34057 27483 34115 27489
rect 34330 27480 34336 27492
rect 34388 27480 34394 27532
rect 35802 27480 35808 27532
rect 35860 27520 35866 27532
rect 35860 27492 36952 27520
rect 35860 27480 35866 27492
rect 23046 27424 23152 27452
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 24394 27412 24400 27464
rect 24452 27412 24458 27464
rect 24946 27412 24952 27464
rect 25004 27412 25010 27464
rect 28350 27412 28356 27464
rect 28408 27412 28414 27464
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 32674 27412 32680 27464
rect 32732 27452 32738 27464
rect 32769 27455 32827 27461
rect 32769 27452 32781 27455
rect 32732 27424 32781 27452
rect 32732 27412 32738 27424
rect 32769 27421 32781 27424
rect 32815 27421 32827 27455
rect 32769 27415 32827 27421
rect 33137 27455 33195 27461
rect 33137 27421 33149 27455
rect 33183 27452 33195 27455
rect 33226 27452 33232 27464
rect 33183 27424 33232 27452
rect 33183 27421 33195 27424
rect 33137 27415 33195 27421
rect 33226 27412 33232 27424
rect 33284 27452 33290 27464
rect 33778 27452 33784 27464
rect 33284 27424 33784 27452
rect 33284 27412 33290 27424
rect 33778 27412 33784 27424
rect 33836 27412 33842 27464
rect 36924 27461 36952 27492
rect 37458 27480 37464 27532
rect 37516 27520 37522 27532
rect 38396 27520 38424 27548
rect 37516 27492 40908 27520
rect 37516 27480 37522 27492
rect 34885 27455 34943 27461
rect 34885 27421 34897 27455
rect 34931 27421 34943 27455
rect 36909 27455 36967 27461
rect 34885 27415 34943 27421
rect 19208 27356 19932 27384
rect 19208 27344 19214 27356
rect 21910 27344 21916 27396
rect 21968 27344 21974 27396
rect 17083 27288 17448 27316
rect 17083 27285 17095 27288
rect 17037 27279 17095 27285
rect 23750 27276 23756 27328
rect 23808 27276 23814 27328
rect 24581 27319 24639 27325
rect 24581 27285 24593 27319
rect 24627 27316 24639 27319
rect 24964 27316 24992 27412
rect 25314 27344 25320 27396
rect 25372 27384 25378 27396
rect 29362 27384 29368 27396
rect 25372 27356 25806 27384
rect 28828 27356 29368 27384
rect 25372 27344 25378 27356
rect 24627 27288 24992 27316
rect 25700 27316 25728 27356
rect 28828 27316 28856 27356
rect 29362 27344 29368 27356
rect 29420 27384 29426 27396
rect 30006 27384 30012 27396
rect 29420 27356 30012 27384
rect 29420 27344 29426 27356
rect 30006 27344 30012 27356
rect 30064 27384 30070 27396
rect 32582 27384 32588 27396
rect 30064 27356 32588 27384
rect 30064 27344 30070 27356
rect 32582 27344 32588 27356
rect 32640 27344 32646 27396
rect 32953 27387 33011 27393
rect 32953 27353 32965 27387
rect 32999 27353 33011 27387
rect 32953 27347 33011 27353
rect 33045 27387 33103 27393
rect 33045 27353 33057 27387
rect 33091 27384 33103 27387
rect 33413 27387 33471 27393
rect 33413 27384 33425 27387
rect 33091 27356 33425 27384
rect 33091 27353 33103 27356
rect 33045 27347 33103 27353
rect 33413 27353 33425 27356
rect 33459 27353 33471 27387
rect 33413 27347 33471 27353
rect 25700 27288 28856 27316
rect 28905 27319 28963 27325
rect 24627 27285 24639 27288
rect 24581 27279 24639 27285
rect 28905 27285 28917 27319
rect 28951 27316 28963 27319
rect 29454 27316 29460 27328
rect 28951 27288 29460 27316
rect 28951 27285 28963 27288
rect 28905 27279 28963 27285
rect 29454 27276 29460 27288
rect 29512 27276 29518 27328
rect 31938 27276 31944 27328
rect 31996 27276 32002 27328
rect 32398 27276 32404 27328
rect 32456 27316 32462 27328
rect 32858 27316 32864 27328
rect 32456 27288 32864 27316
rect 32456 27276 32462 27288
rect 32858 27276 32864 27288
rect 32916 27316 32922 27328
rect 32968 27316 32996 27347
rect 32916 27288 32996 27316
rect 32916 27276 32922 27288
rect 33870 27276 33876 27328
rect 33928 27316 33934 27328
rect 34900 27316 34928 27415
rect 35158 27344 35164 27396
rect 35216 27344 35222 27396
rect 35342 27316 35348 27328
rect 33928 27288 35348 27316
rect 33928 27276 33934 27288
rect 35342 27276 35348 27288
rect 35400 27276 35406 27328
rect 35986 27276 35992 27328
rect 36044 27316 36050 27328
rect 36280 27316 36308 27438
rect 36909 27421 36921 27455
rect 36955 27452 36967 27455
rect 38654 27452 38660 27464
rect 36955 27424 38660 27452
rect 36955 27421 36967 27424
rect 36909 27415 36967 27421
rect 38654 27412 38660 27424
rect 38712 27412 38718 27464
rect 38749 27455 38807 27461
rect 38749 27421 38761 27455
rect 38795 27452 38807 27455
rect 38838 27452 38844 27464
rect 38795 27424 38844 27452
rect 38795 27421 38807 27424
rect 38749 27415 38807 27421
rect 38838 27412 38844 27424
rect 38896 27412 38902 27464
rect 39114 27412 39120 27464
rect 39172 27412 39178 27464
rect 40497 27455 40555 27461
rect 40497 27421 40509 27455
rect 40543 27452 40555 27455
rect 40770 27452 40776 27464
rect 40543 27424 40776 27452
rect 40543 27421 40555 27424
rect 40497 27415 40555 27421
rect 37734 27344 37740 27396
rect 37792 27384 37798 27396
rect 38470 27384 38476 27396
rect 37792 27356 38476 27384
rect 37792 27344 37798 27356
rect 38470 27344 38476 27356
rect 38528 27384 38534 27396
rect 38933 27387 38991 27393
rect 38933 27384 38945 27387
rect 38528 27356 38945 27384
rect 38528 27344 38534 27356
rect 38933 27353 38945 27356
rect 38979 27353 38991 27387
rect 38933 27347 38991 27353
rect 39025 27387 39083 27393
rect 39025 27353 39037 27387
rect 39071 27384 39083 27387
rect 39206 27384 39212 27396
rect 39071 27356 39212 27384
rect 39071 27353 39083 27356
rect 39025 27347 39083 27353
rect 39206 27344 39212 27356
rect 39264 27384 39270 27396
rect 40512 27384 40540 27415
rect 40770 27412 40776 27424
rect 40828 27412 40834 27464
rect 40880 27452 40908 27492
rect 41046 27480 41052 27532
rect 41104 27520 41110 27532
rect 42628 27529 42656 27560
rect 41417 27523 41475 27529
rect 41104 27492 41276 27520
rect 41104 27480 41110 27492
rect 41248 27461 41276 27492
rect 41417 27489 41429 27523
rect 41463 27489 41475 27523
rect 41417 27483 41475 27489
rect 42613 27523 42671 27529
rect 42613 27489 42625 27523
rect 42659 27489 42671 27523
rect 42613 27483 42671 27489
rect 42705 27523 42763 27529
rect 42705 27489 42717 27523
rect 42751 27520 42763 27523
rect 42794 27520 42800 27532
rect 42751 27492 42800 27520
rect 42751 27489 42763 27492
rect 42705 27483 42763 27489
rect 41141 27455 41199 27461
rect 41141 27452 41153 27455
rect 40880 27424 41153 27452
rect 41141 27421 41153 27424
rect 41187 27421 41199 27455
rect 41141 27415 41199 27421
rect 41233 27455 41291 27461
rect 41233 27421 41245 27455
rect 41279 27421 41291 27455
rect 41233 27415 41291 27421
rect 39264 27356 40540 27384
rect 39264 27344 39270 27356
rect 36044 27288 36308 27316
rect 36633 27319 36691 27325
rect 36044 27276 36050 27288
rect 36633 27285 36645 27319
rect 36679 27316 36691 27319
rect 36722 27316 36728 27328
rect 36679 27288 36728 27316
rect 36679 27285 36691 27288
rect 36633 27279 36691 27285
rect 36722 27276 36728 27288
rect 36780 27276 36786 27328
rect 38102 27276 38108 27328
rect 38160 27316 38166 27328
rect 38197 27319 38255 27325
rect 38197 27316 38209 27319
rect 38160 27288 38209 27316
rect 38160 27276 38166 27288
rect 38197 27285 38209 27288
rect 38243 27285 38255 27319
rect 38197 27279 38255 27285
rect 39850 27276 39856 27328
rect 39908 27276 39914 27328
rect 41156 27316 41184 27415
rect 41322 27344 41328 27396
rect 41380 27384 41386 27396
rect 41432 27384 41460 27483
rect 41509 27455 41567 27461
rect 41509 27421 41521 27455
rect 41555 27452 41567 27455
rect 42720 27452 42748 27483
rect 42794 27480 42800 27492
rect 42852 27480 42858 27532
rect 41555 27424 42748 27452
rect 42904 27452 42932 27560
rect 43165 27557 43177 27591
rect 43211 27557 43223 27591
rect 43165 27551 43223 27557
rect 43180 27520 43208 27551
rect 43180 27492 44220 27520
rect 43162 27452 43168 27464
rect 42904 27424 43168 27452
rect 41555 27421 41567 27424
rect 41509 27415 41567 27421
rect 43162 27412 43168 27424
rect 43220 27412 43226 27464
rect 43806 27412 43812 27464
rect 43864 27412 43870 27464
rect 44192 27461 44220 27492
rect 44177 27455 44235 27461
rect 44177 27421 44189 27455
rect 44223 27421 44235 27455
rect 44177 27415 44235 27421
rect 41380 27356 41460 27384
rect 41380 27344 41386 27356
rect 41230 27316 41236 27328
rect 41156 27288 41236 27316
rect 41230 27276 41236 27288
rect 41288 27276 41294 27328
rect 42794 27276 42800 27328
rect 42852 27276 42858 27328
rect 42886 27276 42892 27328
rect 42944 27316 42950 27328
rect 43257 27319 43315 27325
rect 43257 27316 43269 27319
rect 42944 27288 43269 27316
rect 42944 27276 42950 27288
rect 43257 27285 43269 27288
rect 43303 27285 43315 27319
rect 43257 27279 43315 27285
rect 43990 27276 43996 27328
rect 44048 27276 44054 27328
rect 1104 27226 44620 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 44620 27226
rect 1104 27152 44620 27174
rect 10318 27072 10324 27124
rect 10376 27112 10382 27124
rect 14918 27112 14924 27124
rect 10376 27084 14924 27112
rect 10376 27072 10382 27084
rect 14918 27072 14924 27084
rect 14976 27072 14982 27124
rect 16758 27072 16764 27124
rect 16816 27072 16822 27124
rect 17126 27112 17132 27124
rect 16960 27084 17132 27112
rect 8478 27004 8484 27056
rect 8536 27044 8542 27056
rect 8849 27047 8907 27053
rect 8849 27044 8861 27047
rect 8536 27016 8861 27044
rect 8536 27004 8542 27016
rect 8849 27013 8861 27016
rect 8895 27013 8907 27047
rect 12434 27044 12440 27056
rect 10074 27030 12440 27044
rect 8849 27007 8907 27013
rect 10060 27016 12440 27030
rect 6638 26868 6644 26920
rect 6696 26908 6702 26920
rect 8570 26908 8576 26920
rect 6696 26880 8576 26908
rect 6696 26868 6702 26880
rect 8570 26868 8576 26880
rect 8628 26868 8634 26920
rect 9582 26868 9588 26920
rect 9640 26908 9646 26920
rect 10060 26908 10088 27016
rect 12434 27004 12440 27016
rect 12492 27004 12498 27056
rect 16776 27044 16804 27072
rect 16960 27053 16988 27084
rect 17126 27072 17132 27084
rect 17184 27072 17190 27124
rect 18417 27115 18475 27121
rect 18417 27081 18429 27115
rect 18463 27112 18475 27115
rect 18506 27112 18512 27124
rect 18463 27084 18512 27112
rect 18463 27081 18475 27084
rect 18417 27075 18475 27081
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 21910 27072 21916 27124
rect 21968 27112 21974 27124
rect 22005 27115 22063 27121
rect 22005 27112 22017 27115
rect 21968 27084 22017 27112
rect 21968 27072 21974 27084
rect 22005 27081 22017 27084
rect 22051 27081 22063 27115
rect 22005 27075 22063 27081
rect 22094 27072 22100 27124
rect 22152 27072 22158 27124
rect 24394 27072 24400 27124
rect 24452 27112 24458 27124
rect 24765 27115 24823 27121
rect 24765 27112 24777 27115
rect 24452 27084 24777 27112
rect 24452 27072 24458 27084
rect 24765 27081 24777 27084
rect 24811 27081 24823 27115
rect 24765 27075 24823 27081
rect 26234 27072 26240 27124
rect 26292 27072 26298 27124
rect 29638 27072 29644 27124
rect 29696 27112 29702 27124
rect 31849 27115 31907 27121
rect 29696 27084 31524 27112
rect 29696 27072 29702 27084
rect 16500 27016 16804 27044
rect 16945 27047 17003 27053
rect 16500 26985 16528 27016
rect 16945 27013 16957 27047
rect 16991 27013 17003 27047
rect 16945 27007 17003 27013
rect 16485 26979 16543 26985
rect 16485 26945 16497 26979
rect 16531 26945 16543 26979
rect 16485 26939 16543 26945
rect 18046 26936 18052 26988
rect 18104 26936 18110 26988
rect 19426 26936 19432 26988
rect 19484 26976 19490 26988
rect 20441 26979 20499 26985
rect 20441 26976 20453 26979
rect 19484 26948 20453 26976
rect 19484 26936 19490 26948
rect 20441 26945 20453 26948
rect 20487 26976 20499 26979
rect 20622 26976 20628 26988
rect 20487 26948 20628 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 20622 26936 20628 26948
rect 20680 26936 20686 26988
rect 22112 26976 22140 27072
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 22112 26948 22201 26976
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 24397 26979 24455 26985
rect 24397 26945 24409 26979
rect 24443 26976 24455 26979
rect 26252 26976 26280 27072
rect 28445 27047 28503 27053
rect 28445 27013 28457 27047
rect 28491 27044 28503 27047
rect 28813 27047 28871 27053
rect 28813 27044 28825 27047
rect 28491 27016 28825 27044
rect 28491 27013 28503 27016
rect 28445 27007 28503 27013
rect 28813 27013 28825 27016
rect 28859 27013 28871 27047
rect 28813 27007 28871 27013
rect 29319 27047 29377 27053
rect 29319 27013 29331 27047
rect 29365 27044 29377 27047
rect 30190 27044 30196 27056
rect 29365 27016 30196 27044
rect 29365 27013 29377 27016
rect 29319 27007 29377 27013
rect 30190 27004 30196 27016
rect 30248 27004 30254 27056
rect 28997 26979 29055 26985
rect 24443 26948 26280 26976
rect 26896 26948 27370 26976
rect 24443 26945 24455 26948
rect 24397 26939 24455 26945
rect 9640 26880 10088 26908
rect 9640 26868 9646 26880
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 13722 26908 13728 26920
rect 11480 26880 13728 26908
rect 11480 26868 11486 26880
rect 13722 26868 13728 26880
rect 13780 26908 13786 26920
rect 16209 26911 16267 26917
rect 16209 26908 16221 26911
rect 13780 26880 16221 26908
rect 13780 26868 13786 26880
rect 16209 26877 16221 26880
rect 16255 26877 16267 26911
rect 16209 26871 16267 26877
rect 16574 26868 16580 26920
rect 16632 26908 16638 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 16632 26880 16681 26908
rect 16632 26868 16638 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 18064 26908 18092 26936
rect 16669 26871 16727 26877
rect 16776 26880 18092 26908
rect 15654 26800 15660 26852
rect 15712 26840 15718 26852
rect 16776 26840 16804 26880
rect 18322 26868 18328 26920
rect 18380 26908 18386 26920
rect 20165 26911 20223 26917
rect 20165 26908 20177 26911
rect 18380 26880 20177 26908
rect 18380 26868 18386 26880
rect 20165 26877 20177 26880
rect 20211 26877 20223 26911
rect 20165 26871 20223 26877
rect 20254 26868 20260 26920
rect 20312 26908 20318 26920
rect 20349 26911 20407 26917
rect 20349 26908 20361 26911
rect 20312 26880 20361 26908
rect 20312 26868 20318 26880
rect 20349 26877 20361 26880
rect 20395 26877 20407 26911
rect 20349 26871 20407 26877
rect 23474 26868 23480 26920
rect 23532 26908 23538 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 23532 26880 24133 26908
rect 23532 26868 23538 26880
rect 24121 26877 24133 26880
rect 24167 26877 24179 26911
rect 24121 26871 24179 26877
rect 24302 26868 24308 26920
rect 24360 26868 24366 26920
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 26896 26908 26924 26948
rect 28997 26945 29009 26979
rect 29043 26945 29055 26979
rect 28997 26939 29055 26945
rect 25372 26880 26924 26908
rect 26973 26911 27031 26917
rect 25372 26868 25378 26880
rect 26973 26877 26985 26911
rect 27019 26908 27031 26911
rect 28350 26908 28356 26920
rect 27019 26880 28356 26908
rect 27019 26877 27031 26880
rect 26973 26871 27031 26877
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 28718 26868 28724 26920
rect 28776 26868 28782 26920
rect 29012 26908 29040 26939
rect 29086 26936 29092 26988
rect 29144 26936 29150 26988
rect 29178 26936 29184 26988
rect 29236 26936 29242 26988
rect 29454 26936 29460 26988
rect 29512 26936 29518 26988
rect 29546 26936 29552 26988
rect 29604 26936 29610 26988
rect 29730 26936 29736 26988
rect 29788 26936 29794 26988
rect 31496 26985 31524 27084
rect 31849 27081 31861 27115
rect 31895 27112 31907 27115
rect 32030 27112 32036 27124
rect 31895 27084 32036 27112
rect 31895 27081 31907 27084
rect 31849 27075 31907 27081
rect 32030 27072 32036 27084
rect 32088 27072 32094 27124
rect 32306 27072 32312 27124
rect 32364 27072 32370 27124
rect 34514 27072 34520 27124
rect 34572 27072 34578 27124
rect 35158 27072 35164 27124
rect 35216 27112 35222 27124
rect 35621 27115 35679 27121
rect 35621 27112 35633 27115
rect 35216 27084 35633 27112
rect 35216 27072 35222 27084
rect 35621 27081 35633 27084
rect 35667 27081 35679 27115
rect 37458 27112 37464 27124
rect 35621 27075 35679 27081
rect 36648 27084 37464 27112
rect 31665 27047 31723 27053
rect 31665 27013 31677 27047
rect 31711 27044 31723 27047
rect 34532 27044 34560 27072
rect 31711 27016 32352 27044
rect 31711 27013 31723 27016
rect 31665 27007 31723 27013
rect 32324 26985 32352 27016
rect 34256 27016 34744 27044
rect 34256 26988 34284 27016
rect 31481 26979 31539 26985
rect 31481 26945 31493 26979
rect 31527 26976 31539 26979
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 31527 26948 32137 26976
rect 31527 26945 31539 26948
rect 31481 26939 31539 26945
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26976 32367 26979
rect 32858 26976 32864 26988
rect 32355 26948 32864 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 32858 26936 32864 26948
rect 32916 26936 32922 26988
rect 34238 26936 34244 26988
rect 34296 26936 34302 26988
rect 34333 26979 34391 26985
rect 34333 26945 34345 26979
rect 34379 26945 34391 26979
rect 34333 26939 34391 26945
rect 34517 26979 34575 26985
rect 34517 26945 34529 26979
rect 34563 26945 34575 26979
rect 34517 26939 34575 26945
rect 29641 26911 29699 26917
rect 29641 26908 29653 26911
rect 29012 26880 29653 26908
rect 29641 26877 29653 26880
rect 29687 26877 29699 26911
rect 34348 26908 34376 26939
rect 34422 26908 34428 26920
rect 34348 26880 34428 26908
rect 29641 26871 29699 26877
rect 34422 26868 34428 26880
rect 34480 26868 34486 26920
rect 15712 26812 16804 26840
rect 15712 26800 15718 26812
rect 17954 26800 17960 26852
rect 18012 26840 18018 26852
rect 18414 26840 18420 26852
rect 18012 26812 18420 26840
rect 18012 26800 18018 26812
rect 18414 26800 18420 26812
rect 18472 26800 18478 26852
rect 25406 26800 25412 26852
rect 25464 26800 25470 26852
rect 28736 26840 28764 26868
rect 31294 26840 31300 26852
rect 28736 26812 31300 26840
rect 31294 26800 31300 26812
rect 31352 26840 31358 26852
rect 31938 26840 31944 26852
rect 31352 26812 31944 26840
rect 31352 26800 31358 26812
rect 31938 26800 31944 26812
rect 31996 26800 32002 26852
rect 34054 26800 34060 26852
rect 34112 26840 34118 26852
rect 34532 26840 34560 26939
rect 34606 26936 34612 26988
rect 34664 26936 34670 26988
rect 34716 26985 34744 27016
rect 36648 26985 36676 27084
rect 37458 27072 37464 27084
rect 37516 27072 37522 27124
rect 37550 27072 37556 27124
rect 37608 27112 37614 27124
rect 37921 27115 37979 27121
rect 37921 27112 37933 27115
rect 37608 27084 37933 27112
rect 37608 27072 37614 27084
rect 37921 27081 37933 27084
rect 37967 27081 37979 27115
rect 37921 27075 37979 27081
rect 38120 27084 38332 27112
rect 37016 27016 37688 27044
rect 34701 26979 34759 26985
rect 34701 26945 34713 26979
rect 34747 26945 34759 26979
rect 36633 26979 36691 26985
rect 34701 26939 34759 26945
rect 34900 26948 35388 26976
rect 34624 26908 34652 26936
rect 34900 26908 34928 26948
rect 34624 26880 34928 26908
rect 34977 26911 35035 26917
rect 34977 26877 34989 26911
rect 35023 26877 35035 26911
rect 35360 26908 35388 26948
rect 36633 26945 36645 26979
rect 36679 26945 36691 26979
rect 36633 26939 36691 26945
rect 36722 26936 36728 26988
rect 36780 26936 36786 26988
rect 37016 26985 37044 27016
rect 37660 26988 37688 27016
rect 37734 27004 37740 27056
rect 37792 27044 37798 27056
rect 38120 27044 38148 27084
rect 37792 27016 38148 27044
rect 37792 27004 37798 27016
rect 38194 27004 38200 27056
rect 38252 27004 38258 27056
rect 38304 27053 38332 27084
rect 38654 27072 38660 27124
rect 38712 27112 38718 27124
rect 42518 27112 42524 27124
rect 38712 27084 42524 27112
rect 38712 27072 38718 27084
rect 42518 27072 42524 27084
rect 42576 27072 42582 27124
rect 38289 27047 38347 27053
rect 38289 27013 38301 27047
rect 38335 27013 38347 27047
rect 39114 27044 39120 27056
rect 38289 27007 38347 27013
rect 38396 27016 39120 27044
rect 37001 26979 37059 26985
rect 37001 26945 37013 26979
rect 37047 26945 37059 26979
rect 37001 26939 37059 26945
rect 37277 26979 37335 26985
rect 37277 26945 37289 26979
rect 37323 26976 37335 26979
rect 37366 26976 37372 26988
rect 37323 26948 37372 26976
rect 37323 26945 37335 26948
rect 37277 26939 37335 26945
rect 37366 26936 37372 26948
rect 37424 26936 37430 26988
rect 37458 26936 37464 26988
rect 37516 26936 37522 26988
rect 37553 26979 37611 26985
rect 37553 26945 37565 26979
rect 37599 26945 37611 26979
rect 37553 26939 37611 26945
rect 36740 26908 36768 26936
rect 35360 26880 36768 26908
rect 37568 26908 37596 26939
rect 37642 26936 37648 26988
rect 37700 26936 37706 26988
rect 37826 26936 37832 26988
rect 37884 26936 37890 26988
rect 37918 26936 37924 26988
rect 37976 26936 37982 26988
rect 38105 26979 38163 26985
rect 38105 26945 38117 26979
rect 38151 26976 38163 26979
rect 38396 26976 38424 27016
rect 39114 27004 39120 27016
rect 39172 27004 39178 27056
rect 39850 27004 39856 27056
rect 39908 27004 39914 27056
rect 39942 27004 39948 27056
rect 40000 27044 40006 27056
rect 40000 27016 41184 27044
rect 40000 27004 40006 27016
rect 38151 26948 38424 26976
rect 38473 26979 38531 26985
rect 38151 26945 38163 26948
rect 38105 26939 38163 26945
rect 38473 26945 38485 26979
rect 38519 26976 38531 26979
rect 39868 26976 39896 27004
rect 41156 26985 41184 27016
rect 43254 27004 43260 27056
rect 43312 27004 43318 27056
rect 38519 26948 39896 26976
rect 40865 26979 40923 26985
rect 38519 26945 38531 26948
rect 38473 26939 38531 26945
rect 40865 26945 40877 26979
rect 40911 26945 40923 26979
rect 40865 26939 40923 26945
rect 41141 26979 41199 26985
rect 41141 26945 41153 26979
rect 41187 26945 41199 26979
rect 41141 26939 41199 26945
rect 37936 26908 37964 26936
rect 37568 26880 37964 26908
rect 34977 26871 35035 26877
rect 34112 26812 34560 26840
rect 34112 26800 34118 26812
rect 14642 26732 14648 26784
rect 14700 26772 14706 26784
rect 17972 26772 18000 26800
rect 14700 26744 18000 26772
rect 20809 26775 20867 26781
rect 14700 26732 14706 26744
rect 20809 26741 20821 26775
rect 20855 26772 20867 26775
rect 21266 26772 21272 26784
rect 20855 26744 21272 26772
rect 20855 26741 20867 26744
rect 20809 26735 20867 26741
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 25424 26772 25452 26800
rect 29270 26772 29276 26784
rect 25424 26744 29276 26772
rect 29270 26732 29276 26744
rect 29328 26732 29334 26784
rect 34532 26772 34560 26812
rect 34885 26843 34943 26849
rect 34885 26809 34897 26843
rect 34931 26840 34943 26843
rect 34992 26840 35020 26871
rect 34931 26812 35020 26840
rect 34931 26809 34943 26812
rect 34885 26803 34943 26809
rect 35894 26800 35900 26852
rect 35952 26840 35958 26852
rect 38120 26840 38148 26939
rect 40678 26868 40684 26920
rect 40736 26868 40742 26920
rect 40880 26840 40908 26939
rect 41230 26936 41236 26988
rect 41288 26936 41294 26988
rect 44266 26936 44272 26988
rect 44324 26936 44330 26988
rect 40954 26868 40960 26920
rect 41012 26908 41018 26920
rect 41322 26908 41328 26920
rect 41012 26880 41328 26908
rect 41012 26868 41018 26880
rect 41322 26868 41328 26880
rect 41380 26868 41386 26920
rect 41417 26911 41475 26917
rect 41417 26877 41429 26911
rect 41463 26908 41475 26911
rect 41509 26911 41567 26917
rect 41509 26908 41521 26911
rect 41463 26880 41521 26908
rect 41463 26877 41475 26880
rect 41417 26871 41475 26877
rect 41509 26877 41521 26880
rect 41555 26877 41567 26911
rect 41509 26871 41567 26877
rect 42521 26911 42579 26917
rect 42521 26877 42533 26911
rect 42567 26908 42579 26911
rect 42794 26908 42800 26920
rect 42567 26880 42800 26908
rect 42567 26877 42579 26880
rect 42521 26871 42579 26877
rect 42794 26868 42800 26880
rect 42852 26868 42858 26920
rect 43990 26868 43996 26920
rect 44048 26868 44054 26920
rect 42886 26840 42892 26852
rect 35952 26812 38148 26840
rect 40052 26812 40264 26840
rect 40880 26812 42892 26840
rect 35952 26800 35958 26812
rect 36170 26772 36176 26784
rect 34532 26744 36176 26772
rect 36170 26732 36176 26744
rect 36228 26732 36234 26784
rect 36446 26732 36452 26784
rect 36504 26732 36510 26784
rect 36909 26775 36967 26781
rect 36909 26741 36921 26775
rect 36955 26772 36967 26775
rect 37737 26775 37795 26781
rect 37737 26772 37749 26775
rect 36955 26744 37749 26772
rect 36955 26741 36967 26744
rect 36909 26735 36967 26741
rect 37737 26741 37749 26744
rect 37783 26772 37795 26775
rect 40052 26772 40080 26812
rect 37783 26744 40080 26772
rect 37783 26741 37795 26744
rect 37737 26735 37795 26741
rect 40126 26732 40132 26784
rect 40184 26732 40190 26784
rect 40236 26772 40264 26812
rect 42886 26800 42892 26812
rect 42944 26800 42950 26852
rect 40954 26772 40960 26784
rect 40236 26744 40960 26772
rect 40954 26732 40960 26744
rect 41012 26732 41018 26784
rect 42150 26732 42156 26784
rect 42208 26732 42214 26784
rect 1104 26682 44620 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 44620 26682
rect 1104 26608 44620 26630
rect 1578 26528 1584 26580
rect 1636 26568 1642 26580
rect 1636 26540 2774 26568
rect 1636 26528 1642 26540
rect 2746 26500 2774 26540
rect 8570 26528 8576 26580
rect 8628 26568 8634 26580
rect 9674 26568 9680 26580
rect 8628 26540 9680 26568
rect 8628 26528 8634 26540
rect 9674 26528 9680 26540
rect 9732 26528 9738 26580
rect 13262 26568 13268 26580
rect 11164 26540 13268 26568
rect 4985 26503 5043 26509
rect 4985 26500 4997 26503
rect 2746 26472 4997 26500
rect 4985 26469 4997 26472
rect 5031 26469 5043 26503
rect 4985 26463 5043 26469
rect 9398 26460 9404 26512
rect 9456 26460 9462 26512
rect 4893 26435 4951 26441
rect 4893 26401 4905 26435
rect 4939 26432 4951 26435
rect 5718 26432 5724 26444
rect 4939 26404 5724 26432
rect 4939 26401 4951 26404
rect 4893 26395 4951 26401
rect 5718 26392 5724 26404
rect 5776 26392 5782 26444
rect 6270 26392 6276 26444
rect 6328 26392 6334 26444
rect 9416 26432 9444 26460
rect 9048 26404 9444 26432
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26364 5411 26367
rect 6288 26364 6316 26392
rect 9048 26376 9076 26404
rect 5399 26336 6316 26364
rect 5399 26333 5411 26336
rect 5353 26327 5411 26333
rect 9030 26324 9036 26376
rect 9088 26324 9094 26376
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26364 9275 26367
rect 9490 26364 9496 26376
rect 9263 26336 9496 26364
rect 9263 26333 9275 26336
rect 9217 26327 9275 26333
rect 9490 26324 9496 26336
rect 9548 26324 9554 26376
rect 11164 26373 11192 26540
rect 13262 26528 13268 26540
rect 13320 26568 13326 26580
rect 13320 26540 18000 26568
rect 13320 26528 13326 26540
rect 12345 26503 12403 26509
rect 12345 26469 12357 26503
rect 12391 26469 12403 26503
rect 12345 26463 12403 26469
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26333 11207 26367
rect 11149 26327 11207 26333
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12360 26364 12388 26463
rect 12526 26460 12532 26512
rect 12584 26500 12590 26512
rect 15102 26500 15108 26512
rect 12584 26472 13032 26500
rect 12584 26460 12590 26472
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 13004 26441 13032 26472
rect 14752 26472 15108 26500
rect 14752 26441 14780 26472
rect 15102 26460 15108 26472
rect 15160 26500 15166 26512
rect 17402 26500 17408 26512
rect 15160 26472 17408 26500
rect 15160 26460 15166 26472
rect 17402 26460 17408 26472
rect 17460 26460 17466 26512
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12676 26404 12817 26432
rect 12676 26392 12682 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 12989 26435 13047 26441
rect 12989 26401 13001 26435
rect 13035 26432 13047 26435
rect 14737 26435 14795 26441
rect 14737 26432 14749 26435
rect 13035 26404 14749 26432
rect 13035 26401 13047 26404
rect 12989 26395 13047 26401
rect 14737 26401 14749 26404
rect 14783 26401 14795 26435
rect 14737 26395 14795 26401
rect 15838 26392 15844 26444
rect 15896 26432 15902 26444
rect 16390 26432 16396 26444
rect 15896 26404 16396 26432
rect 15896 26392 15902 26404
rect 16390 26392 16396 26404
rect 16448 26392 16454 26444
rect 12299 26336 12388 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 9125 26299 9183 26305
rect 9125 26265 9137 26299
rect 9171 26296 9183 26299
rect 9766 26296 9772 26308
rect 9171 26268 9772 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 10594 26256 10600 26308
rect 10652 26296 10658 26308
rect 12636 26296 12664 26392
rect 13817 26367 13875 26373
rect 13817 26333 13829 26367
rect 13863 26364 13875 26367
rect 13906 26364 13912 26376
rect 13863 26336 13912 26364
rect 13863 26333 13875 26336
rect 13817 26327 13875 26333
rect 13906 26324 13912 26336
rect 13964 26324 13970 26376
rect 17972 26373 18000 26540
rect 19426 26528 19432 26580
rect 19484 26528 19490 26580
rect 28350 26528 28356 26580
rect 28408 26528 28414 26580
rect 30101 26571 30159 26577
rect 30101 26537 30113 26571
rect 30147 26568 30159 26571
rect 31110 26568 31116 26580
rect 30147 26540 31116 26568
rect 30147 26537 30159 26540
rect 30101 26531 30159 26537
rect 31110 26528 31116 26540
rect 31168 26528 31174 26580
rect 36446 26528 36452 26580
rect 36504 26528 36510 26580
rect 37826 26528 37832 26580
rect 37884 26568 37890 26580
rect 37921 26571 37979 26577
rect 37921 26568 37933 26571
rect 37884 26540 37933 26568
rect 37884 26528 37890 26540
rect 37921 26537 37933 26540
rect 37967 26537 37979 26571
rect 37921 26531 37979 26537
rect 41956 26571 42014 26577
rect 41956 26537 41968 26571
rect 42002 26568 42014 26571
rect 42150 26568 42156 26580
rect 42002 26540 42156 26568
rect 42002 26537 42014 26540
rect 41956 26531 42014 26537
rect 42150 26528 42156 26540
rect 42208 26528 42214 26580
rect 43441 26571 43499 26577
rect 43441 26537 43453 26571
rect 43487 26568 43499 26571
rect 43806 26568 43812 26580
rect 43487 26540 43812 26568
rect 43487 26537 43499 26540
rect 43441 26531 43499 26537
rect 43806 26528 43812 26540
rect 43864 26528 43870 26580
rect 21269 26503 21327 26509
rect 21269 26500 21281 26503
rect 21100 26472 21281 26500
rect 20901 26435 20959 26441
rect 20901 26401 20913 26435
rect 20947 26432 20959 26435
rect 21100 26432 21128 26472
rect 21269 26469 21281 26472
rect 21315 26469 21327 26503
rect 23106 26500 23112 26512
rect 21269 26463 21327 26469
rect 21928 26472 23112 26500
rect 20947 26404 21128 26432
rect 21177 26435 21235 26441
rect 20947 26401 20959 26404
rect 20901 26395 20959 26401
rect 21177 26401 21189 26435
rect 21223 26432 21235 26435
rect 21634 26432 21640 26444
rect 21223 26404 21640 26432
rect 21223 26401 21235 26404
rect 21177 26395 21235 26401
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26364 14519 26367
rect 15197 26367 15255 26373
rect 15197 26364 15209 26367
rect 14507 26336 15209 26364
rect 14507 26333 14519 26336
rect 14461 26327 14519 26333
rect 15197 26333 15209 26336
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 17957 26367 18015 26373
rect 17957 26333 17969 26367
rect 18003 26333 18015 26367
rect 17957 26327 18015 26333
rect 21266 26324 21272 26376
rect 21324 26364 21330 26376
rect 21453 26367 21511 26373
rect 21453 26364 21465 26367
rect 21324 26336 21465 26364
rect 21324 26324 21330 26336
rect 21453 26333 21465 26336
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 10652 26268 12664 26296
rect 12713 26299 12771 26305
rect 10652 26256 10658 26268
rect 12713 26265 12725 26299
rect 12759 26296 12771 26299
rect 13173 26299 13231 26305
rect 13173 26296 13185 26299
rect 12759 26268 13185 26296
rect 12759 26265 12771 26268
rect 12713 26259 12771 26265
rect 13173 26265 13185 26268
rect 13219 26265 13231 26299
rect 16209 26299 16267 26305
rect 16209 26296 16221 26299
rect 13173 26259 13231 26265
rect 14016 26268 16221 26296
rect 12066 26188 12072 26240
rect 12124 26188 12130 26240
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 14016 26228 14044 26268
rect 16209 26265 16221 26268
rect 16255 26296 16267 26299
rect 16574 26296 16580 26308
rect 16255 26268 16580 26296
rect 16255 26265 16267 26268
rect 16209 26259 16267 26265
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 16942 26256 16948 26308
rect 17000 26296 17006 26308
rect 21928 26296 21956 26472
rect 23106 26460 23112 26472
rect 23164 26460 23170 26512
rect 23474 26392 23480 26444
rect 23532 26392 23538 26444
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 23624 26336 23704 26364
rect 23624 26324 23630 26336
rect 23676 26305 23704 26336
rect 28258 26324 28264 26376
rect 28316 26324 28322 26376
rect 28368 26373 28396 26528
rect 29086 26460 29092 26512
rect 29144 26500 29150 26512
rect 29454 26500 29460 26512
rect 29144 26472 29460 26500
rect 29144 26460 29150 26472
rect 29454 26460 29460 26472
rect 29512 26460 29518 26512
rect 29730 26460 29736 26512
rect 29788 26500 29794 26512
rect 29825 26503 29883 26509
rect 29825 26500 29837 26503
rect 29788 26472 29837 26500
rect 29788 26460 29794 26472
rect 29825 26469 29837 26472
rect 29871 26469 29883 26503
rect 29825 26463 29883 26469
rect 30745 26503 30803 26509
rect 30745 26469 30757 26503
rect 30791 26500 30803 26503
rect 32122 26500 32128 26512
rect 30791 26472 32128 26500
rect 30791 26469 30803 26472
rect 30745 26463 30803 26469
rect 32122 26460 32128 26472
rect 32180 26460 32186 26512
rect 35437 26503 35495 26509
rect 35437 26469 35449 26503
rect 35483 26469 35495 26503
rect 35437 26463 35495 26469
rect 29546 26392 29552 26444
rect 29604 26432 29610 26444
rect 29604 26404 29960 26432
rect 29604 26392 29610 26404
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 28813 26367 28871 26373
rect 28813 26333 28825 26367
rect 28859 26333 28871 26367
rect 28813 26327 28871 26333
rect 17000 26268 19656 26296
rect 20470 26268 21956 26296
rect 23661 26299 23719 26305
rect 17000 26256 17006 26268
rect 13872 26200 14044 26228
rect 13872 26188 13878 26200
rect 14090 26188 14096 26240
rect 14148 26188 14154 26240
rect 14550 26188 14556 26240
rect 14608 26188 14614 26240
rect 19628 26228 19656 26268
rect 20548 26228 20576 26268
rect 23661 26265 23673 26299
rect 23707 26296 23719 26299
rect 25406 26296 25412 26308
rect 23707 26268 25412 26296
rect 23707 26265 23719 26268
rect 23661 26259 23719 26265
rect 25406 26256 25412 26268
rect 25464 26256 25470 26308
rect 28169 26299 28227 26305
rect 28169 26265 28181 26299
rect 28215 26296 28227 26299
rect 28828 26296 28856 26327
rect 28994 26324 29000 26376
rect 29052 26364 29058 26376
rect 29932 26373 29960 26404
rect 30466 26392 30472 26444
rect 30524 26392 30530 26444
rect 33870 26392 33876 26444
rect 33928 26392 33934 26444
rect 35452 26432 35480 26463
rect 34256 26404 35480 26432
rect 36464 26432 36492 26528
rect 36725 26435 36783 26441
rect 36725 26432 36737 26435
rect 36464 26404 36737 26432
rect 29089 26367 29147 26373
rect 29089 26364 29101 26367
rect 29052 26336 29101 26364
rect 29052 26324 29058 26336
rect 29089 26333 29101 26336
rect 29135 26333 29147 26367
rect 29089 26327 29147 26333
rect 29273 26367 29331 26373
rect 29273 26333 29285 26367
rect 29319 26364 29331 26367
rect 29641 26367 29699 26373
rect 29641 26364 29653 26367
rect 29319 26336 29653 26364
rect 29319 26333 29331 26336
rect 29273 26327 29331 26333
rect 29641 26333 29653 26336
rect 29687 26333 29699 26367
rect 29641 26327 29699 26333
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 30377 26367 30435 26373
rect 30377 26333 30389 26367
rect 30423 26333 30435 26367
rect 30377 26327 30435 26333
rect 31481 26367 31539 26373
rect 31481 26333 31493 26367
rect 31527 26364 31539 26367
rect 31527 26336 32168 26364
rect 31527 26333 31539 26336
rect 31481 26327 31539 26333
rect 28215 26268 28856 26296
rect 28905 26299 28963 26305
rect 28215 26265 28227 26268
rect 28169 26259 28227 26265
rect 28905 26265 28917 26299
rect 28951 26296 28963 26299
rect 29178 26296 29184 26308
rect 28951 26268 29184 26296
rect 28951 26265 28963 26268
rect 28905 26259 28963 26265
rect 29178 26256 29184 26268
rect 29236 26256 29242 26308
rect 29748 26296 29776 26327
rect 30392 26296 30420 26327
rect 29288 26268 30420 26296
rect 29288 26240 29316 26268
rect 19628 26200 20576 26228
rect 21634 26188 21640 26240
rect 21692 26228 21698 26240
rect 23290 26228 23296 26240
rect 21692 26200 23296 26228
rect 21692 26188 21698 26200
rect 23290 26188 23296 26200
rect 23348 26188 23354 26240
rect 23566 26188 23572 26240
rect 23624 26188 23630 26240
rect 24026 26188 24032 26240
rect 24084 26188 24090 26240
rect 28442 26188 28448 26240
rect 28500 26188 28506 26240
rect 29270 26188 29276 26240
rect 29328 26188 29334 26240
rect 32030 26188 32036 26240
rect 32088 26188 32094 26240
rect 32140 26237 32168 26336
rect 33962 26324 33968 26376
rect 34020 26324 34026 26376
rect 34256 26373 34284 26404
rect 36725 26401 36737 26404
rect 36771 26401 36783 26435
rect 36725 26395 36783 26401
rect 40126 26392 40132 26444
rect 40184 26392 40190 26444
rect 41693 26435 41751 26441
rect 41693 26401 41705 26435
rect 41739 26432 41751 26435
rect 42334 26432 42340 26444
rect 41739 26404 42340 26432
rect 41739 26401 41751 26404
rect 41693 26395 41751 26401
rect 42334 26392 42340 26404
rect 42392 26432 42398 26444
rect 44266 26432 44272 26444
rect 42392 26404 44272 26432
rect 42392 26392 42398 26404
rect 44266 26392 44272 26404
rect 44324 26392 44330 26444
rect 34241 26367 34299 26373
rect 34241 26333 34253 26367
rect 34287 26333 34299 26367
rect 34241 26327 34299 26333
rect 34333 26367 34391 26373
rect 34333 26333 34345 26367
rect 34379 26333 34391 26367
rect 35253 26367 35311 26373
rect 35253 26364 35265 26367
rect 34333 26327 34391 26333
rect 34532 26336 35265 26364
rect 32582 26256 32588 26308
rect 32640 26256 32646 26308
rect 33594 26256 33600 26308
rect 33652 26256 33658 26308
rect 34054 26256 34060 26308
rect 34112 26296 34118 26308
rect 34149 26299 34207 26305
rect 34149 26296 34161 26299
rect 34112 26268 34161 26296
rect 34112 26256 34118 26268
rect 34149 26265 34161 26268
rect 34195 26265 34207 26299
rect 34348 26296 34376 26327
rect 34149 26259 34207 26265
rect 34256 26268 34376 26296
rect 34256 26240 34284 26268
rect 32125 26231 32183 26237
rect 32125 26197 32137 26231
rect 32171 26228 32183 26231
rect 32766 26228 32772 26240
rect 32171 26200 32772 26228
rect 32171 26197 32183 26200
rect 32125 26191 32183 26197
rect 32766 26188 32772 26200
rect 32824 26188 32830 26240
rect 34238 26188 34244 26240
rect 34296 26188 34302 26240
rect 34532 26237 34560 26336
rect 35253 26333 35265 26336
rect 35299 26333 35311 26367
rect 35253 26327 35311 26333
rect 35434 26324 35440 26376
rect 35492 26364 35498 26376
rect 35989 26367 36047 26373
rect 35989 26364 36001 26367
rect 35492 26336 36001 26364
rect 35492 26324 35498 26336
rect 35989 26333 36001 26336
rect 36035 26333 36047 26367
rect 35989 26327 36047 26333
rect 37090 26324 37096 26376
rect 37148 26324 37154 26376
rect 38010 26324 38016 26376
rect 38068 26364 38074 26376
rect 38473 26367 38531 26373
rect 38473 26364 38485 26367
rect 38068 26336 38485 26364
rect 38068 26324 38074 26336
rect 38473 26333 38485 26336
rect 38519 26333 38531 26367
rect 38473 26327 38531 26333
rect 39853 26367 39911 26373
rect 39853 26333 39865 26367
rect 39899 26333 39911 26367
rect 39853 26327 39911 26333
rect 37642 26256 37648 26308
rect 37700 26296 37706 26308
rect 37737 26299 37795 26305
rect 37737 26296 37749 26299
rect 37700 26268 37749 26296
rect 37700 26256 37706 26268
rect 37737 26265 37749 26268
rect 37783 26265 37795 26299
rect 37737 26259 37795 26265
rect 38102 26256 38108 26308
rect 38160 26296 38166 26308
rect 39868 26296 39896 26327
rect 41138 26324 41144 26376
rect 41196 26364 41202 26376
rect 41196 26336 41736 26364
rect 41196 26324 41202 26336
rect 40034 26296 40040 26308
rect 38160 26268 40040 26296
rect 38160 26256 38166 26268
rect 40034 26256 40040 26268
rect 40092 26256 40098 26308
rect 41708 26296 41736 26336
rect 43254 26296 43260 26308
rect 41708 26268 42380 26296
rect 43194 26268 43260 26296
rect 34517 26231 34575 26237
rect 34517 26197 34529 26231
rect 34563 26197 34575 26231
rect 34517 26191 34575 26197
rect 34698 26188 34704 26240
rect 34756 26188 34762 26240
rect 35894 26188 35900 26240
rect 35952 26228 35958 26240
rect 36173 26231 36231 26237
rect 36173 26228 36185 26231
rect 35952 26200 36185 26228
rect 35952 26188 35958 26200
rect 36173 26197 36185 26200
rect 36219 26197 36231 26231
rect 36173 26191 36231 26197
rect 41598 26188 41604 26240
rect 41656 26188 41662 26240
rect 42352 26228 42380 26268
rect 43254 26256 43260 26268
rect 43312 26256 43318 26308
rect 43272 26228 43300 26256
rect 42352 26200 43300 26228
rect 1104 26138 44620 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 44620 26138
rect 1104 26064 44620 26086
rect 5718 25984 5724 26036
rect 5776 25984 5782 26036
rect 7834 25984 7840 26036
rect 7892 26024 7898 26036
rect 7892 25996 9720 26024
rect 7892 25984 7898 25996
rect 5736 25888 5764 25984
rect 9582 25956 9588 25968
rect 8602 25928 9588 25956
rect 9582 25916 9588 25928
rect 9640 25916 9646 25968
rect 9692 25956 9720 25996
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 10061 26027 10119 26033
rect 10061 26024 10073 26027
rect 9824 25996 10073 26024
rect 9824 25984 9830 25996
rect 10061 25993 10073 25996
rect 10107 25993 10119 26027
rect 10061 25987 10119 25993
rect 10229 26027 10287 26033
rect 10229 25993 10241 26027
rect 10275 25993 10287 26027
rect 10229 25987 10287 25993
rect 9861 25959 9919 25965
rect 9861 25956 9873 25959
rect 9692 25928 9873 25956
rect 9861 25925 9873 25928
rect 9907 25925 9919 25959
rect 10244 25956 10272 25987
rect 12066 25984 12072 26036
rect 12124 25984 12130 26036
rect 13357 26027 13415 26033
rect 13357 25993 13369 26027
rect 13403 26024 13415 26027
rect 13906 26024 13912 26036
rect 13403 25996 13912 26024
rect 13403 25993 13415 25996
rect 13357 25987 13415 25993
rect 11885 25959 11943 25965
rect 10244 25928 11008 25956
rect 9861 25919 9919 25925
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 5736 25860 6561 25888
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 9030 25848 9036 25900
rect 9088 25888 9094 25900
rect 9769 25891 9827 25897
rect 9769 25888 9781 25891
rect 9088 25860 9781 25888
rect 9088 25848 9094 25860
rect 9769 25857 9781 25860
rect 9815 25888 9827 25891
rect 10505 25891 10563 25897
rect 10505 25888 10517 25891
rect 9815 25860 10517 25888
rect 9815 25857 9827 25860
rect 9769 25851 9827 25857
rect 10505 25857 10517 25860
rect 10551 25888 10563 25891
rect 10594 25888 10600 25900
rect 10551 25860 10600 25888
rect 10551 25857 10563 25860
rect 10505 25851 10563 25857
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 10980 25897 11008 25928
rect 11885 25925 11897 25959
rect 11931 25956 11943 25959
rect 12084 25956 12112 25984
rect 11931 25928 12112 25956
rect 11931 25925 11943 25928
rect 11885 25919 11943 25925
rect 12434 25916 12440 25968
rect 12492 25916 12498 25968
rect 13556 25897 13584 25996
rect 13906 25984 13912 25996
rect 13964 25984 13970 26036
rect 14550 25984 14556 26036
rect 14608 25984 14614 26036
rect 15838 25984 15844 26036
rect 15896 25984 15902 26036
rect 22373 26027 22431 26033
rect 19996 25996 22324 26024
rect 14568 25956 14596 25984
rect 15654 25956 15660 25968
rect 13648 25928 14596 25956
rect 15594 25928 15660 25956
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25857 10747 25891
rect 10689 25851 10747 25857
rect 10965 25891 11023 25897
rect 10965 25857 10977 25891
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 13541 25891 13599 25897
rect 13541 25857 13553 25891
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 5810 25780 5816 25832
rect 5868 25820 5874 25832
rect 6638 25820 6644 25832
rect 5868 25792 6644 25820
rect 5868 25780 5874 25792
rect 6638 25780 6644 25792
rect 6696 25820 6702 25832
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6696 25792 7205 25820
rect 6696 25780 6702 25792
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25820 7619 25823
rect 7926 25820 7932 25832
rect 7607 25792 7932 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 7926 25780 7932 25792
rect 7984 25780 7990 25832
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 10704 25820 10732 25851
rect 9548 25792 10732 25820
rect 9548 25780 9554 25792
rect 10321 25755 10379 25761
rect 10321 25752 10333 25755
rect 10060 25724 10333 25752
rect 6178 25644 6184 25696
rect 6236 25684 6242 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 6236 25656 6377 25684
rect 6236 25644 6242 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 9122 25644 9128 25696
rect 9180 25644 9186 25696
rect 10060 25693 10088 25724
rect 10321 25721 10333 25724
rect 10367 25721 10379 25755
rect 10704 25752 10732 25792
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 11609 25823 11667 25829
rect 11609 25820 11621 25823
rect 11112 25792 11621 25820
rect 11112 25780 11118 25792
rect 11609 25789 11621 25792
rect 11655 25789 11667 25823
rect 12342 25820 12348 25832
rect 11609 25783 11667 25789
rect 11716 25792 12348 25820
rect 11716 25752 11744 25792
rect 12342 25780 12348 25792
rect 12400 25820 12406 25832
rect 13648 25820 13676 25928
rect 15654 25916 15660 25928
rect 15712 25916 15718 25968
rect 16758 25916 16764 25968
rect 16816 25956 16822 25968
rect 16816 25928 17540 25956
rect 16816 25916 16822 25928
rect 13722 25848 13728 25900
rect 13780 25848 13786 25900
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 17512 25897 17540 25928
rect 18046 25916 18052 25968
rect 18104 25956 18110 25968
rect 19996 25956 20024 25996
rect 18104 25928 20102 25956
rect 18104 25916 18110 25928
rect 17497 25891 17555 25897
rect 16632 25860 17448 25888
rect 16632 25848 16638 25860
rect 12400 25792 13676 25820
rect 12400 25780 12406 25792
rect 13814 25780 13820 25832
rect 13872 25820 13878 25832
rect 14093 25823 14151 25829
rect 14093 25820 14105 25823
rect 13872 25792 14105 25820
rect 13872 25780 13878 25792
rect 14093 25789 14105 25792
rect 14139 25789 14151 25823
rect 14093 25783 14151 25789
rect 14366 25780 14372 25832
rect 14424 25780 14430 25832
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25789 17371 25823
rect 17420 25820 17448 25860
rect 17497 25857 17509 25891
rect 17543 25857 17555 25891
rect 17497 25851 17555 25857
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22189 25891 22247 25897
rect 22189 25888 22201 25891
rect 22152 25860 22201 25888
rect 22152 25848 22158 25860
rect 22189 25857 22201 25860
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 19337 25823 19395 25829
rect 19337 25820 19349 25823
rect 17420 25792 19349 25820
rect 17313 25783 17371 25789
rect 19337 25789 19349 25792
rect 19383 25789 19395 25823
rect 19337 25783 19395 25789
rect 10704 25724 11744 25752
rect 17328 25752 17356 25783
rect 19610 25780 19616 25832
rect 19668 25780 19674 25832
rect 17402 25752 17408 25764
rect 17328 25724 17408 25752
rect 10321 25715 10379 25721
rect 17402 25712 17408 25724
rect 17460 25712 17466 25764
rect 22296 25752 22324 25996
rect 22373 25993 22385 26027
rect 22419 26024 22431 26027
rect 22649 26027 22707 26033
rect 22649 26024 22661 26027
rect 22419 25996 22661 26024
rect 22419 25993 22431 25996
rect 22373 25987 22431 25993
rect 22649 25993 22661 25996
rect 22695 26024 22707 26027
rect 23566 26024 23572 26036
rect 22695 25996 23572 26024
rect 22695 25993 22707 25996
rect 22649 25987 22707 25993
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 23842 25984 23848 26036
rect 23900 25984 23906 26036
rect 28258 25984 28264 26036
rect 28316 26024 28322 26036
rect 28721 26027 28779 26033
rect 28721 26024 28733 26027
rect 28316 25996 28733 26024
rect 28316 25984 28322 25996
rect 28721 25993 28733 25996
rect 28767 26024 28779 26027
rect 29365 26027 29423 26033
rect 28767 25996 29132 26024
rect 28767 25993 28779 25996
rect 28721 25987 28779 25993
rect 23860 25956 23888 25984
rect 25314 25956 25320 25968
rect 22480 25928 23888 25956
rect 24886 25928 25320 25956
rect 22480 25900 22508 25928
rect 25314 25916 25320 25928
rect 25372 25916 25378 25968
rect 25406 25916 25412 25968
rect 25464 25916 25470 25968
rect 28537 25959 28595 25965
rect 28537 25925 28549 25959
rect 28583 25956 28595 25959
rect 28905 25959 28963 25965
rect 28905 25956 28917 25959
rect 28583 25928 28917 25956
rect 28583 25925 28595 25928
rect 28537 25919 28595 25925
rect 28905 25925 28917 25928
rect 28951 25956 28963 25959
rect 28994 25956 29000 25968
rect 28951 25928 29000 25956
rect 28951 25925 28963 25928
rect 28905 25919 28963 25925
rect 28994 25916 29000 25928
rect 29052 25916 29058 25968
rect 22462 25848 22468 25900
rect 22520 25848 22526 25900
rect 23290 25848 23296 25900
rect 23348 25888 23354 25900
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 23348 25860 23397 25888
rect 23348 25848 23354 25860
rect 23385 25857 23397 25860
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 26142 25848 26148 25900
rect 26200 25848 26206 25900
rect 28353 25891 28411 25897
rect 28353 25888 28365 25891
rect 26712 25860 28365 25888
rect 23198 25780 23204 25832
rect 23256 25780 23262 25832
rect 23658 25780 23664 25832
rect 23716 25780 23722 25832
rect 25866 25780 25872 25832
rect 25924 25780 25930 25832
rect 22296 25724 23520 25752
rect 23492 25696 23520 25724
rect 26712 25696 26740 25860
rect 28092 25752 28120 25860
rect 28353 25857 28365 25860
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 28442 25848 28448 25900
rect 28500 25888 28506 25900
rect 29104 25897 29132 25996
rect 29365 25993 29377 26027
rect 29411 26024 29423 26027
rect 29454 26024 29460 26036
rect 29411 25996 29460 26024
rect 29411 25993 29423 25996
rect 29365 25987 29423 25993
rect 29454 25984 29460 25996
rect 29512 25984 29518 26036
rect 30101 26027 30159 26033
rect 30101 25993 30113 26027
rect 30147 26024 30159 26027
rect 30466 26024 30472 26036
rect 30147 25996 30472 26024
rect 30147 25993 30159 25996
rect 30101 25987 30159 25993
rect 30466 25984 30472 25996
rect 30524 25984 30530 26036
rect 31938 25984 31944 26036
rect 31996 26024 32002 26036
rect 32677 26027 32735 26033
rect 31996 25996 32628 26024
rect 31996 25984 32002 25996
rect 29270 25916 29276 25968
rect 29328 25916 29334 25968
rect 29546 25916 29552 25968
rect 29604 25956 29610 25968
rect 29604 25928 29868 25956
rect 29604 25916 29610 25928
rect 28629 25891 28687 25897
rect 28629 25888 28641 25891
rect 28500 25860 28641 25888
rect 28500 25848 28506 25860
rect 28629 25857 28641 25860
rect 28675 25857 28687 25891
rect 28629 25851 28687 25857
rect 28813 25891 28871 25897
rect 28813 25857 28825 25891
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 29089 25891 29147 25897
rect 29089 25857 29101 25891
rect 29135 25857 29147 25891
rect 29089 25851 29147 25857
rect 28169 25823 28227 25829
rect 28169 25789 28181 25823
rect 28215 25820 28227 25823
rect 28460 25820 28488 25848
rect 28215 25792 28488 25820
rect 28215 25789 28227 25792
rect 28169 25783 28227 25789
rect 28828 25752 28856 25851
rect 29730 25848 29736 25900
rect 29788 25848 29794 25900
rect 29840 25897 29868 25928
rect 32030 25916 32036 25968
rect 32088 25956 32094 25968
rect 32401 25959 32459 25965
rect 32401 25956 32413 25959
rect 32088 25928 32413 25956
rect 32088 25916 32094 25928
rect 32401 25925 32413 25928
rect 32447 25925 32459 25959
rect 32401 25919 32459 25925
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 31570 25848 31576 25900
rect 31628 25848 31634 25900
rect 32122 25848 32128 25900
rect 32180 25848 32186 25900
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 29178 25780 29184 25832
rect 29236 25820 29242 25832
rect 30101 25823 30159 25829
rect 30101 25820 30113 25823
rect 29236 25792 30113 25820
rect 29236 25780 29242 25792
rect 30101 25789 30113 25792
rect 30147 25789 30159 25823
rect 31588 25820 31616 25848
rect 32324 25820 32352 25851
rect 32398 25820 32404 25832
rect 31588 25792 32404 25820
rect 30101 25783 30159 25789
rect 32398 25780 32404 25792
rect 32456 25780 32462 25832
rect 28092 25724 28856 25752
rect 32306 25712 32312 25764
rect 32364 25752 32370 25764
rect 32508 25752 32536 25851
rect 32600 25820 32628 25996
rect 32677 25993 32689 26027
rect 32723 26024 32735 26027
rect 33594 26024 33600 26036
rect 32723 25996 33600 26024
rect 32723 25993 32735 25996
rect 32677 25987 32735 25993
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 34698 26024 34704 26036
rect 33796 25996 34704 26024
rect 32858 25916 32864 25968
rect 32916 25916 32922 25968
rect 33796 25965 33824 25996
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 35253 26027 35311 26033
rect 35253 25993 35265 26027
rect 35299 26024 35311 26027
rect 35434 26024 35440 26036
rect 35299 25996 35440 26024
rect 35299 25993 35311 25996
rect 35253 25987 35311 25993
rect 35434 25984 35440 25996
rect 35492 25984 35498 26036
rect 35986 26024 35992 26036
rect 35544 25996 35992 26024
rect 33781 25959 33839 25965
rect 33781 25925 33793 25959
rect 33827 25925 33839 25959
rect 35544 25956 35572 25996
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 37090 25984 37096 26036
rect 37148 25984 37154 26036
rect 42705 26027 42763 26033
rect 42705 25993 42717 26027
rect 42751 26024 42763 26027
rect 42886 26024 42892 26036
rect 42751 25996 42892 26024
rect 42751 25993 42763 25996
rect 42705 25987 42763 25993
rect 42886 25984 42892 25996
rect 42944 25984 42950 26036
rect 43165 26027 43223 26033
rect 43165 25993 43177 26027
rect 43211 25993 43223 26027
rect 43165 25987 43223 25993
rect 33781 25919 33839 25925
rect 35268 25928 35572 25956
rect 35621 25959 35679 25965
rect 32766 25848 32772 25900
rect 32824 25848 32830 25900
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 35268 25888 35296 25928
rect 35621 25925 35633 25959
rect 35667 25956 35679 25959
rect 35894 25956 35900 25968
rect 35667 25928 35900 25956
rect 35667 25925 35679 25928
rect 35621 25919 35679 25925
rect 35894 25916 35900 25928
rect 35952 25916 35958 25968
rect 36004 25956 36032 25984
rect 40126 25956 40132 25968
rect 36004 25928 36110 25956
rect 39606 25928 40132 25956
rect 40126 25916 40132 25928
rect 40184 25956 40190 25968
rect 41138 25956 41144 25968
rect 40184 25928 41144 25956
rect 40184 25916 40190 25928
rect 41138 25916 41144 25928
rect 41196 25916 41202 25968
rect 34848 25860 35296 25888
rect 34848 25848 34854 25860
rect 35342 25848 35348 25900
rect 35400 25848 35406 25900
rect 37366 25848 37372 25900
rect 37424 25888 37430 25900
rect 37829 25891 37887 25897
rect 37829 25888 37841 25891
rect 37424 25860 37841 25888
rect 37424 25848 37430 25860
rect 37829 25857 37841 25860
rect 37875 25857 37887 25891
rect 37829 25851 37887 25857
rect 41598 25848 41604 25900
rect 41656 25888 41662 25900
rect 41693 25891 41751 25897
rect 41693 25888 41705 25891
rect 41656 25860 41705 25888
rect 41656 25848 41662 25860
rect 41693 25857 41705 25860
rect 41739 25857 41751 25891
rect 41693 25851 41751 25857
rect 42797 25891 42855 25897
rect 42797 25857 42809 25891
rect 42843 25888 42855 25891
rect 43070 25888 43076 25900
rect 42843 25860 43076 25888
rect 42843 25857 42855 25860
rect 42797 25851 42855 25857
rect 43070 25848 43076 25860
rect 43128 25848 43134 25900
rect 43180 25888 43208 25987
rect 43257 25891 43315 25897
rect 43257 25888 43269 25891
rect 43180 25860 43269 25888
rect 43257 25857 43269 25860
rect 43303 25857 43315 25891
rect 43257 25851 43315 25857
rect 32674 25820 32680 25832
rect 32600 25792 32680 25820
rect 32674 25780 32680 25792
rect 32732 25820 32738 25832
rect 33505 25823 33563 25829
rect 33505 25820 33517 25823
rect 32732 25792 33517 25820
rect 32732 25780 32738 25792
rect 33505 25789 33517 25792
rect 33551 25789 33563 25823
rect 35360 25820 35388 25848
rect 35710 25820 35716 25832
rect 35360 25792 35716 25820
rect 33505 25783 33563 25789
rect 35710 25780 35716 25792
rect 35768 25780 35774 25832
rect 38102 25780 38108 25832
rect 38160 25780 38166 25832
rect 38378 25780 38384 25832
rect 38436 25780 38442 25832
rect 39853 25823 39911 25829
rect 39853 25789 39865 25823
rect 39899 25820 39911 25823
rect 39945 25823 40003 25829
rect 39945 25820 39957 25823
rect 39899 25792 39957 25820
rect 39899 25789 39911 25792
rect 39853 25783 39911 25789
rect 39945 25789 39957 25792
rect 39991 25789 40003 25823
rect 39945 25783 40003 25789
rect 42613 25823 42671 25829
rect 42613 25789 42625 25823
rect 42659 25820 42671 25823
rect 42886 25820 42892 25832
rect 42659 25792 42892 25820
rect 42659 25789 42671 25792
rect 42613 25783 42671 25789
rect 42886 25780 42892 25792
rect 42944 25820 42950 25832
rect 43162 25820 43168 25832
rect 42944 25792 43168 25820
rect 42944 25780 42950 25792
rect 43162 25780 43168 25792
rect 43220 25780 43226 25832
rect 33226 25752 33232 25764
rect 32364 25724 33232 25752
rect 32364 25712 32370 25724
rect 33226 25712 33232 25724
rect 33284 25712 33290 25764
rect 10045 25687 10103 25693
rect 10045 25653 10057 25687
rect 10091 25653 10103 25687
rect 10045 25647 10103 25653
rect 10686 25644 10692 25696
rect 10744 25684 10750 25696
rect 10781 25687 10839 25693
rect 10781 25684 10793 25687
rect 10744 25656 10793 25684
rect 10744 25644 10750 25656
rect 10781 25653 10793 25656
rect 10827 25653 10839 25687
rect 10781 25647 10839 25653
rect 13906 25644 13912 25696
rect 13964 25644 13970 25696
rect 21082 25644 21088 25696
rect 21140 25644 21146 25696
rect 22002 25644 22008 25696
rect 22060 25644 22066 25696
rect 23474 25644 23480 25696
rect 23532 25644 23538 25696
rect 25961 25687 26019 25693
rect 25961 25653 25973 25687
rect 26007 25684 26019 25687
rect 26050 25684 26056 25696
rect 26007 25656 26056 25684
rect 26007 25653 26019 25656
rect 25961 25647 26019 25653
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 26326 25644 26332 25696
rect 26384 25644 26390 25696
rect 26694 25644 26700 25696
rect 26752 25644 26758 25696
rect 28994 25644 29000 25696
rect 29052 25684 29058 25696
rect 29638 25684 29644 25696
rect 29052 25656 29644 25684
rect 29052 25644 29058 25656
rect 29638 25644 29644 25656
rect 29696 25644 29702 25696
rect 29730 25644 29736 25696
rect 29788 25684 29794 25696
rect 29917 25687 29975 25693
rect 29917 25684 29929 25687
rect 29788 25656 29929 25684
rect 29788 25644 29794 25656
rect 29917 25653 29929 25656
rect 29963 25653 29975 25687
rect 29917 25647 29975 25653
rect 37274 25644 37280 25696
rect 37332 25644 37338 25696
rect 40586 25644 40592 25696
rect 40644 25644 40650 25696
rect 41046 25644 41052 25696
rect 41104 25684 41110 25696
rect 41141 25687 41199 25693
rect 41141 25684 41153 25687
rect 41104 25656 41153 25684
rect 41104 25644 41110 25656
rect 41141 25653 41153 25656
rect 41187 25653 41199 25687
rect 41141 25647 41199 25653
rect 43438 25644 43444 25696
rect 43496 25644 43502 25696
rect 1104 25594 44620 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 44620 25594
rect 1104 25520 44620 25542
rect 7926 25440 7932 25492
rect 7984 25440 7990 25492
rect 9122 25440 9128 25492
rect 9180 25440 9186 25492
rect 9582 25440 9588 25492
rect 9640 25440 9646 25492
rect 10686 25440 10692 25492
rect 10744 25489 10750 25492
rect 10744 25483 10759 25489
rect 10747 25449 10759 25483
rect 10744 25443 10759 25449
rect 10744 25440 10750 25443
rect 13906 25440 13912 25492
rect 13964 25440 13970 25492
rect 14277 25483 14335 25489
rect 14277 25449 14289 25483
rect 14323 25480 14335 25483
rect 14366 25480 14372 25492
rect 14323 25452 14372 25480
rect 14323 25449 14335 25452
rect 14277 25443 14335 25449
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 18874 25440 18880 25492
rect 18932 25440 18938 25492
rect 19610 25440 19616 25492
rect 19668 25480 19674 25492
rect 19981 25483 20039 25489
rect 19981 25480 19993 25483
rect 19668 25452 19993 25480
rect 19668 25440 19674 25452
rect 19981 25449 19993 25452
rect 20027 25449 20039 25483
rect 19981 25443 20039 25449
rect 21082 25440 21088 25492
rect 21140 25440 21146 25492
rect 22462 25480 22468 25492
rect 21376 25452 22468 25480
rect 5810 25304 5816 25356
rect 5868 25304 5874 25356
rect 6089 25347 6147 25353
rect 6089 25313 6101 25347
rect 6135 25344 6147 25347
rect 6178 25344 6184 25356
rect 6135 25316 6184 25344
rect 6135 25313 6147 25316
rect 6089 25307 6147 25313
rect 6178 25304 6184 25316
rect 6236 25304 6242 25356
rect 7834 25236 7840 25288
rect 7892 25236 7898 25288
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25276 8079 25279
rect 9140 25276 9168 25440
rect 9490 25304 9496 25356
rect 9548 25304 9554 25356
rect 9508 25276 9536 25304
rect 8067 25248 9168 25276
rect 9416 25248 9536 25276
rect 8067 25245 8079 25248
rect 8021 25239 8079 25245
rect 8941 25211 8999 25217
rect 7314 25180 8432 25208
rect 7561 25143 7619 25149
rect 7561 25109 7573 25143
rect 7607 25140 7619 25143
rect 8294 25140 8300 25152
rect 7607 25112 8300 25140
rect 7607 25109 7619 25112
rect 7561 25103 7619 25109
rect 8294 25100 8300 25112
rect 8352 25100 8358 25152
rect 8404 25140 8432 25180
rect 8941 25177 8953 25211
rect 8987 25208 8999 25211
rect 9416 25208 9444 25248
rect 8987 25180 9444 25208
rect 8987 25177 8999 25180
rect 8941 25171 8999 25177
rect 9600 25140 9628 25440
rect 13924 25412 13952 25440
rect 13924 25384 19380 25412
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 10965 25347 11023 25353
rect 10965 25344 10977 25347
rect 9732 25316 10977 25344
rect 9732 25304 9738 25316
rect 10965 25313 10977 25316
rect 11011 25344 11023 25347
rect 11054 25344 11060 25356
rect 11011 25316 11060 25344
rect 11011 25313 11023 25316
rect 10965 25307 11023 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 11698 25304 11704 25356
rect 11756 25344 11762 25356
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 11756 25316 12817 25344
rect 11756 25304 11762 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 12805 25307 12863 25313
rect 17770 25304 17776 25356
rect 17828 25304 17834 25356
rect 17880 25316 19288 25344
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 14090 25236 14096 25288
rect 14148 25236 14154 25288
rect 14734 25236 14740 25288
rect 14792 25276 14798 25288
rect 17880 25276 17908 25316
rect 14792 25248 17908 25276
rect 14792 25236 14798 25248
rect 18414 25236 18420 25288
rect 18472 25276 18478 25288
rect 19260 25285 19288 25316
rect 18601 25279 18659 25285
rect 18601 25276 18613 25279
rect 18472 25248 18613 25276
rect 18472 25236 18478 25248
rect 18601 25245 18613 25248
rect 18647 25276 18659 25279
rect 18785 25279 18843 25285
rect 18785 25276 18797 25279
rect 18647 25248 18797 25276
rect 18647 25245 18659 25248
rect 18601 25239 18659 25245
rect 18785 25245 18797 25248
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 19352 25276 19380 25384
rect 20717 25347 20775 25353
rect 20717 25344 20729 25347
rect 20364 25316 20729 25344
rect 20165 25279 20223 25285
rect 20165 25276 20177 25279
rect 19352 25248 20177 25276
rect 19245 25239 19303 25245
rect 20165 25245 20177 25248
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 11330 25168 11336 25220
rect 11388 25168 11394 25220
rect 17497 25211 17555 25217
rect 17497 25177 17509 25211
rect 17543 25208 17555 25211
rect 18049 25211 18107 25217
rect 18049 25208 18061 25211
rect 17543 25180 18061 25208
rect 17543 25177 17555 25180
rect 17497 25171 17555 25177
rect 18049 25177 18061 25180
rect 18095 25177 18107 25211
rect 18049 25171 18107 25177
rect 8404 25112 9628 25140
rect 17126 25100 17132 25152
rect 17184 25100 17190 25152
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25140 17647 25143
rect 19242 25140 19248 25152
rect 17635 25112 19248 25140
rect 17635 25109 17647 25112
rect 17589 25103 17647 25109
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 19426 25100 19432 25152
rect 19484 25100 19490 25152
rect 20180 25140 20208 25239
rect 20254 25236 20260 25288
rect 20312 25276 20318 25288
rect 20364 25285 20392 25316
rect 20717 25313 20729 25316
rect 20763 25313 20775 25347
rect 21100 25344 21128 25440
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 21100 25316 21281 25344
rect 20717 25307 20775 25313
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 21269 25307 21327 25313
rect 20349 25279 20407 25285
rect 20349 25276 20361 25279
rect 20312 25248 20361 25276
rect 20312 25236 20318 25248
rect 20349 25245 20361 25248
rect 20395 25245 20407 25279
rect 20349 25239 20407 25245
rect 20441 25279 20499 25285
rect 20441 25245 20453 25279
rect 20487 25276 20499 25279
rect 21376 25276 21404 25452
rect 22462 25440 22468 25452
rect 22520 25440 22526 25492
rect 23198 25440 23204 25492
rect 23256 25480 23262 25492
rect 23477 25483 23535 25489
rect 23477 25480 23489 25483
rect 23256 25452 23489 25480
rect 23256 25440 23262 25452
rect 23477 25449 23489 25452
rect 23523 25449 23535 25483
rect 23477 25443 23535 25449
rect 23569 25483 23627 25489
rect 23569 25449 23581 25483
rect 23615 25480 23627 25483
rect 23658 25480 23664 25492
rect 23615 25452 23664 25480
rect 23615 25449 23627 25452
rect 23569 25443 23627 25449
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 26053 25483 26111 25489
rect 26053 25449 26065 25483
rect 26099 25480 26111 25483
rect 26099 25452 26648 25480
rect 26099 25449 26111 25452
rect 26053 25443 26111 25449
rect 26234 25412 26240 25424
rect 23584 25384 26240 25412
rect 21634 25304 21640 25356
rect 21692 25344 21698 25356
rect 21729 25347 21787 25353
rect 21729 25344 21741 25347
rect 21692 25316 21741 25344
rect 21692 25304 21698 25316
rect 21729 25313 21741 25316
rect 21775 25313 21787 25347
rect 21729 25307 21787 25313
rect 22002 25304 22008 25356
rect 22060 25304 22066 25356
rect 20487 25248 21404 25276
rect 20487 25245 20499 25248
rect 20441 25239 20499 25245
rect 23474 25208 23480 25220
rect 23230 25180 23480 25208
rect 23474 25168 23480 25180
rect 23532 25168 23538 25220
rect 23584 25140 23612 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 26326 25372 26332 25424
rect 26384 25412 26390 25424
rect 26620 25412 26648 25452
rect 26694 25440 26700 25492
rect 26752 25440 26758 25492
rect 28629 25483 28687 25489
rect 28629 25449 28641 25483
rect 28675 25480 28687 25483
rect 28675 25452 29132 25480
rect 28675 25449 28687 25452
rect 28629 25443 28687 25449
rect 28994 25412 29000 25424
rect 26384 25384 26556 25412
rect 26620 25384 29000 25412
rect 26384 25372 26390 25384
rect 25682 25304 25688 25356
rect 25740 25304 25746 25356
rect 26528 25353 26556 25384
rect 28994 25372 29000 25384
rect 29052 25372 29058 25424
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25313 26571 25347
rect 26513 25307 26571 25313
rect 27157 25347 27215 25353
rect 27157 25313 27169 25347
rect 27203 25313 27215 25347
rect 27157 25307 27215 25313
rect 27433 25347 27491 25353
rect 27433 25313 27445 25347
rect 27479 25344 27491 25347
rect 27479 25316 28856 25344
rect 27479 25313 27491 25316
rect 27433 25307 27491 25313
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25276 23811 25279
rect 24026 25276 24032 25288
rect 23799 25248 24032 25276
rect 23799 25245 23811 25248
rect 23753 25239 23811 25245
rect 24026 25236 24032 25248
rect 24084 25236 24090 25288
rect 24210 25236 24216 25288
rect 24268 25276 24274 25288
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 24268 25248 24961 25276
rect 24268 25236 24274 25248
rect 24949 25245 24961 25248
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 25130 25236 25136 25288
rect 25188 25276 25194 25288
rect 25777 25279 25835 25285
rect 25777 25276 25789 25279
rect 25188 25248 25789 25276
rect 25188 25236 25194 25248
rect 25777 25245 25789 25248
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 26234 25236 26240 25288
rect 26292 25276 26298 25288
rect 26421 25279 26479 25285
rect 26421 25276 26433 25279
rect 26292 25248 26433 25276
rect 26292 25236 26298 25248
rect 26421 25245 26433 25248
rect 26467 25245 26479 25279
rect 26421 25239 26479 25245
rect 27065 25279 27123 25285
rect 27065 25245 27077 25279
rect 27111 25245 27123 25279
rect 27172 25276 27200 25307
rect 27706 25276 27712 25288
rect 27172 25248 27712 25276
rect 27065 25239 27123 25245
rect 20180 25112 23612 25140
rect 23658 25100 23664 25152
rect 23716 25140 23722 25152
rect 24397 25143 24455 25149
rect 24397 25140 24409 25143
rect 23716 25112 24409 25140
rect 23716 25100 23722 25112
rect 24397 25109 24409 25112
rect 24443 25109 24455 25143
rect 24397 25103 24455 25109
rect 25866 25100 25872 25152
rect 25924 25140 25930 25152
rect 27080 25140 27108 25239
rect 27706 25236 27712 25248
rect 27764 25236 27770 25288
rect 28552 25285 28580 25316
rect 28828 25285 28856 25316
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25245 28595 25279
rect 28537 25239 28595 25245
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25245 28871 25279
rect 29104 25276 29132 25452
rect 29178 25440 29184 25492
rect 29236 25440 29242 25492
rect 29546 25440 29552 25492
rect 29604 25480 29610 25492
rect 29641 25483 29699 25489
rect 29641 25480 29653 25483
rect 29604 25452 29653 25480
rect 29604 25440 29610 25452
rect 29641 25449 29653 25452
rect 29687 25449 29699 25483
rect 29641 25443 29699 25449
rect 36620 25483 36678 25489
rect 36620 25449 36632 25483
rect 36666 25480 36678 25483
rect 37274 25480 37280 25492
rect 36666 25452 37280 25480
rect 36666 25449 36678 25452
rect 36620 25443 36678 25449
rect 37274 25440 37280 25452
rect 37332 25440 37338 25492
rect 38378 25440 38384 25492
rect 38436 25480 38442 25492
rect 38473 25483 38531 25489
rect 38473 25480 38485 25483
rect 38436 25452 38485 25480
rect 38436 25440 38442 25452
rect 38473 25449 38485 25452
rect 38519 25449 38531 25483
rect 38473 25443 38531 25449
rect 39393 25483 39451 25489
rect 39393 25449 39405 25483
rect 39439 25480 39451 25483
rect 40126 25480 40132 25492
rect 39439 25452 40132 25480
rect 39439 25449 39451 25452
rect 39393 25443 39451 25449
rect 40126 25440 40132 25452
rect 40184 25440 40190 25492
rect 40497 25483 40555 25489
rect 40497 25449 40509 25483
rect 40543 25480 40555 25483
rect 40678 25480 40684 25492
rect 40543 25452 40684 25480
rect 40543 25449 40555 25452
rect 40497 25443 40555 25449
rect 40678 25440 40684 25452
rect 40736 25440 40742 25492
rect 40954 25440 40960 25492
rect 41012 25440 41018 25492
rect 29196 25344 29224 25440
rect 40313 25415 40371 25421
rect 40313 25381 40325 25415
rect 40359 25412 40371 25415
rect 40972 25412 41000 25440
rect 40359 25384 41000 25412
rect 40359 25381 40371 25384
rect 40313 25375 40371 25381
rect 29196 25316 29776 25344
rect 29748 25285 29776 25316
rect 35710 25304 35716 25356
rect 35768 25344 35774 25356
rect 36357 25347 36415 25353
rect 36357 25344 36369 25347
rect 35768 25316 36369 25344
rect 35768 25304 35774 25316
rect 36357 25313 36369 25316
rect 36403 25344 36415 25347
rect 38102 25344 38108 25356
rect 36403 25316 38108 25344
rect 36403 25313 36415 25316
rect 36357 25307 36415 25313
rect 38102 25304 38108 25316
rect 38160 25304 38166 25356
rect 39117 25347 39175 25353
rect 39117 25313 39129 25347
rect 39163 25344 39175 25347
rect 39853 25347 39911 25353
rect 39853 25344 39865 25347
rect 39163 25316 39865 25344
rect 39163 25313 39175 25316
rect 39117 25307 39175 25313
rect 39853 25313 39865 25316
rect 39899 25313 39911 25347
rect 39853 25307 39911 25313
rect 43438 25304 43444 25356
rect 43496 25344 43502 25356
rect 43901 25347 43959 25353
rect 43901 25344 43913 25347
rect 43496 25316 43913 25344
rect 43496 25304 43502 25316
rect 43901 25313 43913 25316
rect 43947 25313 43959 25347
rect 43901 25307 43959 25313
rect 44177 25347 44235 25353
rect 44177 25313 44189 25347
rect 44223 25344 44235 25347
rect 44266 25344 44272 25356
rect 44223 25316 44272 25344
rect 44223 25313 44235 25316
rect 44177 25307 44235 25313
rect 44266 25304 44272 25316
rect 44324 25304 44330 25356
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29104 25248 29561 25276
rect 28813 25239 28871 25245
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 31757 25279 31815 25285
rect 31757 25245 31769 25279
rect 31803 25276 31815 25279
rect 32122 25276 32128 25288
rect 31803 25248 32128 25276
rect 31803 25245 31815 25248
rect 31757 25239 31815 25245
rect 28736 25208 28764 25239
rect 32122 25236 32128 25248
rect 32180 25276 32186 25288
rect 32493 25279 32551 25285
rect 32493 25276 32505 25279
rect 32180 25248 32505 25276
rect 32180 25236 32186 25248
rect 32493 25245 32505 25248
rect 32539 25245 32551 25279
rect 32493 25239 32551 25245
rect 35986 25236 35992 25288
rect 36044 25236 36050 25288
rect 39574 25236 39580 25288
rect 39632 25236 39638 25288
rect 40037 25279 40095 25285
rect 40037 25245 40049 25279
rect 40083 25245 40095 25279
rect 40037 25239 40095 25245
rect 40129 25279 40187 25285
rect 40129 25245 40141 25279
rect 40175 25276 40187 25279
rect 40218 25276 40224 25288
rect 40175 25248 40224 25276
rect 40175 25245 40187 25248
rect 40129 25239 40187 25245
rect 28997 25211 29055 25217
rect 28997 25208 29009 25211
rect 28736 25180 29009 25208
rect 28997 25177 29009 25180
rect 29043 25208 29055 25211
rect 31665 25211 31723 25217
rect 31665 25208 31677 25211
rect 29043 25180 31677 25208
rect 29043 25177 29055 25180
rect 28997 25171 29055 25177
rect 31665 25177 31677 25180
rect 31711 25177 31723 25211
rect 36004 25208 36032 25236
rect 40052 25208 40080 25239
rect 40218 25236 40224 25248
rect 40276 25236 40282 25288
rect 40405 25279 40463 25285
rect 40405 25245 40417 25279
rect 40451 25276 40463 25279
rect 40586 25276 40592 25288
rect 40451 25248 40592 25276
rect 40451 25245 40463 25248
rect 40405 25239 40463 25245
rect 40586 25236 40592 25248
rect 40644 25236 40650 25288
rect 40681 25279 40739 25285
rect 40681 25245 40693 25279
rect 40727 25245 40739 25279
rect 40681 25239 40739 25245
rect 40696 25208 40724 25239
rect 40770 25236 40776 25288
rect 40828 25236 40834 25288
rect 41046 25236 41052 25288
rect 41104 25236 41110 25288
rect 41230 25236 41236 25288
rect 41288 25236 41294 25288
rect 41248 25208 41276 25236
rect 36004 25180 37122 25208
rect 40052 25180 41276 25208
rect 31665 25171 31723 25177
rect 43254 25168 43260 25220
rect 43312 25168 43318 25220
rect 27154 25140 27160 25152
rect 25924 25112 27160 25140
rect 25924 25100 25930 25112
rect 27154 25100 27160 25112
rect 27212 25100 27218 25152
rect 31938 25100 31944 25152
rect 31996 25100 32002 25152
rect 38010 25100 38016 25152
rect 38068 25140 38074 25152
rect 38105 25143 38163 25149
rect 38105 25140 38117 25143
rect 38068 25112 38117 25140
rect 38068 25100 38074 25112
rect 38105 25109 38117 25112
rect 38151 25109 38163 25143
rect 38105 25103 38163 25109
rect 42429 25143 42487 25149
rect 42429 25109 42441 25143
rect 42475 25140 42487 25143
rect 43070 25140 43076 25152
rect 42475 25112 43076 25140
rect 42475 25109 42487 25112
rect 42429 25103 42487 25109
rect 43070 25100 43076 25112
rect 43128 25100 43134 25152
rect 1104 25050 44620 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 44620 25050
rect 1104 24976 44620 24998
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 11885 24939 11943 24945
rect 11885 24936 11897 24939
rect 11756 24908 11897 24936
rect 11756 24896 11762 24908
rect 11885 24905 11897 24908
rect 11931 24905 11943 24939
rect 11885 24899 11943 24905
rect 15562 24896 15568 24948
rect 15620 24936 15626 24948
rect 16117 24939 16175 24945
rect 16117 24936 16129 24939
rect 15620 24908 16129 24936
rect 15620 24896 15626 24908
rect 16117 24905 16129 24908
rect 16163 24905 16175 24939
rect 16117 24899 16175 24905
rect 18414 24896 18420 24948
rect 18472 24896 18478 24948
rect 25682 24896 25688 24948
rect 25740 24896 25746 24948
rect 26142 24896 26148 24948
rect 26200 24936 26206 24948
rect 26200 24908 27476 24936
rect 26200 24896 26206 24908
rect 15654 24868 15660 24880
rect 15318 24840 15660 24868
rect 15654 24828 15660 24840
rect 15712 24868 15718 24880
rect 15712 24840 17434 24868
rect 15712 24828 15718 24840
rect 21634 24828 21640 24880
rect 21692 24868 21698 24880
rect 21692 24840 22508 24868
rect 21692 24828 21698 24840
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 11977 24803 12035 24809
rect 10735 24772 11560 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 11330 24692 11336 24744
rect 11388 24692 11394 24744
rect 10873 24667 10931 24673
rect 10873 24633 10885 24667
rect 10919 24664 10931 24667
rect 11348 24664 11376 24692
rect 11532 24673 11560 24772
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 12023 24772 13216 24800
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 12986 24732 12992 24744
rect 12207 24704 12992 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 13188 24732 13216 24772
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 16574 24760 16580 24812
rect 16632 24800 16638 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16632 24772 16681 24800
rect 16632 24760 16638 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19061 24803 19119 24809
rect 19061 24800 19073 24803
rect 19024 24772 19073 24800
rect 19024 24760 19030 24772
rect 19061 24769 19073 24772
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 13188 24704 13860 24732
rect 13832 24676 13860 24704
rect 14090 24692 14096 24744
rect 14148 24692 14154 24744
rect 16206 24692 16212 24744
rect 16264 24692 16270 24744
rect 16393 24735 16451 24741
rect 16393 24701 16405 24735
rect 16439 24732 16451 24735
rect 16439 24704 16528 24732
rect 16439 24701 16451 24704
rect 16393 24695 16451 24701
rect 10919 24636 11376 24664
rect 11517 24667 11575 24673
rect 10919 24633 10931 24636
rect 10873 24627 10931 24633
rect 11517 24633 11529 24667
rect 11563 24633 11575 24667
rect 11517 24627 11575 24633
rect 13814 24624 13820 24676
rect 13872 24624 13878 24676
rect 15746 24556 15752 24608
rect 15804 24556 15810 24608
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 16500 24596 16528 24704
rect 16942 24692 16948 24744
rect 17000 24692 17006 24744
rect 19168 24608 19196 24763
rect 22186 24760 22192 24812
rect 22244 24760 22250 24812
rect 22480 24809 22508 24840
rect 23474 24828 23480 24880
rect 23532 24828 23538 24880
rect 27062 24868 27068 24880
rect 26068 24840 27068 24868
rect 22465 24803 22523 24809
rect 22465 24769 22477 24803
rect 22511 24769 22523 24803
rect 22465 24763 22523 24769
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24800 25927 24803
rect 26068 24800 26096 24840
rect 26252 24812 26280 24840
rect 27062 24828 27068 24840
rect 27120 24828 27126 24880
rect 27448 24868 27476 24908
rect 27706 24896 27712 24948
rect 27764 24896 27770 24948
rect 32122 24896 32128 24948
rect 32180 24896 32186 24948
rect 40586 24896 40592 24948
rect 40644 24896 40650 24948
rect 44634 24896 44640 24948
rect 44692 24896 44698 24948
rect 31938 24868 31944 24880
rect 27172 24840 27384 24868
rect 27448 24840 27752 24868
rect 25915 24772 26096 24800
rect 25915 24769 25927 24772
rect 25869 24763 25927 24769
rect 26142 24760 26148 24812
rect 26200 24760 26206 24812
rect 26234 24760 26240 24812
rect 26292 24760 26298 24812
rect 26973 24803 27031 24809
rect 26973 24769 26985 24803
rect 27019 24800 27031 24803
rect 27172 24800 27200 24840
rect 27019 24772 27200 24800
rect 27249 24803 27307 24809
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 27249 24769 27261 24803
rect 27295 24769 27307 24803
rect 27356 24800 27384 24840
rect 27617 24803 27675 24809
rect 27617 24800 27629 24803
rect 27356 24772 27629 24800
rect 27249 24763 27307 24769
rect 27617 24769 27629 24772
rect 27663 24769 27675 24803
rect 27724 24800 27752 24840
rect 31680 24840 31944 24868
rect 27798 24800 27804 24812
rect 27724 24772 27804 24800
rect 27617 24763 27675 24769
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22388 24704 22753 24732
rect 22388 24673 22416 24704
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 26988 24732 27016 24763
rect 22741 24695 22799 24701
rect 26068 24704 27016 24732
rect 26068 24676 26096 24704
rect 27154 24692 27160 24744
rect 27212 24692 27218 24744
rect 22373 24667 22431 24673
rect 22373 24633 22385 24667
rect 22419 24633 22431 24667
rect 22373 24627 22431 24633
rect 23750 24624 23756 24676
rect 23808 24664 23814 24676
rect 25866 24664 25872 24676
rect 23808 24636 25872 24664
rect 23808 24624 23814 24636
rect 25866 24624 25872 24636
rect 25924 24664 25930 24676
rect 25961 24667 26019 24673
rect 25961 24664 25973 24667
rect 25924 24636 25973 24664
rect 25924 24624 25930 24636
rect 25961 24633 25973 24636
rect 26007 24633 26019 24667
rect 25961 24627 26019 24633
rect 26050 24624 26056 24676
rect 26108 24624 26114 24676
rect 27264 24664 27292 24763
rect 27798 24760 27804 24772
rect 27856 24760 27862 24812
rect 31386 24760 31392 24812
rect 31444 24760 31450 24812
rect 31570 24760 31576 24812
rect 31628 24760 31634 24812
rect 31680 24809 31708 24840
rect 31938 24828 31944 24840
rect 31996 24828 32002 24880
rect 32582 24828 32588 24880
rect 32640 24828 32646 24880
rect 39393 24871 39451 24877
rect 36556 24840 36860 24868
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24769 31723 24803
rect 31665 24763 31723 24769
rect 31757 24803 31815 24809
rect 31757 24769 31769 24803
rect 31803 24800 31815 24803
rect 32030 24800 32036 24812
rect 31803 24772 32036 24800
rect 31803 24769 31815 24772
rect 31757 24763 31815 24769
rect 32030 24760 32036 24772
rect 32088 24800 32094 24812
rect 32306 24800 32312 24812
rect 32088 24772 32312 24800
rect 32088 24760 32094 24772
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 33873 24803 33931 24809
rect 33873 24769 33885 24803
rect 33919 24800 33931 24803
rect 35710 24800 35716 24812
rect 33919 24772 35716 24800
rect 33919 24769 33931 24772
rect 33873 24763 33931 24769
rect 35710 24760 35716 24772
rect 35768 24760 35774 24812
rect 36173 24803 36231 24809
rect 36173 24769 36185 24803
rect 36219 24800 36231 24803
rect 36556 24800 36584 24840
rect 36725 24803 36783 24809
rect 36725 24800 36737 24803
rect 36219 24772 36584 24800
rect 36648 24772 36737 24800
rect 36219 24769 36231 24772
rect 36173 24763 36231 24769
rect 36648 24741 36676 24772
rect 36725 24769 36737 24772
rect 36771 24769 36783 24803
rect 36832 24800 36860 24840
rect 39393 24837 39405 24871
rect 39439 24868 39451 24871
rect 40126 24868 40132 24880
rect 39439 24840 40132 24868
rect 39439 24837 39451 24840
rect 39393 24831 39451 24837
rect 40126 24828 40132 24840
rect 40184 24828 40190 24880
rect 36998 24800 37004 24812
rect 36832 24772 37004 24800
rect 36725 24763 36783 24769
rect 36998 24760 37004 24772
rect 37056 24760 37062 24812
rect 39485 24803 39543 24809
rect 39485 24769 39497 24803
rect 39531 24800 39543 24803
rect 40604 24800 40632 24896
rect 39531 24772 40632 24800
rect 44269 24803 44327 24809
rect 39531 24769 39543 24772
rect 39485 24763 39543 24769
rect 44269 24769 44281 24803
rect 44315 24800 44327 24803
rect 44652 24800 44680 24896
rect 44315 24772 44680 24800
rect 44315 24769 44327 24772
rect 44269 24763 44327 24769
rect 33597 24735 33655 24741
rect 33597 24732 33609 24735
rect 31956 24704 33609 24732
rect 26896 24636 27292 24664
rect 27433 24667 27491 24673
rect 17678 24596 17684 24608
rect 15896 24568 17684 24596
rect 15896 24556 15902 24568
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 19150 24556 19156 24608
rect 19208 24556 19214 24608
rect 19242 24556 19248 24608
rect 19300 24596 19306 24608
rect 22002 24596 22008 24608
rect 19300 24568 22008 24596
rect 19300 24556 19306 24568
rect 22002 24556 22008 24568
rect 22060 24596 22066 24608
rect 24213 24599 24271 24605
rect 24213 24596 24225 24599
rect 22060 24568 24225 24596
rect 22060 24556 22066 24568
rect 24213 24565 24225 24568
rect 24259 24596 24271 24599
rect 25130 24596 25136 24608
rect 24259 24568 25136 24596
rect 24259 24565 24271 24568
rect 24213 24559 24271 24565
rect 25130 24556 25136 24568
rect 25188 24596 25194 24608
rect 26896 24596 26924 24636
rect 27433 24633 27445 24667
rect 27479 24664 27491 24667
rect 27522 24664 27528 24676
rect 27479 24636 27528 24664
rect 27479 24633 27491 24636
rect 27433 24627 27491 24633
rect 27522 24624 27528 24636
rect 27580 24624 27586 24676
rect 31956 24673 31984 24704
rect 33597 24701 33609 24704
rect 33643 24701 33655 24735
rect 33597 24695 33655 24701
rect 36633 24735 36691 24741
rect 36633 24701 36645 24735
rect 36679 24701 36691 24735
rect 36633 24695 36691 24701
rect 39298 24692 39304 24744
rect 39356 24732 39362 24744
rect 39577 24735 39635 24741
rect 39577 24732 39589 24735
rect 39356 24704 39589 24732
rect 39356 24692 39362 24704
rect 39577 24701 39589 24704
rect 39623 24701 39635 24735
rect 39577 24695 39635 24701
rect 31941 24667 31999 24673
rect 31941 24633 31953 24667
rect 31987 24633 31999 24667
rect 31941 24627 31999 24633
rect 36541 24667 36599 24673
rect 36541 24633 36553 24667
rect 36587 24664 36599 24667
rect 44085 24667 44143 24673
rect 44085 24664 44097 24667
rect 36587 24636 44097 24664
rect 36587 24633 36599 24636
rect 36541 24627 36599 24633
rect 44085 24633 44097 24636
rect 44131 24633 44143 24667
rect 44085 24627 44143 24633
rect 25188 24568 26924 24596
rect 25188 24556 25194 24568
rect 27062 24556 27068 24608
rect 27120 24556 27126 24608
rect 28534 24556 28540 24608
rect 28592 24596 28598 24608
rect 34422 24596 34428 24608
rect 28592 24568 34428 24596
rect 28592 24556 28598 24568
rect 34422 24556 34428 24568
rect 34480 24556 34486 24608
rect 36906 24556 36912 24608
rect 36964 24556 36970 24608
rect 39022 24556 39028 24608
rect 39080 24556 39086 24608
rect 1104 24506 44620 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 44620 24506
rect 1104 24432 44620 24454
rect 12894 24352 12900 24404
rect 12952 24392 12958 24404
rect 13357 24395 13415 24401
rect 13357 24392 13369 24395
rect 12952 24364 13369 24392
rect 12952 24352 12958 24364
rect 13357 24361 13369 24364
rect 13403 24361 13415 24395
rect 13357 24355 13415 24361
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 14461 24395 14519 24401
rect 14461 24392 14473 24395
rect 14148 24364 14473 24392
rect 14148 24352 14154 24364
rect 14461 24361 14473 24364
rect 14507 24361 14519 24395
rect 14461 24355 14519 24361
rect 15746 24352 15752 24404
rect 15804 24352 15810 24404
rect 16853 24395 16911 24401
rect 16853 24361 16865 24395
rect 16899 24392 16911 24395
rect 16942 24392 16948 24404
rect 16899 24364 16948 24392
rect 16899 24361 16911 24364
rect 16853 24355 16911 24361
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22186 24392 22192 24404
rect 22143 24364 22192 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 31113 24395 31171 24401
rect 31113 24361 31125 24395
rect 31159 24392 31171 24395
rect 31386 24392 31392 24404
rect 31159 24364 31392 24392
rect 31159 24361 31171 24364
rect 31113 24355 31171 24361
rect 31386 24352 31392 24364
rect 31444 24352 31450 24404
rect 39390 24392 39396 24404
rect 31726 24364 39396 24392
rect 13078 24284 13084 24336
rect 13136 24324 13142 24336
rect 14185 24327 14243 24333
rect 14185 24324 14197 24327
rect 13136 24296 14197 24324
rect 13136 24284 13142 24296
rect 14185 24293 14197 24296
rect 14231 24293 14243 24327
rect 14185 24287 14243 24293
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11609 24259 11667 24265
rect 11609 24256 11621 24259
rect 11112 24228 11621 24256
rect 11112 24216 11118 24228
rect 11609 24225 11621 24228
rect 11655 24225 11667 24259
rect 15764 24256 15792 24352
rect 19061 24327 19119 24333
rect 19061 24293 19073 24327
rect 19107 24324 19119 24327
rect 19150 24324 19156 24336
rect 19107 24296 19156 24324
rect 19107 24293 19119 24296
rect 19061 24287 19119 24293
rect 19150 24284 19156 24296
rect 19208 24324 19214 24336
rect 19208 24296 20668 24324
rect 19208 24284 19214 24296
rect 11609 24219 11667 24225
rect 14660 24228 15792 24256
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 14550 24188 14556 24200
rect 14323 24160 14556 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 14660 24197 14688 24228
rect 16574 24216 16580 24268
rect 16632 24256 16638 24268
rect 17313 24259 17371 24265
rect 17313 24256 17325 24259
rect 16632 24228 17325 24256
rect 16632 24216 16638 24228
rect 17313 24225 17325 24228
rect 17359 24225 17371 24259
rect 17313 24219 17371 24225
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24256 19855 24259
rect 19978 24256 19984 24268
rect 19843 24228 19984 24256
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20640 24265 20668 24296
rect 20732 24296 28994 24324
rect 20625 24259 20683 24265
rect 20625 24225 20637 24259
rect 20671 24225 20683 24259
rect 20625 24219 20683 24225
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24157 14703 24191
rect 14645 24151 14703 24157
rect 14734 24148 14740 24200
rect 14792 24188 14798 24200
rect 14829 24191 14887 24197
rect 14829 24188 14841 24191
rect 14792 24160 14841 24188
rect 14792 24148 14798 24160
rect 14829 24157 14841 24160
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24188 16727 24191
rect 17126 24188 17132 24200
rect 16715 24160 17132 24188
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 20732 24188 20760 24296
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 23566 24256 23572 24268
rect 22704 24228 23572 24256
rect 22704 24216 22710 24228
rect 23566 24216 23572 24228
rect 23624 24216 23630 24268
rect 28966 24256 28994 24296
rect 29546 24284 29552 24336
rect 29604 24284 29610 24336
rect 31726 24324 31754 24364
rect 39390 24352 39396 24364
rect 39448 24352 39454 24404
rect 42889 24395 42947 24401
rect 42889 24361 42901 24395
rect 42935 24392 42947 24395
rect 42978 24392 42984 24404
rect 42935 24364 42984 24392
rect 42935 24361 42947 24364
rect 42889 24355 42947 24361
rect 42978 24352 42984 24364
rect 43036 24352 43042 24404
rect 29656 24296 31754 24324
rect 29656 24256 29684 24296
rect 39022 24284 39028 24336
rect 39080 24284 39086 24336
rect 28966 24228 29684 24256
rect 30193 24259 30251 24265
rect 30193 24225 30205 24259
rect 30239 24256 30251 24259
rect 30745 24259 30803 24265
rect 30745 24256 30757 24259
rect 30239 24228 30757 24256
rect 30239 24225 30251 24228
rect 30193 24219 30251 24225
rect 30745 24225 30757 24228
rect 30791 24225 30803 24259
rect 30745 24219 30803 24225
rect 32674 24216 32680 24268
rect 32732 24256 32738 24268
rect 32769 24259 32827 24265
rect 32769 24256 32781 24259
rect 32732 24228 32781 24256
rect 32732 24216 32738 24228
rect 32769 24225 32781 24228
rect 32815 24225 32827 24259
rect 32769 24219 32827 24225
rect 34514 24216 34520 24268
rect 34572 24256 34578 24268
rect 35253 24259 35311 24265
rect 35253 24256 35265 24259
rect 34572 24228 35265 24256
rect 34572 24216 34578 24228
rect 35253 24225 35265 24228
rect 35299 24225 35311 24259
rect 35253 24219 35311 24225
rect 18892 24160 20760 24188
rect 11882 24080 11888 24132
rect 11940 24080 11946 24132
rect 12434 24080 12440 24132
rect 12492 24080 12498 24132
rect 13188 24092 15424 24120
rect 12618 24012 12624 24064
rect 12676 24052 12682 24064
rect 13188 24052 13216 24092
rect 12676 24024 13216 24052
rect 15013 24055 15071 24061
rect 12676 24012 12682 24024
rect 15013 24021 15025 24055
rect 15059 24052 15071 24055
rect 15286 24052 15292 24064
rect 15059 24024 15292 24052
rect 15059 24021 15071 24024
rect 15013 24015 15071 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 15396 24052 15424 24092
rect 17586 24080 17592 24132
rect 17644 24080 17650 24132
rect 18046 24080 18052 24132
rect 18104 24080 18110 24132
rect 18892 24052 18920 24160
rect 20990 24148 20996 24200
rect 21048 24148 21054 24200
rect 22002 24148 22008 24200
rect 22060 24188 22066 24200
rect 22465 24191 22523 24197
rect 22465 24188 22477 24191
rect 22060 24160 22477 24188
rect 22060 24148 22066 24160
rect 22465 24157 22477 24160
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 24578 24148 24584 24200
rect 24636 24188 24642 24200
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 24636 24160 24961 24188
rect 24636 24148 24642 24160
rect 24949 24157 24961 24160
rect 24995 24157 25007 24191
rect 24949 24151 25007 24157
rect 29549 24191 29607 24197
rect 29549 24157 29561 24191
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 29825 24191 29883 24197
rect 29825 24157 29837 24191
rect 29871 24188 29883 24191
rect 29914 24188 29920 24200
rect 29871 24160 29920 24188
rect 29871 24157 29883 24160
rect 29825 24151 29883 24157
rect 19613 24123 19671 24129
rect 19613 24089 19625 24123
rect 19659 24120 19671 24123
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19659 24092 20085 24120
rect 19659 24089 19671 24092
rect 19613 24083 19671 24089
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 22186 24120 22192 24132
rect 20073 24083 20131 24089
rect 20732 24092 22192 24120
rect 15396 24024 18920 24052
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19705 24055 19763 24061
rect 19705 24021 19717 24055
rect 19751 24052 19763 24055
rect 20732 24052 20760 24092
rect 22186 24080 22192 24092
rect 22244 24080 22250 24132
rect 29564 24120 29592 24151
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 30006 24148 30012 24200
rect 30064 24148 30070 24200
rect 30098 24148 30104 24200
rect 30156 24148 30162 24200
rect 30282 24148 30288 24200
rect 30340 24148 30346 24200
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 30432 24160 30696 24188
rect 30432 24148 30438 24160
rect 30024 24120 30052 24148
rect 29564 24092 30052 24120
rect 30668 24064 30696 24160
rect 30834 24148 30840 24200
rect 30892 24148 30898 24200
rect 36354 24148 36360 24200
rect 36412 24188 36418 24200
rect 36909 24191 36967 24197
rect 36909 24188 36921 24191
rect 36412 24160 36921 24188
rect 36412 24148 36418 24160
rect 36909 24157 36921 24160
rect 36955 24157 36967 24191
rect 36909 24151 36967 24157
rect 37550 24148 37556 24200
rect 37608 24148 37614 24200
rect 38841 24191 38899 24197
rect 38841 24157 38853 24191
rect 38887 24188 38899 24191
rect 39040 24188 39068 24284
rect 40034 24216 40040 24268
rect 40092 24256 40098 24268
rect 40497 24259 40555 24265
rect 40497 24256 40509 24259
rect 40092 24228 40509 24256
rect 40092 24216 40098 24228
rect 40497 24225 40509 24228
rect 40543 24225 40555 24259
rect 40497 24219 40555 24225
rect 43073 24259 43131 24265
rect 43073 24225 43085 24259
rect 43119 24256 43131 24259
rect 43530 24256 43536 24268
rect 43119 24228 43536 24256
rect 43119 24225 43131 24228
rect 43073 24219 43131 24225
rect 43530 24216 43536 24228
rect 43588 24216 43594 24268
rect 38887 24160 39068 24188
rect 38887 24157 38899 24160
rect 38841 24151 38899 24157
rect 40218 24148 40224 24200
rect 40276 24148 40282 24200
rect 42797 24191 42855 24197
rect 42797 24157 42809 24191
rect 42843 24188 42855 24191
rect 43346 24188 43352 24200
rect 42843 24160 43352 24188
rect 42843 24157 42855 24160
rect 42797 24151 42855 24157
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 33042 24080 33048 24132
rect 33100 24080 33106 24132
rect 34790 24120 34796 24132
rect 34270 24092 34796 24120
rect 34790 24080 34796 24092
rect 34848 24080 34854 24132
rect 40773 24123 40831 24129
rect 40773 24120 40785 24123
rect 40420 24092 40785 24120
rect 19751 24024 20760 24052
rect 19751 24021 19763 24024
rect 19705 24015 19763 24021
rect 20806 24012 20812 24064
rect 20864 24012 20870 24064
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 22094 24052 22100 24064
rect 21140 24024 22100 24052
rect 21140 24012 21146 24024
rect 22094 24012 22100 24024
rect 22152 24012 22158 24064
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 22557 24055 22615 24061
rect 22557 24052 22569 24055
rect 22336 24024 22569 24052
rect 22336 24012 22342 24024
rect 22557 24021 22569 24024
rect 22603 24021 22615 24055
rect 22557 24015 22615 24021
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 24302 24052 24308 24064
rect 23532 24024 24308 24052
rect 23532 24012 23538 24024
rect 24302 24012 24308 24024
rect 24360 24052 24366 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 24360 24024 24409 24052
rect 24360 24012 24366 24024
rect 24397 24021 24409 24024
rect 24443 24021 24455 24055
rect 24397 24015 24455 24021
rect 29178 24012 29184 24064
rect 29236 24052 29242 24064
rect 29733 24055 29791 24061
rect 29733 24052 29745 24055
rect 29236 24024 29745 24052
rect 29236 24012 29242 24024
rect 29733 24021 29745 24024
rect 29779 24052 29791 24055
rect 30098 24052 30104 24064
rect 29779 24024 30104 24052
rect 29779 24021 29791 24024
rect 29733 24015 29791 24021
rect 30098 24012 30104 24024
rect 30156 24012 30162 24064
rect 30466 24012 30472 24064
rect 30524 24012 30530 24064
rect 30650 24012 30656 24064
rect 30708 24012 30714 24064
rect 34698 24012 34704 24064
rect 34756 24012 34762 24064
rect 35802 24012 35808 24064
rect 35860 24052 35866 24064
rect 37093 24055 37151 24061
rect 37093 24052 37105 24055
rect 35860 24024 37105 24052
rect 35860 24012 35866 24024
rect 37093 24021 37105 24024
rect 37139 24052 37151 24055
rect 37274 24052 37280 24064
rect 37139 24024 37280 24052
rect 37139 24021 37151 24024
rect 37093 24015 37151 24021
rect 37274 24012 37280 24024
rect 37332 24012 37338 24064
rect 37366 24012 37372 24064
rect 37424 24012 37430 24064
rect 39025 24055 39083 24061
rect 39025 24021 39037 24055
rect 39071 24052 39083 24055
rect 39206 24052 39212 24064
rect 39071 24024 39212 24052
rect 39071 24021 39083 24024
rect 39025 24015 39083 24021
rect 39206 24012 39212 24024
rect 39264 24012 39270 24064
rect 40420 24061 40448 24092
rect 40773 24089 40785 24092
rect 40819 24089 40831 24123
rect 40773 24083 40831 24089
rect 41156 24092 41262 24120
rect 41156 24064 41184 24092
rect 40405 24055 40463 24061
rect 40405 24021 40417 24055
rect 40451 24021 40463 24055
rect 40405 24015 40463 24021
rect 41138 24012 41144 24064
rect 41196 24012 41202 24064
rect 42242 24012 42248 24064
rect 42300 24012 42306 24064
rect 43073 24055 43131 24061
rect 43073 24021 43085 24055
rect 43119 24052 43131 24055
rect 43162 24052 43168 24064
rect 43119 24024 43168 24052
rect 43119 24021 43131 24024
rect 43073 24015 43131 24021
rect 43162 24012 43168 24024
rect 43220 24012 43226 24064
rect 1104 23962 44620 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 44620 23962
rect 1104 23888 44620 23910
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 12069 23851 12127 23857
rect 12069 23848 12081 23851
rect 11940 23820 12081 23848
rect 11940 23808 11946 23820
rect 12069 23817 12081 23820
rect 12115 23817 12127 23851
rect 12069 23811 12127 23817
rect 12345 23851 12403 23857
rect 12345 23817 12357 23851
rect 12391 23817 12403 23851
rect 12345 23811 12403 23817
rect 12713 23851 12771 23857
rect 12713 23817 12725 23851
rect 12759 23848 12771 23851
rect 12894 23848 12900 23860
rect 12759 23820 12900 23848
rect 12759 23817 12771 23820
rect 12713 23811 12771 23817
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 12360 23712 12388 23811
rect 12894 23808 12900 23820
rect 12952 23808 12958 23860
rect 14550 23808 14556 23860
rect 14608 23848 14614 23860
rect 15289 23851 15347 23857
rect 15289 23848 15301 23851
rect 14608 23820 15301 23848
rect 14608 23808 14614 23820
rect 15289 23817 15301 23820
rect 15335 23817 15347 23851
rect 15289 23811 15347 23817
rect 15102 23780 15108 23792
rect 15042 23752 15108 23780
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 12299 23684 12388 23712
rect 15304 23712 15332 23811
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 18141 23851 18199 23857
rect 18141 23848 18153 23851
rect 17644 23820 18153 23848
rect 17644 23808 17650 23820
rect 18141 23817 18153 23820
rect 18187 23817 18199 23851
rect 18141 23811 18199 23817
rect 19242 23808 19248 23860
rect 19300 23808 19306 23860
rect 20806 23848 20812 23860
rect 20180 23820 20812 23848
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15304 23684 15945 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 18325 23715 18383 23721
rect 18325 23681 18337 23715
rect 18371 23712 18383 23715
rect 19260 23712 19288 23808
rect 20180 23789 20208 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 25038 23808 25044 23860
rect 25096 23848 25102 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 25096 23820 25145 23848
rect 25096 23808 25102 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25133 23811 25191 23817
rect 29546 23808 29552 23860
rect 29604 23808 29610 23860
rect 30466 23808 30472 23860
rect 30524 23808 30530 23860
rect 30834 23808 30840 23860
rect 30892 23848 30898 23860
rect 31389 23851 31447 23857
rect 31389 23848 31401 23851
rect 30892 23820 31401 23848
rect 30892 23808 30898 23820
rect 31389 23817 31401 23820
rect 31435 23817 31447 23851
rect 31389 23811 31447 23817
rect 33042 23808 33048 23860
rect 33100 23848 33106 23860
rect 33689 23851 33747 23857
rect 33689 23848 33701 23851
rect 33100 23820 33701 23848
rect 33100 23808 33106 23820
rect 33689 23817 33701 23820
rect 33735 23817 33747 23851
rect 34425 23851 34483 23857
rect 34425 23848 34437 23851
rect 33689 23811 33747 23817
rect 33888 23820 34437 23848
rect 20165 23783 20223 23789
rect 20165 23749 20177 23783
rect 20211 23749 20223 23783
rect 20165 23743 20223 23749
rect 20898 23740 20904 23792
rect 20956 23740 20962 23792
rect 18371 23684 19288 23712
rect 23124 23684 26372 23712
rect 18371 23681 18383 23684
rect 18325 23675 18383 23681
rect 12805 23647 12863 23653
rect 12805 23613 12817 23647
rect 12851 23613 12863 23647
rect 12805 23607 12863 23613
rect 12820 23576 12848 23607
rect 12986 23604 12992 23656
rect 13044 23604 13050 23656
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 13814 23604 13820 23656
rect 13872 23604 13878 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 19889 23647 19947 23653
rect 19889 23644 19901 23647
rect 19392 23616 19901 23644
rect 19392 23604 19398 23616
rect 19889 23613 19901 23616
rect 19935 23613 19947 23647
rect 23124 23644 23152 23684
rect 19889 23607 19947 23613
rect 19996 23616 23152 23644
rect 12820 23548 12940 23576
rect 12912 23508 12940 23548
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 19996 23576 20024 23616
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 26234 23576 26240 23588
rect 19484 23548 20024 23576
rect 21192 23548 26240 23576
rect 19484 23536 19490 23548
rect 14458 23508 14464 23520
rect 12912 23480 14464 23508
rect 14458 23468 14464 23480
rect 14516 23468 14522 23520
rect 15378 23468 15384 23520
rect 15436 23468 15442 23520
rect 16206 23468 16212 23520
rect 16264 23508 16270 23520
rect 21192 23508 21220 23548
rect 26234 23536 26240 23548
rect 26292 23536 26298 23588
rect 26344 23576 26372 23684
rect 26418 23672 26424 23724
rect 26476 23672 26482 23724
rect 29564 23721 29592 23808
rect 29730 23740 29736 23792
rect 29788 23740 29794 23792
rect 30484 23780 30512 23808
rect 30484 23752 31616 23780
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 29914 23672 29920 23724
rect 29972 23672 29978 23724
rect 30098 23672 30104 23724
rect 30156 23672 30162 23724
rect 30466 23672 30472 23724
rect 30524 23672 30530 23724
rect 31036 23721 31064 23752
rect 31588 23721 31616 23752
rect 33888 23721 33916 23820
rect 34425 23817 34437 23820
rect 34471 23817 34483 23851
rect 34425 23811 34483 23817
rect 34698 23808 34704 23860
rect 34756 23808 34762 23860
rect 35434 23808 35440 23860
rect 35492 23808 35498 23860
rect 36906 23848 36912 23860
rect 36832 23820 36912 23848
rect 34716 23780 34744 23808
rect 34348 23752 34744 23780
rect 34793 23783 34851 23789
rect 30653 23715 30711 23721
rect 30653 23681 30665 23715
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 31021 23715 31079 23721
rect 31021 23681 31033 23715
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 31389 23715 31447 23721
rect 31389 23681 31401 23715
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23681 31631 23715
rect 31573 23675 31631 23681
rect 33873 23715 33931 23721
rect 33873 23681 33885 23715
rect 33919 23681 33931 23715
rect 33873 23675 33931 23681
rect 33965 23715 34023 23721
rect 33965 23681 33977 23715
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 29932 23644 29960 23672
rect 30668 23644 30696 23675
rect 31404 23644 31432 23675
rect 29932 23616 31432 23644
rect 32490 23576 32496 23588
rect 26344 23548 32496 23576
rect 32490 23536 32496 23548
rect 32548 23536 32554 23588
rect 33980 23576 34008 23675
rect 34054 23672 34060 23724
rect 34112 23672 34118 23724
rect 34146 23672 34152 23724
rect 34204 23721 34210 23724
rect 34348 23721 34376 23752
rect 34793 23749 34805 23783
rect 34839 23780 34851 23783
rect 34839 23752 35112 23780
rect 34839 23749 34851 23752
rect 34793 23743 34851 23749
rect 34204 23715 34233 23721
rect 34221 23681 34233 23715
rect 34204 23675 34233 23681
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23681 34391 23715
rect 34333 23675 34391 23681
rect 34204 23672 34210 23675
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 35084 23721 35112 23752
rect 34885 23715 34943 23721
rect 34885 23712 34897 23715
rect 34664 23684 34897 23712
rect 34664 23672 34670 23684
rect 34885 23681 34897 23684
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 35069 23715 35127 23721
rect 35069 23681 35081 23715
rect 35115 23712 35127 23715
rect 35452 23712 35480 23808
rect 35802 23740 35808 23792
rect 35860 23740 35866 23792
rect 36832 23789 36860 23820
rect 36906 23808 36912 23820
rect 36964 23808 36970 23860
rect 39206 23808 39212 23860
rect 39264 23848 39270 23860
rect 39264 23820 39436 23848
rect 39264 23808 39270 23820
rect 36817 23783 36875 23789
rect 36817 23749 36829 23783
rect 36863 23749 36875 23783
rect 36817 23743 36875 23749
rect 38654 23740 38660 23792
rect 38712 23780 38718 23792
rect 39408 23789 39436 23820
rect 40218 23808 40224 23860
rect 40276 23848 40282 23860
rect 40957 23851 41015 23857
rect 40957 23848 40969 23851
rect 40276 23820 40969 23848
rect 40276 23808 40282 23820
rect 40957 23817 40969 23820
rect 41003 23817 41015 23851
rect 40957 23811 41015 23817
rect 41046 23808 41052 23860
rect 41104 23848 41110 23860
rect 41417 23851 41475 23857
rect 41417 23848 41429 23851
rect 41104 23820 41429 23848
rect 41104 23808 41110 23820
rect 41417 23817 41429 23820
rect 41463 23817 41475 23851
rect 41417 23811 41475 23817
rect 42242 23808 42248 23860
rect 42300 23808 42306 23860
rect 42794 23808 42800 23860
rect 42852 23848 42858 23860
rect 42852 23820 43484 23848
rect 42852 23808 42858 23820
rect 39025 23783 39083 23789
rect 39025 23780 39037 23783
rect 38712 23752 39037 23780
rect 38712 23740 38718 23752
rect 39025 23749 39037 23752
rect 39071 23749 39083 23783
rect 39025 23743 39083 23749
rect 39393 23783 39451 23789
rect 39393 23749 39405 23783
rect 39439 23749 39451 23783
rect 41138 23780 41144 23792
rect 40618 23752 41144 23780
rect 39393 23743 39451 23749
rect 41138 23740 41144 23752
rect 41196 23740 41202 23792
rect 41325 23783 41383 23789
rect 41325 23749 41337 23783
rect 41371 23780 41383 23783
rect 41506 23780 41512 23792
rect 41371 23752 41512 23780
rect 41371 23749 41383 23752
rect 41325 23743 41383 23749
rect 41506 23740 41512 23752
rect 41564 23780 41570 23792
rect 42260 23780 42288 23808
rect 42886 23780 42892 23792
rect 41564 23752 42288 23780
rect 42720 23752 42892 23780
rect 41564 23740 41570 23752
rect 35115 23684 35480 23712
rect 35115 23681 35127 23684
rect 35069 23675 35127 23681
rect 37090 23604 37096 23656
rect 37148 23644 37154 23656
rect 39117 23647 39175 23653
rect 39117 23644 39129 23647
rect 37148 23616 39129 23644
rect 37148 23604 37154 23616
rect 34698 23576 34704 23588
rect 33980 23548 34704 23576
rect 34698 23536 34704 23548
rect 34756 23576 34762 23588
rect 37752 23585 37780 23616
rect 39117 23613 39129 23616
rect 39163 23613 39175 23647
rect 39117 23607 39175 23613
rect 39390 23604 39396 23656
rect 39448 23644 39454 23656
rect 41509 23647 41567 23653
rect 41509 23644 41521 23647
rect 39448 23616 41521 23644
rect 39448 23604 39454 23616
rect 41509 23613 41521 23616
rect 41555 23644 41567 23647
rect 42720 23644 42748 23752
rect 42886 23740 42892 23752
rect 42944 23740 42950 23792
rect 43346 23780 43352 23792
rect 43272 23752 43352 23780
rect 42797 23715 42855 23721
rect 42797 23681 42809 23715
rect 42843 23681 42855 23715
rect 42797 23675 42855 23681
rect 41555 23616 42748 23644
rect 41555 23613 41567 23616
rect 41509 23607 41567 23613
rect 34977 23579 35035 23585
rect 34977 23576 34989 23579
rect 34756 23548 34989 23576
rect 34756 23536 34762 23548
rect 34977 23545 34989 23548
rect 35023 23545 35035 23579
rect 34977 23539 35035 23545
rect 37737 23579 37795 23585
rect 37737 23545 37749 23579
rect 37783 23545 37795 23579
rect 42812 23576 42840 23675
rect 42978 23672 42984 23724
rect 43036 23712 43042 23724
rect 43272 23721 43300 23752
rect 43346 23740 43352 23752
rect 43404 23740 43410 23792
rect 43456 23721 43484 23820
rect 43257 23715 43315 23721
rect 43036 23684 43208 23712
rect 43036 23672 43042 23684
rect 42889 23647 42947 23653
rect 42889 23613 42901 23647
rect 42935 23644 42947 23647
rect 43073 23647 43131 23653
rect 43073 23644 43085 23647
rect 42935 23616 43085 23644
rect 42935 23613 42947 23616
rect 42889 23607 42947 23613
rect 43073 23613 43085 23616
rect 43119 23613 43131 23647
rect 43180 23644 43208 23684
rect 43257 23681 43269 23715
rect 43303 23681 43315 23715
rect 43257 23675 43315 23681
rect 43441 23715 43499 23721
rect 43441 23681 43453 23715
rect 43487 23681 43499 23715
rect 43441 23675 43499 23681
rect 43530 23672 43536 23724
rect 43588 23672 43594 23724
rect 43346 23644 43352 23656
rect 43180 23616 43352 23644
rect 43073 23607 43131 23613
rect 43346 23604 43352 23616
rect 43404 23604 43410 23656
rect 42812 23548 43116 23576
rect 37737 23539 37795 23545
rect 43088 23520 43116 23548
rect 16264 23480 21220 23508
rect 16264 23468 16270 23480
rect 21542 23468 21548 23520
rect 21600 23508 21606 23520
rect 21637 23511 21695 23517
rect 21637 23508 21649 23511
rect 21600 23480 21649 23508
rect 21600 23468 21606 23480
rect 21637 23477 21649 23480
rect 21683 23477 21695 23511
rect 21637 23471 21695 23477
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 22649 23511 22707 23517
rect 22649 23508 22661 23511
rect 22336 23480 22661 23508
rect 22336 23468 22342 23480
rect 22649 23477 22661 23480
rect 22695 23477 22707 23511
rect 22649 23471 22707 23477
rect 29638 23468 29644 23520
rect 29696 23508 29702 23520
rect 30282 23508 30288 23520
rect 29696 23480 30288 23508
rect 29696 23468 29702 23480
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 35345 23511 35403 23517
rect 35345 23477 35357 23511
rect 35391 23508 35403 23511
rect 35618 23508 35624 23520
rect 35391 23480 35624 23508
rect 35391 23477 35403 23480
rect 35345 23471 35403 23477
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 40126 23468 40132 23520
rect 40184 23508 40190 23520
rect 40865 23511 40923 23517
rect 40865 23508 40877 23511
rect 40184 23480 40877 23508
rect 40184 23468 40190 23480
rect 40865 23477 40877 23480
rect 40911 23477 40923 23511
rect 40865 23471 40923 23477
rect 42426 23468 42432 23520
rect 42484 23468 42490 23520
rect 43070 23468 43076 23520
rect 43128 23468 43134 23520
rect 1104 23418 44620 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 44620 23418
rect 1104 23344 44620 23366
rect 13814 23264 13820 23316
rect 13872 23304 13878 23316
rect 14093 23307 14151 23313
rect 14093 23304 14105 23307
rect 13872 23276 14105 23304
rect 13872 23264 13878 23276
rect 14093 23273 14105 23276
rect 14139 23273 14151 23307
rect 14093 23267 14151 23273
rect 14366 23264 14372 23316
rect 14424 23304 14430 23316
rect 15102 23304 15108 23316
rect 14424 23276 15108 23304
rect 14424 23264 14430 23276
rect 15102 23264 15108 23276
rect 15160 23304 15166 23316
rect 15565 23307 15623 23313
rect 15565 23304 15577 23307
rect 15160 23276 15577 23304
rect 15160 23264 15166 23276
rect 15565 23273 15577 23276
rect 15611 23304 15623 23307
rect 17402 23304 17408 23316
rect 15611 23276 17408 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 17494 23264 17500 23316
rect 17552 23304 17558 23316
rect 17552 23276 20852 23304
rect 17552 23264 17558 23276
rect 14553 23239 14611 23245
rect 14553 23205 14565 23239
rect 14599 23205 14611 23239
rect 14553 23199 14611 23205
rect 15028 23208 19334 23236
rect 11609 23171 11667 23177
rect 11609 23137 11621 23171
rect 11655 23168 11667 23171
rect 12986 23168 12992 23180
rect 11655 23140 12992 23168
rect 11655 23137 11667 23140
rect 11609 23131 11667 23137
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23100 10839 23103
rect 11333 23103 11391 23109
rect 10827 23072 11008 23100
rect 10827 23069 10839 23072
rect 10781 23063 10839 23069
rect 10042 22924 10048 22976
rect 10100 22964 10106 22976
rect 10321 22967 10379 22973
rect 10321 22964 10333 22967
rect 10100 22936 10333 22964
rect 10100 22924 10106 22936
rect 10321 22933 10333 22936
rect 10367 22933 10379 22967
rect 10321 22927 10379 22933
rect 10594 22924 10600 22976
rect 10652 22924 10658 22976
rect 10980 22973 11008 23072
rect 11333 23069 11345 23103
rect 11379 23100 11391 23103
rect 11790 23100 11796 23112
rect 11379 23072 11796 23100
rect 11379 23069 11391 23072
rect 11333 23063 11391 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14568 23100 14596 23199
rect 15028 23177 15056 23208
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23137 15071 23171
rect 15013 23131 15071 23137
rect 15102 23128 15108 23180
rect 15160 23128 15166 23180
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 19306 23168 19334 23208
rect 20070 23168 20076 23180
rect 15344 23140 15516 23168
rect 15344 23128 15350 23140
rect 14323 23072 14596 23100
rect 14921 23103 14979 23109
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14921 23069 14933 23103
rect 14967 23100 14979 23103
rect 15378 23100 15384 23112
rect 14967 23072 15384 23100
rect 14967 23069 14979 23072
rect 14921 23063 14979 23069
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15488 23109 15516 23140
rect 16408 23140 18276 23168
rect 19306 23140 20076 23168
rect 16408 23112 16436 23140
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 16390 23100 16396 23112
rect 15519 23072 16396 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17037 23103 17095 23109
rect 17037 23100 17049 23103
rect 16816 23072 17049 23100
rect 16816 23060 16822 23072
rect 17037 23069 17049 23072
rect 17083 23100 17095 23103
rect 17218 23100 17224 23112
rect 17083 23072 17224 23100
rect 17083 23069 17095 23072
rect 17037 23063 17095 23069
rect 17218 23060 17224 23072
rect 17276 23060 17282 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17972 23072 18153 23100
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 17494 23032 17500 23044
rect 14516 23004 17500 23032
rect 14516 22992 14522 23004
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 17972 22976 18000 23072
rect 18141 23069 18153 23072
rect 18187 23069 18199 23103
rect 18141 23063 18199 23069
rect 18046 22992 18052 23044
rect 18104 22992 18110 23044
rect 10965 22967 11023 22973
rect 10965 22933 10977 22967
rect 11011 22933 11023 22967
rect 10965 22927 11023 22933
rect 11422 22924 11428 22976
rect 11480 22924 11486 22976
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 17034 22964 17040 22976
rect 14700 22936 17040 22964
rect 14700 22924 14706 22936
rect 17034 22924 17040 22936
rect 17092 22924 17098 22976
rect 17313 22967 17371 22973
rect 17313 22933 17325 22967
rect 17359 22964 17371 22967
rect 17770 22964 17776 22976
rect 17359 22936 17776 22964
rect 17359 22933 17371 22936
rect 17313 22927 17371 22933
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 17954 22924 17960 22976
rect 18012 22924 18018 22976
rect 18248 22964 18276 23140
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 19242 23060 19248 23112
rect 19300 23060 19306 23112
rect 19518 22992 19524 23044
rect 19576 22992 19582 23044
rect 20824 23032 20852 23276
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 21048 23276 21189 23304
rect 21048 23264 21054 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 21450 23264 21456 23316
rect 21508 23264 21514 23316
rect 24210 23264 24216 23316
rect 24268 23264 24274 23316
rect 29178 23264 29184 23316
rect 29236 23264 29242 23316
rect 30006 23304 30012 23316
rect 29656 23276 30012 23304
rect 21468 23236 21496 23264
rect 21008 23208 21496 23236
rect 23860 23208 25728 23236
rect 21008 23180 21036 23208
rect 20990 23128 20996 23180
rect 21048 23128 21054 23180
rect 21266 23128 21272 23180
rect 21324 23168 21330 23180
rect 21729 23171 21787 23177
rect 21729 23168 21741 23171
rect 21324 23140 21741 23168
rect 21324 23128 21330 23140
rect 21729 23137 21741 23140
rect 21775 23137 21787 23171
rect 23860 23168 23888 23208
rect 21729 23131 21787 23137
rect 22066 23140 23888 23168
rect 21542 23060 21548 23112
rect 21600 23060 21606 23112
rect 22066 23032 22094 23140
rect 22462 23060 22468 23112
rect 22520 23060 22526 23112
rect 25590 23060 25596 23112
rect 25648 23060 25654 23112
rect 25700 23100 25728 23208
rect 26605 23171 26663 23177
rect 26605 23137 26617 23171
rect 26651 23168 26663 23171
rect 27801 23171 27859 23177
rect 27801 23168 27813 23171
rect 26651 23140 27813 23168
rect 26651 23137 26663 23140
rect 26605 23131 26663 23137
rect 27801 23137 27813 23140
rect 27847 23168 27859 23171
rect 29656 23168 29684 23276
rect 30006 23264 30012 23276
rect 30064 23264 30070 23316
rect 30282 23264 30288 23316
rect 30340 23304 30346 23316
rect 32217 23307 32275 23313
rect 32217 23304 32229 23307
rect 30340 23276 32229 23304
rect 30340 23264 30346 23276
rect 32217 23273 32229 23276
rect 32263 23273 32275 23307
rect 33229 23307 33287 23313
rect 33229 23304 33241 23307
rect 32217 23267 32275 23273
rect 32600 23276 33241 23304
rect 30852 23208 32352 23236
rect 27847 23140 28856 23168
rect 27847 23137 27859 23140
rect 27801 23131 27859 23137
rect 25777 23103 25835 23109
rect 25777 23100 25789 23103
rect 25700 23072 25789 23100
rect 25777 23069 25789 23072
rect 25823 23100 25835 23103
rect 25866 23100 25872 23112
rect 25823 23072 25872 23100
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 26786 23060 26792 23112
rect 26844 23060 26850 23112
rect 28074 23060 28080 23112
rect 28132 23060 28138 23112
rect 28828 23109 28856 23140
rect 29472 23140 29684 23168
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23069 28871 23103
rect 29472 23100 29500 23140
rect 30466 23128 30472 23180
rect 30524 23168 30530 23180
rect 30852 23168 30880 23208
rect 30524 23140 30880 23168
rect 30524 23128 30530 23140
rect 31662 23128 31668 23180
rect 31720 23168 31726 23180
rect 31720 23140 32168 23168
rect 31720 23128 31726 23140
rect 28813 23063 28871 23069
rect 28920 23072 29500 23100
rect 19628 23004 20010 23032
rect 20824 23004 22094 23032
rect 19628 22964 19656 23004
rect 18248 22936 19656 22964
rect 19904 22964 19932 23004
rect 22738 22992 22744 23044
rect 22796 22992 22802 23044
rect 24026 23032 24032 23044
rect 23966 23004 24032 23032
rect 24026 22992 24032 23004
rect 24084 22992 24090 23044
rect 24118 22992 24124 23044
rect 24176 23032 24182 23044
rect 24486 23032 24492 23044
rect 24176 23004 24492 23032
rect 24176 22992 24182 23004
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 28721 23035 28779 23041
rect 28721 23001 28733 23035
rect 28767 23032 28779 23035
rect 28920 23032 28948 23072
rect 29546 23060 29552 23112
rect 29604 23060 29610 23112
rect 32140 23109 32168 23140
rect 32324 23109 32352 23208
rect 31941 23103 31999 23109
rect 31941 23100 31953 23103
rect 31312 23072 31953 23100
rect 28767 23004 28948 23032
rect 28767 23001 28779 23004
rect 28721 22995 28779 23001
rect 28994 22992 29000 23044
rect 29052 22992 29058 23044
rect 29822 22992 29828 23044
rect 29880 22992 29886 23044
rect 29932 23004 30314 23032
rect 20346 22964 20352 22976
rect 19904 22936 20352 22964
rect 20346 22924 20352 22936
rect 20404 22964 20410 22976
rect 20898 22964 20904 22976
rect 20404 22936 20904 22964
rect 20404 22924 20410 22936
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 21910 22964 21916 22976
rect 21683 22936 21916 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 24044 22964 24072 22992
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24044 22936 24593 22964
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 26881 22967 26939 22973
rect 26881 22933 26893 22967
rect 26927 22964 26939 22967
rect 29086 22964 29092 22976
rect 26927 22936 29092 22964
rect 26927 22933 26939 22936
rect 26881 22927 26939 22933
rect 29086 22924 29092 22936
rect 29144 22924 29150 22976
rect 29178 22924 29184 22976
rect 29236 22964 29242 22976
rect 29932 22964 29960 23004
rect 29236 22936 29960 22964
rect 29236 22924 29242 22936
rect 30190 22924 30196 22976
rect 30248 22964 30254 22976
rect 31312 22973 31340 23072
rect 31941 23069 31953 23072
rect 31987 23069 31999 23103
rect 31941 23063 31999 23069
rect 32125 23103 32183 23109
rect 32125 23069 32137 23103
rect 32171 23069 32183 23103
rect 32125 23063 32183 23069
rect 32309 23103 32367 23109
rect 32309 23069 32321 23103
rect 32355 23069 32367 23103
rect 32309 23063 32367 23069
rect 32600 22976 32628 23276
rect 33229 23273 33241 23276
rect 33275 23273 33287 23307
rect 33229 23267 33287 23273
rect 33413 23307 33471 23313
rect 33413 23273 33425 23307
rect 33459 23304 33471 23307
rect 33459 23276 34100 23304
rect 33459 23273 33471 23276
rect 33413 23267 33471 23273
rect 33244 23168 33272 23267
rect 33781 23239 33839 23245
rect 33781 23205 33793 23239
rect 33827 23236 33839 23239
rect 33827 23208 33916 23236
rect 33827 23205 33839 23208
rect 33781 23199 33839 23205
rect 33244 23140 33640 23168
rect 33612 23109 33640 23140
rect 33888 23112 33916 23208
rect 34072 23112 34100 23276
rect 37090 23264 37096 23316
rect 37148 23264 37154 23316
rect 37001 23171 37059 23177
rect 37001 23137 37013 23171
rect 37047 23168 37059 23171
rect 37108 23168 37136 23264
rect 37047 23140 37136 23168
rect 37277 23171 37335 23177
rect 37047 23137 37059 23140
rect 37001 23131 37059 23137
rect 37277 23137 37289 23171
rect 37323 23168 37335 23171
rect 37366 23168 37372 23180
rect 37323 23140 37372 23168
rect 37323 23137 37335 23140
rect 37277 23131 37335 23137
rect 37366 23128 37372 23140
rect 37424 23128 37430 23180
rect 43162 23128 43168 23180
rect 43220 23128 43226 23180
rect 33505 23103 33563 23109
rect 33505 23100 33517 23103
rect 32968 23072 33517 23100
rect 32968 22976 32996 23072
rect 33505 23069 33517 23072
rect 33551 23069 33563 23103
rect 33505 23063 33563 23069
rect 33597 23103 33655 23109
rect 33597 23069 33609 23103
rect 33643 23069 33655 23103
rect 33597 23063 33655 23069
rect 33870 23060 33876 23112
rect 33928 23060 33934 23112
rect 34054 23060 34060 23112
rect 34112 23060 34118 23112
rect 34514 23060 34520 23112
rect 34572 23060 34578 23112
rect 35342 23060 35348 23112
rect 35400 23100 35406 23112
rect 35713 23103 35771 23109
rect 35713 23100 35725 23103
rect 35400 23072 35725 23100
rect 35400 23060 35406 23072
rect 35713 23069 35725 23072
rect 35759 23069 35771 23103
rect 35713 23063 35771 23069
rect 42794 23060 42800 23112
rect 42852 23100 42858 23112
rect 43073 23103 43131 23109
rect 43073 23100 43085 23103
rect 42852 23072 43085 23100
rect 42852 23060 42858 23072
rect 43073 23069 43085 23072
rect 43119 23100 43131 23103
rect 43254 23100 43260 23112
rect 43119 23072 43260 23100
rect 43119 23069 43131 23072
rect 43073 23063 43131 23069
rect 43254 23060 43260 23072
rect 43312 23060 43318 23112
rect 33045 23035 33103 23041
rect 33045 23001 33057 23035
rect 33091 23032 33103 23035
rect 33781 23035 33839 23041
rect 33781 23032 33793 23035
rect 33091 23004 33793 23032
rect 33091 23001 33103 23004
rect 33045 22995 33103 23001
rect 33781 23001 33793 23004
rect 33827 23032 33839 23035
rect 34532 23032 34560 23060
rect 33827 23004 34560 23032
rect 33827 23001 33839 23004
rect 33781 22995 33839 23001
rect 37274 22992 37280 23044
rect 37332 23032 37338 23044
rect 37332 23004 37766 23032
rect 37332 22992 37338 23004
rect 31297 22967 31355 22973
rect 31297 22964 31309 22967
rect 30248 22936 31309 22964
rect 30248 22924 30254 22936
rect 31297 22933 31309 22936
rect 31343 22933 31355 22967
rect 31297 22927 31355 22933
rect 31386 22924 31392 22976
rect 31444 22924 31450 22976
rect 32582 22924 32588 22976
rect 32640 22924 32646 22976
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 33245 22967 33303 22973
rect 33245 22964 33257 22967
rect 33008 22936 33257 22964
rect 33008 22924 33014 22936
rect 33245 22933 33257 22936
rect 33291 22933 33303 22967
rect 33245 22927 33303 22933
rect 34238 22924 34244 22976
rect 34296 22924 34302 22976
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 35161 22967 35219 22973
rect 35161 22964 35173 22967
rect 34848 22936 35173 22964
rect 34848 22924 34854 22936
rect 35161 22933 35173 22936
rect 35207 22933 35219 22967
rect 35161 22927 35219 22933
rect 38746 22924 38752 22976
rect 38804 22924 38810 22976
rect 42705 22967 42763 22973
rect 42705 22933 42717 22967
rect 42751 22964 42763 22967
rect 42794 22964 42800 22976
rect 42751 22936 42800 22964
rect 42751 22933 42763 22936
rect 42705 22927 42763 22933
rect 42794 22924 42800 22936
rect 42852 22924 42858 22976
rect 1104 22874 44620 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 44620 22874
rect 1104 22800 44620 22822
rect 10042 22760 10048 22772
rect 9784 22732 10048 22760
rect 9784 22701 9812 22732
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 10502 22720 10508 22772
rect 10560 22760 10566 22772
rect 11517 22763 11575 22769
rect 11517 22760 11529 22763
rect 10560 22732 11529 22760
rect 10560 22720 10566 22732
rect 11517 22729 11529 22732
rect 11563 22729 11575 22763
rect 16485 22763 16543 22769
rect 11517 22723 11575 22729
rect 11992 22732 16436 22760
rect 9769 22695 9827 22701
rect 9769 22661 9781 22695
rect 9815 22661 9827 22695
rect 9769 22655 9827 22661
rect 10870 22584 10876 22636
rect 10928 22584 10934 22636
rect 11882 22584 11888 22636
rect 11940 22584 11946 22636
rect 7742 22516 7748 22568
rect 7800 22556 7806 22568
rect 9493 22559 9551 22565
rect 9493 22556 9505 22559
rect 7800 22528 9505 22556
rect 7800 22516 7806 22528
rect 9493 22525 9505 22528
rect 9539 22525 9551 22559
rect 9493 22519 9551 22525
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22556 11299 22559
rect 11900 22556 11928 22584
rect 11992 22568 12020 22732
rect 13357 22695 13415 22701
rect 13357 22661 13369 22695
rect 13403 22692 13415 22695
rect 14918 22692 14924 22704
rect 13403 22664 14924 22692
rect 13403 22661 13415 22664
rect 13357 22655 13415 22661
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22624 13323 22627
rect 13446 22624 13452 22636
rect 13311 22596 13452 22624
rect 13311 22593 13323 22596
rect 13265 22587 13323 22593
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22593 16359 22627
rect 16301 22587 16359 22593
rect 11287 22528 11928 22556
rect 11287 22525 11299 22528
rect 11241 22519 11299 22525
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 12161 22559 12219 22565
rect 12161 22525 12173 22559
rect 12207 22556 12219 22559
rect 12986 22556 12992 22568
rect 12207 22528 12992 22556
rect 12207 22525 12219 22528
rect 12161 22519 12219 22525
rect 12986 22516 12992 22528
rect 13044 22556 13050 22568
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13044 22528 13553 22556
rect 13044 22516 13050 22528
rect 13541 22525 13553 22528
rect 13587 22556 13599 22559
rect 15838 22556 15844 22568
rect 13587 22528 15844 22556
rect 13587 22525 13599 22528
rect 13541 22519 13599 22525
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 12894 22380 12900 22432
rect 12952 22380 12958 22432
rect 16316 22420 16344 22587
rect 16408 22488 16436 22732
rect 16485 22729 16497 22763
rect 16531 22729 16543 22763
rect 19153 22763 19211 22769
rect 16485 22723 16543 22729
rect 17052 22732 18276 22760
rect 16500 22692 16528 22723
rect 17052 22704 17080 22732
rect 16945 22695 17003 22701
rect 16945 22692 16957 22695
rect 16500 22664 16957 22692
rect 16945 22661 16957 22664
rect 16991 22661 17003 22695
rect 16945 22655 17003 22661
rect 17034 22652 17040 22704
rect 17092 22652 17098 22704
rect 17402 22652 17408 22704
rect 17460 22652 17466 22704
rect 18248 22692 18276 22732
rect 19153 22729 19165 22763
rect 19199 22760 19211 22763
rect 19426 22760 19432 22772
rect 19199 22732 19432 22760
rect 19199 22729 19211 22732
rect 19153 22723 19211 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 20990 22760 20996 22772
rect 19668 22732 20996 22760
rect 19668 22720 19674 22732
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 23017 22763 23075 22769
rect 23017 22760 23029 22763
rect 22796 22732 23029 22760
rect 22796 22720 22802 22732
rect 23017 22729 23029 22732
rect 23063 22729 23075 22763
rect 23017 22723 23075 22729
rect 23658 22720 23664 22772
rect 23716 22720 23722 22772
rect 24673 22763 24731 22769
rect 24673 22729 24685 22763
rect 24719 22760 24731 22763
rect 25590 22760 25596 22772
rect 24719 22732 25596 22760
rect 24719 22729 24731 22732
rect 24673 22723 24731 22729
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 26786 22760 26792 22772
rect 25823 22732 26792 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 26786 22720 26792 22732
rect 26844 22720 26850 22772
rect 28169 22763 28227 22769
rect 28169 22729 28181 22763
rect 28215 22760 28227 22763
rect 28994 22760 29000 22772
rect 28215 22732 29000 22760
rect 28215 22729 28227 22732
rect 28169 22723 28227 22729
rect 28994 22720 29000 22732
rect 29052 22720 29058 22772
rect 29365 22763 29423 22769
rect 29365 22729 29377 22763
rect 29411 22760 29423 22763
rect 29822 22760 29828 22772
rect 29411 22732 29828 22760
rect 29411 22729 29423 22732
rect 29365 22723 29423 22729
rect 29822 22720 29828 22732
rect 29880 22720 29886 22772
rect 31386 22760 31392 22772
rect 30208 22732 31392 22760
rect 24118 22692 24124 22704
rect 18248 22664 24124 22692
rect 24118 22652 24124 22664
rect 24176 22652 24182 22704
rect 24872 22664 25820 22692
rect 19702 22628 19708 22636
rect 19306 22624 19708 22628
rect 18984 22600 19708 22624
rect 18984 22596 19334 22600
rect 16666 22516 16672 22568
rect 16724 22516 16730 22568
rect 18984 22565 19012 22596
rect 19702 22584 19708 22600
rect 19760 22584 19766 22636
rect 19794 22584 19800 22636
rect 19852 22584 19858 22636
rect 22002 22584 22008 22636
rect 22060 22584 22066 22636
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22624 23259 22627
rect 23247 22596 23336 22624
rect 23247 22593 23259 22596
rect 23201 22587 23259 22593
rect 18969 22559 19027 22565
rect 16776 22528 18000 22556
rect 16776 22488 16804 22528
rect 16408 22460 16804 22488
rect 17972 22488 18000 22528
rect 18969 22525 18981 22559
rect 19015 22525 19027 22559
rect 18969 22519 19027 22525
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22556 19119 22559
rect 19107 22528 19656 22556
rect 19107 22525 19119 22528
rect 19061 22519 19119 22525
rect 19288 22488 19294 22500
rect 17972 22460 19294 22488
rect 19288 22448 19294 22460
rect 19346 22448 19352 22500
rect 19628 22488 19656 22528
rect 19702 22488 19708 22500
rect 19628 22460 19708 22488
rect 19702 22448 19708 22460
rect 19760 22448 19766 22500
rect 23308 22497 23336 22596
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 24872 22633 24900 22664
rect 24857 22627 24915 22633
rect 23440 22596 24808 22624
rect 23440 22584 23446 22596
rect 23750 22516 23756 22568
rect 23808 22516 23814 22568
rect 23934 22516 23940 22568
rect 23992 22516 23998 22568
rect 24780 22556 24808 22596
rect 24857 22593 24869 22627
rect 24903 22593 24915 22627
rect 25409 22627 25467 22633
rect 25409 22624 25421 22627
rect 24857 22587 24915 22593
rect 24964 22596 25421 22624
rect 24964 22556 24992 22596
rect 25409 22593 25421 22596
rect 25455 22624 25467 22627
rect 25682 22624 25688 22636
rect 25455 22596 25688 22624
rect 25455 22593 25467 22596
rect 25409 22587 25467 22593
rect 25682 22584 25688 22596
rect 25740 22584 25746 22636
rect 25792 22624 25820 22664
rect 25866 22652 25872 22704
rect 25924 22692 25930 22704
rect 30101 22695 30159 22701
rect 30101 22692 30113 22695
rect 25924 22664 26096 22692
rect 25924 22652 25930 22664
rect 26068 22633 26096 22664
rect 29564 22664 30113 22692
rect 26053 22627 26111 22633
rect 25792 22596 26004 22624
rect 24780 22528 24992 22556
rect 25133 22559 25191 22565
rect 25133 22525 25145 22559
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 25501 22559 25559 22565
rect 25501 22525 25513 22559
rect 25547 22556 25559 22559
rect 25869 22559 25927 22565
rect 25869 22556 25881 22559
rect 25547 22528 25881 22556
rect 25547 22525 25559 22528
rect 25501 22519 25559 22525
rect 25869 22525 25881 22528
rect 25915 22525 25927 22559
rect 25976 22556 26004 22596
rect 26053 22593 26065 22627
rect 26099 22593 26111 22627
rect 26053 22587 26111 22593
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 26329 22627 26387 22633
rect 26329 22624 26341 22627
rect 26200 22596 26341 22624
rect 26200 22584 26206 22596
rect 26329 22593 26341 22596
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 28074 22584 28080 22636
rect 28132 22622 28138 22636
rect 28132 22594 28175 22622
rect 28132 22584 28138 22594
rect 29270 22584 29276 22636
rect 29328 22584 29334 22636
rect 29564 22633 29592 22664
rect 30101 22661 30113 22664
rect 30147 22661 30159 22695
rect 30101 22655 30159 22661
rect 29549 22627 29607 22633
rect 29549 22593 29561 22627
rect 29595 22593 29607 22627
rect 29549 22587 29607 22593
rect 29638 22584 29644 22636
rect 29696 22584 29702 22636
rect 29733 22627 29791 22633
rect 29733 22593 29745 22627
rect 29779 22593 29791 22627
rect 29733 22587 29791 22593
rect 26160 22556 26188 22584
rect 25976 22528 26188 22556
rect 29288 22556 29316 22584
rect 29748 22556 29776 22587
rect 29822 22584 29828 22636
rect 29880 22633 29886 22636
rect 29880 22627 29909 22633
rect 29897 22593 29909 22627
rect 29880 22587 29909 22593
rect 30009 22627 30067 22633
rect 30009 22593 30021 22627
rect 30055 22624 30067 22627
rect 30208 22624 30236 22732
rect 31386 22720 31392 22732
rect 31444 22720 31450 22772
rect 31662 22720 31668 22772
rect 31720 22720 31726 22772
rect 32582 22720 32588 22772
rect 32640 22720 32646 22772
rect 32950 22720 32956 22772
rect 33008 22720 33014 22772
rect 34054 22720 34060 22772
rect 34112 22720 34118 22772
rect 34238 22720 34244 22772
rect 34296 22720 34302 22772
rect 35342 22720 35348 22772
rect 35400 22720 35406 22772
rect 37550 22720 37556 22772
rect 37608 22720 37614 22772
rect 37921 22763 37979 22769
rect 37921 22729 37933 22763
rect 37967 22760 37979 22763
rect 38746 22760 38752 22772
rect 37967 22732 38752 22760
rect 37967 22729 37979 22732
rect 37921 22723 37979 22729
rect 38746 22720 38752 22732
rect 38804 22720 38810 22772
rect 40126 22760 40132 22772
rect 39592 22732 40132 22760
rect 30392 22664 30788 22692
rect 30392 22636 30420 22664
rect 30055 22596 30236 22624
rect 30285 22627 30343 22633
rect 30055 22593 30067 22596
rect 30009 22587 30067 22593
rect 30285 22593 30297 22627
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 29880 22584 29886 22587
rect 29288 22528 29776 22556
rect 25869 22519 25927 22525
rect 23293 22491 23351 22497
rect 23293 22457 23305 22491
rect 23339 22457 23351 22491
rect 25148 22488 25176 22519
rect 30098 22516 30104 22568
rect 30156 22556 30162 22568
rect 30300 22556 30328 22587
rect 30374 22584 30380 22636
rect 30432 22584 30438 22636
rect 30466 22584 30472 22636
rect 30524 22584 30530 22636
rect 30558 22584 30564 22636
rect 30616 22584 30622 22636
rect 30650 22584 30656 22636
rect 30708 22584 30714 22636
rect 30760 22633 30788 22664
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22593 30803 22627
rect 30745 22587 30803 22593
rect 31680 22556 31708 22720
rect 32861 22695 32919 22701
rect 32140 22664 32720 22692
rect 32140 22633 32168 22664
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 30156 22528 31708 22556
rect 30156 22516 30162 22528
rect 31754 22516 31760 22568
rect 31812 22556 31818 22568
rect 32140 22556 32168 22587
rect 32214 22584 32220 22636
rect 32272 22584 32278 22636
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32692 22633 32720 22664
rect 32861 22661 32873 22695
rect 32907 22661 32919 22695
rect 32861 22655 32919 22661
rect 32677 22627 32735 22633
rect 32677 22593 32689 22627
rect 32723 22593 32735 22627
rect 32677 22587 32735 22593
rect 31812 22528 32168 22556
rect 31812 22516 31818 22528
rect 25774 22488 25780 22500
rect 25148 22460 25780 22488
rect 23293 22451 23351 22457
rect 25774 22448 25780 22460
rect 25832 22488 25838 22500
rect 26145 22491 26203 22497
rect 26145 22488 26157 22491
rect 25832 22460 26157 22488
rect 25832 22448 25838 22460
rect 26145 22457 26157 22460
rect 26191 22457 26203 22491
rect 26145 22451 26203 22457
rect 26237 22491 26295 22497
rect 26237 22457 26249 22491
rect 26283 22457 26295 22491
rect 26237 22451 26295 22457
rect 17586 22420 17592 22432
rect 16316 22392 17592 22420
rect 17586 22380 17592 22392
rect 17644 22380 17650 22432
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18417 22423 18475 22429
rect 18417 22420 18429 22423
rect 18012 22392 18429 22420
rect 18012 22380 18018 22392
rect 18417 22389 18429 22392
rect 18463 22389 18475 22423
rect 18417 22383 18475 22389
rect 19518 22380 19524 22432
rect 19576 22380 19582 22432
rect 19613 22423 19671 22429
rect 19613 22389 19625 22423
rect 19659 22420 19671 22423
rect 20162 22420 20168 22432
rect 19659 22392 20168 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 20162 22380 20168 22392
rect 20220 22380 20226 22432
rect 21818 22380 21824 22432
rect 21876 22380 21882 22432
rect 25041 22423 25099 22429
rect 25041 22389 25053 22423
rect 25087 22420 25099 22423
rect 25314 22420 25320 22432
rect 25087 22392 25320 22420
rect 25087 22389 25099 22392
rect 25041 22383 25099 22389
rect 25314 22380 25320 22392
rect 25372 22420 25378 22432
rect 26252 22420 26280 22451
rect 29822 22448 29828 22500
rect 29880 22488 29886 22500
rect 30558 22488 30564 22500
rect 29880 22460 30564 22488
rect 29880 22448 29886 22460
rect 30558 22448 30564 22460
rect 30616 22448 30622 22500
rect 32398 22488 32404 22500
rect 31220 22460 32404 22488
rect 31220 22432 31248 22460
rect 32398 22448 32404 22460
rect 32456 22488 32462 22500
rect 32876 22488 32904 22655
rect 32953 22627 33011 22633
rect 32953 22593 32965 22627
rect 32999 22593 33011 22627
rect 32953 22587 33011 22593
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 32456 22460 32904 22488
rect 32456 22448 32462 22460
rect 25372 22392 26280 22420
rect 25372 22380 25378 22392
rect 31202 22380 31208 22432
rect 31260 22380 31266 22432
rect 32214 22380 32220 22432
rect 32272 22420 32278 22432
rect 32968 22420 32996 22587
rect 33704 22488 33732 22587
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 34072 22624 34100 22720
rect 34149 22627 34207 22633
rect 34149 22624 34161 22627
rect 34072 22596 34161 22624
rect 34149 22593 34161 22596
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34256 22556 34284 22720
rect 35802 22652 35808 22704
rect 35860 22652 35866 22704
rect 38010 22652 38016 22704
rect 38068 22652 38074 22704
rect 34698 22584 34704 22636
rect 34756 22624 34762 22636
rect 35069 22627 35127 22633
rect 35069 22624 35081 22627
rect 34756 22596 35081 22624
rect 34756 22584 34762 22596
rect 35069 22593 35081 22596
rect 35115 22593 35127 22627
rect 35069 22587 35127 22593
rect 34977 22559 35035 22565
rect 34977 22556 34989 22559
rect 34256 22528 34989 22556
rect 34977 22525 34989 22528
rect 35023 22525 35035 22559
rect 34977 22519 35035 22525
rect 35084 22488 35112 22587
rect 37090 22584 37096 22636
rect 37148 22584 37154 22636
rect 39592 22633 39620 22732
rect 40126 22720 40132 22732
rect 40184 22720 40190 22772
rect 40037 22695 40095 22701
rect 40037 22661 40049 22695
rect 40083 22661 40095 22695
rect 40402 22692 40408 22704
rect 40037 22655 40095 22661
rect 40328 22664 40408 22692
rect 39577 22627 39635 22633
rect 39577 22593 39589 22627
rect 39623 22593 39635 22627
rect 40052 22624 40080 22655
rect 40328 22633 40356 22664
rect 40402 22652 40408 22664
rect 40460 22652 40466 22704
rect 43254 22652 43260 22704
rect 43312 22692 43318 22704
rect 43349 22695 43407 22701
rect 43349 22692 43361 22695
rect 43312 22664 43361 22692
rect 43312 22652 43318 22664
rect 43349 22661 43361 22664
rect 43395 22661 43407 22695
rect 43349 22655 43407 22661
rect 39577 22587 39635 22593
rect 39684 22596 40080 22624
rect 40313 22627 40371 22633
rect 36814 22516 36820 22568
rect 36872 22516 36878 22568
rect 38102 22516 38108 22568
rect 38160 22556 38166 22568
rect 39298 22556 39304 22568
rect 38160 22528 39304 22556
rect 38160 22516 38166 22528
rect 39298 22516 39304 22528
rect 39356 22516 39362 22568
rect 39684 22565 39712 22596
rect 40313 22593 40325 22627
rect 40359 22593 40371 22627
rect 40313 22587 40371 22593
rect 43070 22584 43076 22636
rect 43128 22624 43134 22636
rect 43438 22624 43444 22636
rect 43128 22596 43444 22624
rect 43128 22584 43134 22596
rect 43438 22584 43444 22596
rect 43496 22584 43502 22636
rect 39669 22559 39727 22565
rect 39669 22525 39681 22559
rect 39715 22525 39727 22559
rect 39669 22519 39727 22525
rect 39850 22516 39856 22568
rect 39908 22556 39914 22568
rect 40037 22559 40095 22565
rect 40037 22556 40049 22559
rect 39908 22528 40049 22556
rect 39908 22516 39914 22528
rect 40037 22525 40049 22528
rect 40083 22556 40095 22559
rect 40083 22528 41000 22556
rect 40083 22525 40095 22528
rect 40037 22519 40095 22525
rect 40972 22500 41000 22528
rect 43162 22516 43168 22568
rect 43220 22516 43226 22568
rect 33704 22460 35112 22488
rect 39942 22448 39948 22500
rect 40000 22448 40006 22500
rect 40954 22448 40960 22500
rect 41012 22448 41018 22500
rect 32272 22392 32996 22420
rect 34333 22423 34391 22429
rect 32272 22380 32278 22392
rect 34333 22389 34345 22423
rect 34379 22420 34391 22423
rect 34514 22420 34520 22432
rect 34379 22392 34520 22420
rect 34379 22389 34391 22392
rect 34333 22383 34391 22389
rect 34514 22380 34520 22392
rect 34572 22380 34578 22432
rect 34698 22380 34704 22432
rect 34756 22380 34762 22432
rect 40218 22380 40224 22432
rect 40276 22420 40282 22432
rect 41138 22420 41144 22432
rect 40276 22392 41144 22420
rect 40276 22380 40282 22392
rect 41138 22380 41144 22392
rect 41196 22420 41202 22432
rect 41690 22420 41696 22432
rect 41196 22392 41696 22420
rect 41196 22380 41202 22392
rect 41690 22380 41696 22392
rect 41748 22420 41754 22432
rect 42889 22423 42947 22429
rect 42889 22420 42901 22423
rect 41748 22392 42901 22420
rect 41748 22380 41754 22392
rect 42889 22389 42901 22392
rect 42935 22389 42947 22423
rect 42889 22383 42947 22389
rect 43346 22380 43352 22432
rect 43404 22380 43410 22432
rect 1104 22330 44620 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 44620 22330
rect 1104 22256 44620 22278
rect 10124 22219 10182 22225
rect 10124 22185 10136 22219
rect 10170 22216 10182 22219
rect 10594 22216 10600 22228
rect 10170 22188 10600 22216
rect 10170 22185 10182 22188
rect 10124 22179 10182 22185
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 11609 22219 11667 22225
rect 11609 22185 11621 22219
rect 11655 22216 11667 22219
rect 11790 22216 11796 22228
rect 11655 22188 11796 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 11790 22176 11796 22188
rect 11848 22176 11854 22228
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 13633 22219 13691 22225
rect 13633 22216 13645 22219
rect 13504 22188 13645 22216
rect 13504 22176 13510 22188
rect 13633 22185 13645 22188
rect 13679 22185 13691 22219
rect 13633 22179 13691 22185
rect 17586 22176 17592 22228
rect 17644 22176 17650 22228
rect 21256 22219 21314 22225
rect 18156 22188 21128 22216
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22080 9919 22083
rect 11146 22080 11152 22092
rect 9907 22052 11152 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 11146 22040 11152 22052
rect 11204 22080 11210 22092
rect 11885 22083 11943 22089
rect 11885 22080 11897 22083
rect 11204 22052 11897 22080
rect 11204 22040 11210 22052
rect 11885 22049 11897 22052
rect 11931 22049 11943 22083
rect 11885 22043 11943 22049
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12308 22052 13308 22080
rect 12308 22040 12314 22052
rect 13280 21998 13308 22052
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 13596 22052 15393 22080
rect 13596 22040 13602 22052
rect 15381 22049 15393 22052
rect 15427 22080 15439 22083
rect 18049 22083 18107 22089
rect 15427 22052 16712 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 16684 22024 16712 22052
rect 18049 22049 18061 22083
rect 18095 22080 18107 22083
rect 18156 22080 18184 22188
rect 19978 22148 19984 22160
rect 18248 22120 19984 22148
rect 18248 22089 18276 22120
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 18095 22052 18184 22080
rect 18233 22083 18291 22089
rect 18095 22049 18107 22052
rect 18049 22043 18107 22049
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 21100 22080 21128 22188
rect 21256 22185 21268 22219
rect 21302 22216 21314 22219
rect 21818 22216 21824 22228
rect 21302 22188 21824 22216
rect 21302 22185 21314 22188
rect 21256 22179 21314 22185
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 22296 22188 25176 22216
rect 22296 22080 22324 22188
rect 25148 22160 25176 22188
rect 25314 22176 25320 22228
rect 25372 22176 25378 22228
rect 25685 22219 25743 22225
rect 25685 22185 25697 22219
rect 25731 22216 25743 22219
rect 25958 22216 25964 22228
rect 25731 22188 25964 22216
rect 25731 22185 25743 22188
rect 25685 22179 25743 22185
rect 25958 22176 25964 22188
rect 26016 22176 26022 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 26513 22219 26571 22225
rect 26513 22216 26525 22219
rect 26292 22188 26525 22216
rect 26292 22176 26298 22188
rect 26513 22185 26525 22188
rect 26559 22185 26571 22219
rect 26513 22179 26571 22185
rect 26789 22219 26847 22225
rect 26789 22185 26801 22219
rect 26835 22216 26847 22219
rect 28074 22216 28080 22228
rect 26835 22188 28080 22216
rect 26835 22185 26847 22188
rect 26789 22179 26847 22185
rect 28074 22176 28080 22188
rect 28132 22176 28138 22228
rect 28534 22176 28540 22228
rect 28592 22216 28598 22228
rect 28902 22216 28908 22228
rect 28592 22188 28908 22216
rect 28592 22176 28598 22188
rect 28902 22176 28908 22188
rect 28960 22176 28966 22228
rect 29914 22176 29920 22228
rect 29972 22176 29978 22228
rect 34422 22176 34428 22228
rect 34480 22216 34486 22228
rect 34480 22188 35756 22216
rect 34480 22176 34486 22188
rect 25130 22108 25136 22160
rect 25188 22108 25194 22160
rect 21100 22052 22324 22080
rect 22741 22083 22799 22089
rect 18233 22043 18291 22049
rect 22741 22049 22753 22083
rect 22787 22080 22799 22083
rect 23014 22080 23020 22092
rect 22787 22052 23020 22080
rect 22787 22049 22799 22052
rect 22741 22043 22799 22049
rect 16666 21972 16672 22024
rect 16724 21972 16730 22024
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 17678 22012 17684 22024
rect 16816 21984 17684 22012
rect 16816 21972 16822 21984
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 17954 21972 17960 22024
rect 18012 21972 18018 22024
rect 10870 21904 10876 21956
rect 10928 21904 10934 21956
rect 12161 21947 12219 21953
rect 12161 21913 12173 21947
rect 12207 21944 12219 21947
rect 12434 21944 12440 21956
rect 12207 21916 12440 21944
rect 12207 21913 12219 21916
rect 12161 21907 12219 21913
rect 12434 21904 12440 21916
rect 12492 21904 12498 21956
rect 15654 21904 15660 21956
rect 15712 21904 15718 21956
rect 17770 21904 17776 21956
rect 17828 21944 17834 21956
rect 18248 21944 18276 22043
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 20993 22015 21051 22021
rect 20993 22012 21005 22015
rect 20036 21984 21005 22012
rect 20036 21972 20042 21984
rect 20993 21981 21005 21984
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 22370 21972 22376 22024
rect 22428 21972 22434 22024
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23842 22012 23848 22024
rect 23440 21984 23848 22012
rect 23440 21972 23446 21984
rect 23842 21972 23848 21984
rect 23900 22012 23906 22024
rect 24949 22015 25007 22021
rect 24949 22012 24961 22015
rect 23900 21984 24961 22012
rect 23900 21972 23906 21984
rect 24949 21981 24961 21984
rect 24995 22012 25007 22015
rect 25038 22012 25044 22024
rect 24995 21984 25044 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 25332 22012 25360 22176
rect 25869 22151 25927 22157
rect 25869 22117 25881 22151
rect 25915 22148 25927 22151
rect 26050 22148 26056 22160
rect 25915 22120 26056 22148
rect 25915 22117 25927 22120
rect 25869 22111 25927 22117
rect 26050 22108 26056 22120
rect 26108 22108 26114 22160
rect 28810 22108 28816 22160
rect 28868 22108 28874 22160
rect 34606 22148 34612 22160
rect 32232 22120 34612 22148
rect 25593 22083 25651 22089
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 28828 22080 28856 22108
rect 32232 22092 32260 22120
rect 34606 22108 34612 22120
rect 34664 22108 34670 22160
rect 35728 22148 35756 22188
rect 35802 22176 35808 22228
rect 35860 22216 35866 22228
rect 36262 22216 36268 22228
rect 35860 22188 36268 22216
rect 35860 22176 35866 22188
rect 36262 22176 36268 22188
rect 36320 22176 36326 22228
rect 40402 22176 40408 22228
rect 40460 22216 40466 22228
rect 41230 22216 41236 22228
rect 40460 22188 41236 22216
rect 40460 22176 40466 22188
rect 41230 22176 41236 22188
rect 41288 22216 41294 22228
rect 41288 22188 41368 22216
rect 41288 22176 41294 22188
rect 38838 22148 38844 22160
rect 35728 22120 38844 22148
rect 38838 22108 38844 22120
rect 38896 22108 38902 22160
rect 40494 22108 40500 22160
rect 40552 22108 40558 22160
rect 25639 22052 25912 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25884 22024 25912 22052
rect 26344 22052 28856 22080
rect 26344 22024 26372 22052
rect 29086 22040 29092 22092
rect 29144 22080 29150 22092
rect 29144 22052 29868 22080
rect 29144 22040 29150 22052
rect 25409 22015 25467 22021
rect 25409 22012 25421 22015
rect 25332 21984 25421 22012
rect 25409 21981 25421 21984
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 25682 21972 25688 22024
rect 25740 21972 25746 22024
rect 25866 21972 25872 22024
rect 25924 21972 25930 22024
rect 26326 21972 26332 22024
rect 26384 21972 26390 22024
rect 28534 21972 28540 22024
rect 28592 21972 28598 22024
rect 28721 22015 28779 22021
rect 28721 22014 28733 22015
rect 28644 21986 28733 22014
rect 28644 21956 28672 21986
rect 28721 21981 28733 21986
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 28948 21974 28954 22026
rect 29006 22012 29012 22026
rect 29840 22024 29868 22052
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 32214 22080 32220 22092
rect 31168 22052 32220 22080
rect 31168 22040 31174 22052
rect 32214 22040 32220 22052
rect 32272 22040 32278 22092
rect 34146 22040 34152 22092
rect 34204 22080 34210 22092
rect 35437 22083 35495 22089
rect 35437 22080 35449 22083
rect 34204 22052 35449 22080
rect 34204 22040 34210 22052
rect 35437 22049 35449 22052
rect 35483 22049 35495 22083
rect 35437 22043 35495 22049
rect 40126 22040 40132 22092
rect 40184 22080 40190 22092
rect 40313 22083 40371 22089
rect 40313 22080 40325 22083
rect 40184 22052 40325 22080
rect 40184 22040 40190 22052
rect 40313 22049 40325 22052
rect 40359 22080 40371 22083
rect 40359 22052 40724 22080
rect 40359 22049 40371 22052
rect 40313 22043 40371 22049
rect 29546 22012 29552 22024
rect 29006 21984 29552 22012
rect 29006 21974 29012 21984
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 29822 21972 29828 22024
rect 29880 21972 29886 22024
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 22012 30159 22015
rect 30282 22012 30288 22024
rect 30147 21984 30288 22012
rect 30147 21981 30159 21984
rect 30101 21975 30159 21981
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 30742 21972 30748 22024
rect 30800 22012 30806 22024
rect 30837 22015 30895 22021
rect 30837 22012 30849 22015
rect 30800 21984 30849 22012
rect 30800 21972 30806 21984
rect 30837 21981 30849 21984
rect 30883 21981 30895 22015
rect 30837 21975 30895 21981
rect 31570 21972 31576 22024
rect 31628 22012 31634 22024
rect 31628 21984 32352 22012
rect 31628 21972 31634 21984
rect 32324 21956 32352 21984
rect 34238 21972 34244 22024
rect 34296 22012 34302 22024
rect 34606 22012 34612 22024
rect 34296 21984 34612 22012
rect 34296 21972 34302 21984
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 34698 21972 34704 22024
rect 34756 21972 34762 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 34977 22015 35035 22021
rect 34977 22012 34989 22015
rect 34848 21984 34989 22012
rect 34848 21972 34854 21984
rect 34977 21981 34989 21984
rect 35023 21981 35035 22015
rect 34977 21975 35035 21981
rect 35069 22015 35127 22021
rect 35069 21981 35081 22015
rect 35115 22012 35127 22015
rect 35342 22012 35348 22024
rect 35115 21984 35348 22012
rect 35115 21981 35127 21984
rect 35069 21975 35127 21981
rect 17828 21916 18276 21944
rect 17828 21904 17834 21916
rect 24854 21904 24860 21956
rect 24912 21944 24918 21956
rect 25133 21947 25191 21953
rect 25133 21944 25145 21947
rect 24912 21916 25145 21944
rect 24912 21904 24918 21916
rect 25133 21913 25145 21916
rect 25179 21913 25191 21947
rect 25133 21907 25191 21913
rect 27798 21904 27804 21956
rect 27856 21944 27862 21956
rect 27856 21916 28212 21944
rect 27856 21904 27862 21916
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 12250 21876 12256 21888
rect 11112 21848 12256 21876
rect 11112 21836 11118 21848
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 17129 21879 17187 21885
rect 17129 21845 17141 21879
rect 17175 21876 17187 21879
rect 17954 21876 17960 21888
rect 17175 21848 17960 21876
rect 17175 21845 17187 21848
rect 17129 21839 17187 21845
rect 17954 21836 17960 21848
rect 18012 21876 18018 21888
rect 19150 21876 19156 21888
rect 18012 21848 19156 21876
rect 18012 21836 18018 21848
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 26510 21876 26516 21888
rect 22244 21848 26516 21876
rect 22244 21836 22250 21848
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 28184 21876 28212 21916
rect 28258 21904 28264 21956
rect 28316 21904 28322 21956
rect 28626 21904 28632 21956
rect 28684 21904 28690 21956
rect 28810 21904 28816 21956
rect 28868 21944 28874 21956
rect 30929 21947 30987 21953
rect 30929 21944 30941 21947
rect 28868 21916 30941 21944
rect 28868 21904 28874 21916
rect 30929 21913 30941 21916
rect 30975 21944 30987 21947
rect 31754 21944 31760 21956
rect 30975 21916 31760 21944
rect 30975 21913 30987 21916
rect 30929 21907 30987 21913
rect 31754 21904 31760 21916
rect 31812 21944 31818 21956
rect 32214 21944 32220 21956
rect 31812 21916 32220 21944
rect 31812 21904 31818 21916
rect 32214 21904 32220 21916
rect 32272 21904 32278 21956
rect 32306 21904 32312 21956
rect 32364 21944 32370 21956
rect 34885 21947 34943 21953
rect 34885 21944 34897 21947
rect 32364 21916 34897 21944
rect 32364 21904 32370 21916
rect 34885 21913 34897 21916
rect 34931 21913 34943 21947
rect 34885 21907 34943 21913
rect 28997 21879 29055 21885
rect 28997 21876 29009 21879
rect 28184 21848 29009 21876
rect 28997 21845 29009 21848
rect 29043 21876 29055 21879
rect 29178 21876 29184 21888
rect 29043 21848 29184 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29178 21836 29184 21848
rect 29236 21836 29242 21888
rect 32030 21836 32036 21888
rect 32088 21876 32094 21888
rect 35084 21876 35112 21975
rect 35342 21972 35348 21984
rect 35400 21972 35406 22024
rect 35526 21972 35532 22024
rect 35584 21972 35590 22024
rect 40218 21972 40224 22024
rect 40276 22012 40282 22024
rect 40696 22021 40724 22052
rect 40954 22040 40960 22092
rect 41012 22080 41018 22092
rect 41049 22083 41107 22089
rect 41049 22080 41061 22083
rect 41012 22052 41061 22080
rect 41012 22040 41018 22052
rect 41049 22049 41061 22052
rect 41095 22049 41107 22083
rect 41049 22043 41107 22049
rect 41138 22040 41144 22092
rect 41196 22040 41202 22092
rect 41230 22040 41236 22092
rect 41288 22040 41294 22092
rect 41340 22080 41368 22188
rect 42886 22108 42892 22160
rect 42944 22148 42950 22160
rect 43346 22148 43352 22160
rect 42944 22120 43352 22148
rect 42944 22108 42950 22120
rect 43346 22108 43352 22120
rect 43404 22108 43410 22160
rect 41340 22052 41552 22080
rect 40405 22015 40463 22021
rect 40405 22012 40417 22015
rect 40276 21984 40417 22012
rect 40276 21972 40282 21984
rect 40405 21981 40417 21984
rect 40451 21981 40463 22015
rect 40405 21975 40463 21981
rect 40681 22015 40739 22021
rect 40681 21981 40693 22015
rect 40727 21981 40739 22015
rect 40681 21975 40739 21981
rect 40770 21972 40776 22024
rect 40828 21972 40834 22024
rect 40310 21944 40316 21956
rect 35268 21916 36860 21944
rect 35268 21885 35296 21916
rect 36832 21888 36860 21916
rect 40052 21916 40316 21944
rect 32088 21848 35112 21876
rect 35253 21879 35311 21885
rect 32088 21836 32094 21848
rect 35253 21845 35265 21879
rect 35299 21845 35311 21879
rect 35253 21839 35311 21845
rect 36814 21836 36820 21888
rect 36872 21836 36878 21888
rect 39482 21836 39488 21888
rect 39540 21876 39546 21888
rect 40052 21885 40080 21916
rect 40310 21904 40316 21916
rect 40368 21904 40374 21956
rect 40497 21947 40555 21953
rect 40497 21913 40509 21947
rect 40543 21913 40555 21947
rect 40972 21944 41000 22040
rect 41524 22024 41552 22052
rect 42150 22040 42156 22092
rect 42208 22080 42214 22092
rect 44085 22083 44143 22089
rect 42208 22052 43392 22080
rect 42208 22040 42214 22052
rect 41322 21972 41328 22024
rect 41380 21972 41386 22024
rect 41506 21972 41512 22024
rect 41564 21972 41570 22024
rect 41690 21972 41696 22024
rect 41748 21972 41754 22024
rect 41785 22015 41843 22021
rect 41785 21981 41797 22015
rect 41831 21981 41843 22015
rect 41785 21975 41843 21981
rect 41800 21944 41828 21975
rect 42058 21972 42064 22024
rect 42116 22012 42122 22024
rect 42337 22015 42395 22021
rect 42337 22012 42349 22015
rect 42116 21984 42349 22012
rect 42116 21972 42122 21984
rect 42337 21981 42349 21984
rect 42383 21981 42395 22015
rect 42337 21975 42395 21981
rect 42610 21972 42616 22024
rect 42668 21972 42674 22024
rect 42794 21972 42800 22024
rect 42852 21972 42858 22024
rect 43162 21972 43168 22024
rect 43220 21972 43226 22024
rect 43364 22021 43392 22052
rect 44085 22049 44097 22083
rect 44131 22080 44143 22083
rect 44358 22080 44364 22092
rect 44131 22052 44364 22080
rect 44131 22049 44143 22052
rect 44085 22043 44143 22049
rect 44358 22040 44364 22052
rect 44416 22040 44422 22092
rect 43349 22015 43407 22021
rect 43349 21981 43361 22015
rect 43395 22012 43407 22015
rect 43530 22012 43536 22024
rect 43395 21984 43536 22012
rect 43395 21981 43407 21984
rect 43349 21975 43407 21981
rect 43530 21972 43536 21984
rect 43588 21972 43594 22024
rect 43622 21972 43628 22024
rect 43680 21972 43686 22024
rect 43640 21944 43668 21972
rect 40972 21916 43668 21944
rect 40497 21907 40555 21913
rect 40037 21879 40095 21885
rect 40037 21876 40049 21879
rect 39540 21848 40049 21876
rect 39540 21836 39546 21848
rect 40037 21845 40049 21848
rect 40083 21845 40095 21879
rect 40037 21839 40095 21845
rect 40218 21836 40224 21888
rect 40276 21876 40282 21888
rect 40512 21876 40540 21907
rect 40276 21848 40540 21876
rect 40276 21836 40282 21848
rect 40862 21836 40868 21888
rect 40920 21836 40926 21888
rect 41138 21836 41144 21888
rect 41196 21876 41202 21888
rect 41607 21879 41665 21885
rect 41607 21876 41619 21879
rect 41196 21848 41619 21876
rect 41196 21836 41202 21848
rect 41607 21845 41619 21848
rect 41653 21845 41665 21879
rect 41607 21839 41665 21845
rect 42334 21836 42340 21888
rect 42392 21876 42398 21888
rect 42429 21879 42487 21885
rect 42429 21876 42441 21879
rect 42392 21848 42441 21876
rect 42392 21836 42398 21848
rect 42429 21845 42441 21848
rect 42475 21845 42487 21879
rect 42429 21839 42487 21845
rect 43441 21879 43499 21885
rect 43441 21845 43453 21879
rect 43487 21876 43499 21879
rect 43898 21876 43904 21888
rect 43487 21848 43904 21876
rect 43487 21845 43499 21848
rect 43441 21839 43499 21845
rect 43898 21836 43904 21848
rect 43956 21836 43962 21888
rect 1104 21786 44620 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 44620 21786
rect 1104 21712 44620 21734
rect 12434 21632 12440 21684
rect 12492 21632 12498 21684
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 15841 21675 15899 21681
rect 15841 21672 15853 21675
rect 15712 21644 15853 21672
rect 15712 21632 15718 21644
rect 15841 21641 15853 21644
rect 15887 21641 15899 21675
rect 15841 21635 15899 21641
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 17497 21675 17555 21681
rect 17497 21672 17509 21675
rect 16724 21644 17509 21672
rect 16724 21632 16730 21644
rect 17497 21641 17509 21644
rect 17543 21672 17555 21675
rect 17862 21672 17868 21684
rect 17543 21644 17868 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17862 21632 17868 21644
rect 17920 21672 17926 21684
rect 17920 21644 19334 21672
rect 17920 21632 17926 21644
rect 13538 21604 13544 21616
rect 13372 21576 13544 21604
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21536 8171 21539
rect 10502 21536 10508 21548
rect 8159 21508 10508 21536
rect 8159 21505 8171 21508
rect 8113 21499 8171 21505
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 12621 21539 12679 21545
rect 12621 21505 12633 21539
rect 12667 21536 12679 21539
rect 12894 21536 12900 21548
rect 12667 21508 12900 21536
rect 12667 21505 12679 21508
rect 12621 21499 12679 21505
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13078 21496 13084 21548
rect 13136 21496 13142 21548
rect 13372 21545 13400 21576
rect 13538 21564 13544 21576
rect 13596 21564 13602 21616
rect 14366 21564 14372 21616
rect 14424 21564 14430 21616
rect 19306 21604 19334 21644
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 21913 21675 21971 21681
rect 21913 21641 21925 21675
rect 21959 21672 21971 21675
rect 22002 21672 22008 21684
rect 21959 21644 22008 21672
rect 21959 21641 21971 21644
rect 21913 21635 21971 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22278 21632 22284 21684
rect 22336 21632 22342 21684
rect 24026 21632 24032 21684
rect 24084 21672 24090 21684
rect 24084 21644 28212 21672
rect 24084 21632 24090 21644
rect 19996 21604 20024 21632
rect 19306 21576 20024 21604
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 16022 21496 16028 21548
rect 16080 21496 16086 21548
rect 18782 21496 18788 21548
rect 18840 21496 18846 21548
rect 19628 21545 19656 21576
rect 20346 21564 20352 21616
rect 20404 21564 20410 21616
rect 21174 21564 21180 21616
rect 21232 21604 21238 21616
rect 21634 21604 21640 21616
rect 21232 21576 21640 21604
rect 21232 21564 21238 21576
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 26234 21604 26240 21616
rect 22066 21576 23612 21604
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21505 19671 21539
rect 22066 21536 22094 21576
rect 23584 21548 23612 21576
rect 25884 21576 26240 21604
rect 19613 21499 19671 21505
rect 21100 21508 22094 21536
rect 22373 21539 22431 21545
rect 13633 21471 13691 21477
rect 13633 21468 13645 21471
rect 13280 21440 13645 21468
rect 13280 21409 13308 21440
rect 13633 21437 13645 21440
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15381 21471 15439 21477
rect 15381 21468 15393 21471
rect 15160 21440 15393 21468
rect 15160 21428 15166 21440
rect 15381 21437 15393 21440
rect 15427 21468 15439 21471
rect 15427 21440 16528 21468
rect 15427 21437 15439 21440
rect 15381 21431 15439 21437
rect 13265 21403 13323 21409
rect 13265 21369 13277 21403
rect 13311 21369 13323 21403
rect 13265 21363 13323 21369
rect 6825 21335 6883 21341
rect 6825 21301 6837 21335
rect 6871 21332 6883 21335
rect 6914 21332 6920 21344
rect 6871 21304 6920 21332
rect 6871 21301 6883 21304
rect 6825 21295 6883 21301
rect 6914 21292 6920 21304
rect 6972 21332 6978 21344
rect 7742 21332 7748 21344
rect 6972 21304 7748 21332
rect 6972 21292 6978 21304
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 16500 21332 16528 21440
rect 19886 21428 19892 21480
rect 19944 21428 19950 21480
rect 21100 21332 21128 21508
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22738 21536 22744 21548
rect 22419 21508 22744 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23290 21496 23296 21548
rect 23348 21496 23354 21548
rect 23566 21496 23572 21548
rect 23624 21496 23630 21548
rect 25884 21545 25912 21576
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 28184 21604 28212 21644
rect 28258 21632 28264 21684
rect 28316 21672 28322 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 28316 21644 28365 21672
rect 28316 21632 28322 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28626 21632 28632 21684
rect 28684 21632 28690 21684
rect 36354 21672 36360 21684
rect 28966 21644 36360 21672
rect 28644 21604 28672 21632
rect 28966 21604 28994 21644
rect 36354 21632 36360 21644
rect 36412 21632 36418 21684
rect 40034 21672 40040 21684
rect 38672 21644 40040 21672
rect 28184 21576 28994 21604
rect 33226 21564 33232 21616
rect 33284 21604 33290 21616
rect 33778 21604 33784 21616
rect 33284 21576 33784 21604
rect 33284 21564 33290 21576
rect 33778 21564 33784 21576
rect 33836 21564 33842 21616
rect 34514 21604 34520 21616
rect 34440 21576 34520 21604
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 26053 21499 26111 21505
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21536 27767 21539
rect 28074 21536 28080 21548
rect 27755 21508 28080 21536
rect 27755 21505 27767 21508
rect 27709 21499 27767 21505
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 22557 21471 22615 21477
rect 22557 21468 22569 21471
rect 21324 21440 22569 21468
rect 21324 21428 21330 21440
rect 22557 21437 22569 21440
rect 22603 21468 22615 21471
rect 23934 21468 23940 21480
rect 22603 21440 23940 21468
rect 22603 21437 22615 21440
rect 22557 21431 22615 21437
rect 23934 21428 23940 21440
rect 23992 21428 23998 21480
rect 26068 21468 26096 21499
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 28350 21496 28356 21548
rect 28408 21536 28414 21548
rect 28537 21539 28595 21545
rect 28537 21536 28549 21539
rect 28408 21508 28549 21536
rect 28408 21496 28414 21508
rect 28537 21505 28549 21508
rect 28583 21505 28595 21539
rect 28537 21499 28595 21505
rect 28629 21539 28687 21545
rect 28629 21505 28641 21539
rect 28675 21505 28687 21539
rect 28629 21499 28687 21505
rect 25884 21440 26096 21468
rect 28261 21471 28319 21477
rect 25884 21344 25912 21440
rect 28261 21437 28273 21471
rect 28307 21468 28319 21471
rect 28644 21468 28672 21499
rect 28718 21496 28724 21548
rect 28776 21496 28782 21548
rect 28902 21496 28908 21548
rect 28960 21496 28966 21548
rect 31938 21496 31944 21548
rect 31996 21496 32002 21548
rect 33962 21496 33968 21548
rect 34020 21536 34026 21548
rect 34440 21545 34468 21576
rect 34514 21564 34520 21576
rect 34572 21564 34578 21616
rect 38672 21545 38700 21644
rect 40034 21632 40040 21644
rect 40092 21632 40098 21684
rect 40862 21632 40868 21684
rect 40920 21632 40926 21684
rect 41138 21632 41144 21684
rect 41196 21632 41202 21684
rect 41506 21632 41512 21684
rect 41564 21632 41570 21684
rect 42978 21632 42984 21684
rect 43036 21672 43042 21684
rect 43441 21675 43499 21681
rect 43441 21672 43453 21675
rect 43036 21644 43453 21672
rect 43036 21632 43042 21644
rect 43441 21641 43453 21644
rect 43487 21641 43499 21675
rect 43441 21635 43499 21641
rect 43530 21632 43536 21684
rect 43588 21632 43594 21684
rect 39853 21607 39911 21613
rect 39853 21604 39865 21607
rect 38764 21576 39865 21604
rect 38764 21548 38792 21576
rect 39853 21573 39865 21576
rect 39899 21573 39911 21607
rect 39853 21567 39911 21573
rect 34241 21539 34299 21545
rect 34241 21536 34253 21539
rect 34020 21508 34253 21536
rect 34020 21496 34026 21508
rect 34241 21505 34253 21508
rect 34287 21505 34299 21539
rect 34241 21499 34299 21505
rect 34425 21539 34483 21545
rect 34425 21505 34437 21539
rect 34471 21505 34483 21539
rect 34425 21499 34483 21505
rect 38657 21539 38715 21545
rect 38657 21505 38669 21539
rect 38703 21505 38715 21539
rect 38657 21499 38715 21505
rect 38746 21496 38752 21548
rect 38804 21496 38810 21548
rect 38933 21539 38991 21545
rect 38933 21505 38945 21539
rect 38979 21536 38991 21539
rect 39482 21536 39488 21548
rect 38979 21508 39488 21536
rect 38979 21505 38991 21508
rect 38933 21499 38991 21505
rect 39482 21496 39488 21508
rect 39540 21496 39546 21548
rect 39574 21496 39580 21548
rect 39632 21536 39638 21548
rect 39761 21539 39819 21545
rect 39761 21536 39773 21539
rect 39632 21508 39773 21536
rect 39632 21496 39638 21508
rect 39761 21505 39773 21508
rect 39807 21505 39819 21539
rect 39761 21499 39819 21505
rect 28307 21440 28672 21468
rect 28307 21437 28319 21440
rect 28261 21431 28319 21437
rect 38838 21428 38844 21480
rect 38896 21468 38902 21480
rect 38896 21440 39252 21468
rect 38896 21428 38902 21440
rect 34054 21360 34060 21412
rect 34112 21400 34118 21412
rect 39224 21400 39252 21440
rect 39298 21428 39304 21480
rect 39356 21468 39362 21480
rect 39669 21471 39727 21477
rect 39669 21468 39681 21471
rect 39356 21440 39681 21468
rect 39356 21428 39362 21440
rect 39669 21437 39681 21440
rect 39715 21437 39727 21471
rect 39868 21468 39896 21567
rect 39942 21564 39948 21616
rect 40000 21564 40006 21616
rect 40126 21496 40132 21548
rect 40184 21496 40190 21548
rect 40218 21496 40224 21548
rect 40276 21496 40282 21548
rect 40586 21496 40592 21548
rect 40644 21496 40650 21548
rect 40773 21539 40831 21545
rect 40773 21505 40785 21539
rect 40819 21536 40831 21539
rect 40880 21536 40908 21632
rect 40819 21508 40908 21536
rect 40819 21505 40831 21508
rect 40773 21499 40831 21505
rect 39942 21468 39948 21480
rect 39868 21440 39948 21468
rect 39669 21431 39727 21437
rect 39942 21428 39948 21440
rect 40000 21428 40006 21480
rect 39850 21400 39856 21412
rect 34112 21372 34468 21400
rect 39224 21372 39856 21400
rect 34112 21360 34118 21372
rect 34440 21344 34468 21372
rect 39850 21360 39856 21372
rect 39908 21360 39914 21412
rect 40144 21400 40172 21496
rect 40865 21471 40923 21477
rect 40865 21437 40877 21471
rect 40911 21468 40923 21471
rect 41156 21468 41184 21632
rect 41233 21539 41291 21545
rect 41233 21505 41245 21539
rect 41279 21536 41291 21539
rect 41524 21536 41552 21632
rect 42812 21576 43116 21604
rect 41279 21508 41552 21536
rect 41601 21539 41659 21545
rect 41279 21505 41291 21508
rect 41233 21499 41291 21505
rect 41601 21505 41613 21539
rect 41647 21536 41659 21539
rect 42426 21536 42432 21548
rect 41647 21508 42432 21536
rect 41647 21505 41659 21508
rect 41601 21499 41659 21505
rect 42426 21496 42432 21508
rect 42484 21496 42490 21548
rect 42518 21496 42524 21548
rect 42576 21536 42582 21548
rect 42812 21545 42840 21576
rect 43088 21548 43116 21576
rect 42797 21539 42855 21545
rect 42797 21536 42809 21539
rect 42576 21508 42809 21536
rect 42576 21496 42582 21508
rect 42797 21505 42809 21508
rect 42843 21505 42855 21539
rect 42797 21499 42855 21505
rect 42886 21496 42892 21548
rect 42944 21496 42950 21548
rect 43070 21496 43076 21548
rect 43128 21496 43134 21548
rect 43257 21539 43315 21545
rect 43257 21505 43269 21539
rect 43303 21536 43315 21539
rect 43438 21536 43444 21548
rect 43303 21508 43444 21536
rect 43303 21505 43315 21508
rect 43257 21499 43315 21505
rect 43438 21496 43444 21508
rect 43496 21496 43502 21548
rect 43548 21545 43576 21632
rect 43533 21539 43591 21545
rect 43533 21505 43545 21539
rect 43579 21505 43591 21539
rect 43533 21499 43591 21505
rect 43622 21496 43628 21548
rect 43680 21496 43686 21548
rect 40911 21440 41184 21468
rect 41325 21471 41383 21477
rect 40911 21437 40923 21440
rect 40865 21431 40923 21437
rect 41325 21437 41337 21471
rect 41371 21468 41383 21471
rect 41414 21468 41420 21480
rect 41371 21440 41420 21468
rect 41371 21437 41383 21440
rect 41325 21431 41383 21437
rect 41414 21428 41420 21440
rect 41472 21428 41478 21480
rect 41509 21471 41567 21477
rect 41509 21437 41521 21471
rect 41555 21437 41567 21471
rect 41509 21431 41567 21437
rect 41230 21400 41236 21412
rect 40144 21372 41236 21400
rect 41230 21360 41236 21372
rect 41288 21400 41294 21412
rect 41524 21400 41552 21431
rect 41690 21428 41696 21480
rect 41748 21468 41754 21480
rect 42058 21468 42064 21480
rect 41748 21440 42064 21468
rect 41748 21428 41754 21440
rect 42058 21428 42064 21440
rect 42116 21428 42122 21480
rect 42705 21471 42763 21477
rect 42705 21437 42717 21471
rect 42751 21437 42763 21471
rect 42705 21431 42763 21437
rect 42981 21471 43039 21477
rect 42981 21437 42993 21471
rect 43027 21468 43039 21471
rect 43640 21468 43668 21496
rect 43027 21440 43668 21468
rect 43027 21437 43039 21440
rect 42981 21431 43039 21437
rect 41288 21372 41552 21400
rect 41288 21360 41294 21372
rect 41966 21360 41972 21412
rect 42024 21360 42030 21412
rect 16500 21304 21128 21332
rect 23106 21292 23112 21344
rect 23164 21292 23170 21344
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 25958 21292 25964 21344
rect 26016 21292 26022 21344
rect 28626 21292 28632 21344
rect 28684 21332 28690 21344
rect 29178 21332 29184 21344
rect 28684 21304 29184 21332
rect 28684 21292 28690 21304
rect 29178 21292 29184 21304
rect 29236 21292 29242 21344
rect 29546 21292 29552 21344
rect 29604 21332 29610 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 29604 21304 30665 21332
rect 29604 21292 29610 21304
rect 30653 21301 30665 21304
rect 30699 21332 30711 21335
rect 30834 21332 30840 21344
rect 30699 21304 30840 21332
rect 30699 21301 30711 21304
rect 30653 21295 30711 21301
rect 30834 21292 30840 21304
rect 30892 21292 30898 21344
rect 34330 21292 34336 21344
rect 34388 21292 34394 21344
rect 34422 21292 34428 21344
rect 34480 21292 34486 21344
rect 39114 21292 39120 21344
rect 39172 21292 39178 21344
rect 39390 21292 39396 21344
rect 39448 21332 39454 21344
rect 40218 21332 40224 21344
rect 39448 21304 40224 21332
rect 39448 21292 39454 21304
rect 40218 21292 40224 21304
rect 40276 21292 40282 21344
rect 40402 21292 40408 21344
rect 40460 21292 40466 21344
rect 41322 21292 41328 21344
rect 41380 21332 41386 21344
rect 42720 21332 42748 21431
rect 41380 21304 42748 21332
rect 41380 21292 41386 21304
rect 43162 21292 43168 21344
rect 43220 21292 43226 21344
rect 43254 21292 43260 21344
rect 43312 21292 43318 21344
rect 1104 21242 44620 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 44620 21242
rect 1104 21168 44620 21190
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 13136 21100 14105 21128
rect 13136 21088 13142 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14093 21091 14151 21097
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 16080 21100 16681 21128
rect 16080 21088 16086 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 19886 21088 19892 21140
rect 19944 21128 19950 21140
rect 20441 21131 20499 21137
rect 20441 21128 20453 21131
rect 19944 21100 20453 21128
rect 19944 21088 19950 21100
rect 20441 21097 20453 21100
rect 20487 21097 20499 21131
rect 20441 21091 20499 21097
rect 24213 21131 24271 21137
rect 24213 21097 24225 21131
rect 24259 21128 24271 21131
rect 24578 21128 24584 21140
rect 24259 21100 24584 21128
rect 24259 21097 24271 21100
rect 24213 21091 24271 21097
rect 24578 21088 24584 21100
rect 24636 21088 24642 21140
rect 25958 21088 25964 21140
rect 26016 21088 26022 21140
rect 28718 21088 28724 21140
rect 28776 21128 28782 21140
rect 29089 21131 29147 21137
rect 29089 21128 29101 21131
rect 28776 21100 29101 21128
rect 28776 21088 28782 21100
rect 29089 21097 29101 21100
rect 29135 21097 29147 21131
rect 29089 21091 29147 21097
rect 29178 21088 29184 21140
rect 29236 21088 29242 21140
rect 33229 21131 33287 21137
rect 33229 21097 33241 21131
rect 33275 21128 33287 21131
rect 33962 21128 33968 21140
rect 33275 21100 33968 21128
rect 33275 21097 33287 21100
rect 33229 21091 33287 21097
rect 33962 21088 33968 21100
rect 34020 21088 34026 21140
rect 34146 21088 34152 21140
rect 34204 21088 34210 21140
rect 34330 21088 34336 21140
rect 34388 21088 34394 21140
rect 39574 21088 39580 21140
rect 39632 21088 39638 21140
rect 40034 21088 40040 21140
rect 40092 21128 40098 21140
rect 40221 21131 40279 21137
rect 40221 21128 40233 21131
rect 40092 21100 40233 21128
rect 40092 21088 40098 21100
rect 40221 21097 40233 21100
rect 40267 21128 40279 21131
rect 41322 21128 41328 21140
rect 40267 21100 41328 21128
rect 40267 21097 40279 21100
rect 40221 21091 40279 21097
rect 41322 21088 41328 21100
rect 41380 21088 41386 21140
rect 42150 21128 42156 21140
rect 41524 21100 42156 21128
rect 20717 21063 20775 21069
rect 20717 21029 20729 21063
rect 20763 21029 20775 21063
rect 20717 21023 20775 21029
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 8941 20995 8999 21001
rect 8941 20992 8953 20995
rect 8352 20964 8953 20992
rect 8352 20952 8358 20964
rect 8941 20961 8953 20964
rect 8987 20961 8999 20995
rect 8941 20955 8999 20961
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 17310 20952 17316 21004
rect 17368 20952 17374 21004
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 13964 20896 14473 20924
rect 13964 20884 13970 20896
rect 14461 20893 14473 20896
rect 14507 20924 14519 20927
rect 15102 20924 15108 20936
rect 14507 20896 15108 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 17037 20927 17095 20933
rect 17037 20893 17049 20927
rect 17083 20924 17095 20927
rect 17954 20924 17960 20936
rect 17083 20896 17960 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 18506 20884 18512 20936
rect 18564 20884 18570 20936
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20924 20683 20927
rect 20732 20924 20760 21023
rect 21266 20992 21272 21004
rect 20671 20896 20760 20924
rect 20824 20964 21272 20992
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 20824 20856 20852 20964
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 22462 20952 22468 21004
rect 22520 20952 22526 21004
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23106 20992 23112 21004
rect 22787 20964 23112 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 25869 20995 25927 21001
rect 25869 20961 25881 20995
rect 25915 20992 25927 20995
rect 25976 20992 26004 21088
rect 28353 21063 28411 21069
rect 28353 21029 28365 21063
rect 28399 21060 28411 21063
rect 28902 21060 28908 21072
rect 28399 21032 28908 21060
rect 28399 21029 28411 21032
rect 28353 21023 28411 21029
rect 28902 21020 28908 21032
rect 28960 21020 28966 21072
rect 30006 21060 30012 21072
rect 29012 21032 30012 21060
rect 25915 20964 26004 20992
rect 26145 20995 26203 21001
rect 25915 20961 25927 20964
rect 25869 20955 25927 20961
rect 26145 20961 26157 20995
rect 26191 20992 26203 20995
rect 28166 20992 28172 21004
rect 26191 20964 28172 20992
rect 26191 20961 26203 20964
rect 26145 20955 26203 20961
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 29012 21001 29040 21032
rect 30006 21020 30012 21032
rect 30064 21020 30070 21072
rect 32401 21063 32459 21069
rect 32401 21029 32413 21063
rect 32447 21060 32459 21063
rect 32447 21032 33732 21060
rect 32447 21029 32459 21032
rect 32401 21023 32459 21029
rect 28997 20995 29055 21001
rect 28997 20992 29009 20995
rect 28736 20964 29009 20992
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20924 21143 20927
rect 21634 20924 21640 20936
rect 21131 20896 21640 20924
rect 21131 20893 21143 20896
rect 21085 20887 21143 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 25038 20884 25044 20936
rect 25096 20924 25102 20936
rect 25777 20927 25835 20933
rect 25777 20924 25789 20927
rect 25096 20896 25789 20924
rect 25096 20884 25102 20896
rect 25777 20893 25789 20896
rect 25823 20924 25835 20927
rect 26050 20924 26056 20936
rect 25823 20896 26056 20924
rect 25823 20893 25835 20896
rect 25777 20887 25835 20893
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 24026 20856 24032 20868
rect 20732 20828 20852 20856
rect 23966 20828 24032 20856
rect 20732 20800 20760 20828
rect 24026 20816 24032 20828
rect 24084 20816 24090 20868
rect 9582 20748 9588 20800
rect 9640 20748 9646 20800
rect 14550 20748 14556 20800
rect 14608 20748 14614 20800
rect 17126 20748 17132 20800
rect 17184 20748 17190 20800
rect 18322 20748 18328 20800
rect 18380 20748 18386 20800
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 21174 20748 21180 20800
rect 21232 20748 21238 20800
rect 25958 20748 25964 20800
rect 26016 20788 26022 20800
rect 26970 20788 26976 20800
rect 26016 20760 26976 20788
rect 26016 20748 26022 20760
rect 26970 20748 26976 20760
rect 27028 20748 27034 20800
rect 28184 20788 28212 20952
rect 28534 20884 28540 20936
rect 28592 20884 28598 20936
rect 28626 20884 28632 20936
rect 28684 20884 28690 20936
rect 28736 20933 28764 20964
rect 28997 20961 29009 20964
rect 29043 20961 29055 20995
rect 29822 20992 29828 21004
rect 28997 20955 29055 20961
rect 29288 20964 29828 20992
rect 28721 20927 28779 20933
rect 28721 20893 28733 20927
rect 28767 20893 28779 20927
rect 28721 20887 28779 20893
rect 28810 20884 28816 20936
rect 28868 20884 28874 20936
rect 29288 20933 29316 20964
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 30742 20952 30748 21004
rect 30800 20992 30806 21004
rect 31757 20995 31815 21001
rect 30800 20964 31616 20992
rect 30800 20952 30806 20964
rect 29273 20927 29331 20933
rect 29273 20893 29285 20927
rect 29319 20893 29331 20927
rect 30193 20927 30251 20933
rect 30193 20924 30205 20927
rect 29273 20887 29331 20893
rect 29380 20896 30205 20924
rect 29380 20856 29408 20896
rect 30193 20893 30205 20896
rect 30239 20893 30251 20927
rect 30193 20887 30251 20893
rect 30374 20884 30380 20936
rect 30432 20924 30438 20936
rect 31018 20924 31024 20936
rect 30432 20896 31024 20924
rect 30432 20884 30438 20896
rect 31018 20884 31024 20896
rect 31076 20884 31082 20936
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 31202 20884 31208 20936
rect 31260 20924 31266 20936
rect 31588 20933 31616 20964
rect 31757 20961 31769 20995
rect 31803 20992 31815 20995
rect 32125 20995 32183 21001
rect 32125 20992 32137 20995
rect 31803 20964 32137 20992
rect 31803 20961 31815 20964
rect 31757 20955 31815 20961
rect 32125 20961 32137 20964
rect 32171 20992 32183 20995
rect 33704 20992 33732 21032
rect 32171 20964 32812 20992
rect 32171 20961 32183 20964
rect 32125 20955 32183 20961
rect 31297 20927 31355 20933
rect 31297 20924 31309 20927
rect 31260 20896 31309 20924
rect 31260 20884 31266 20896
rect 31297 20893 31309 20896
rect 31343 20893 31355 20927
rect 31297 20887 31355 20893
rect 31573 20927 31631 20933
rect 31573 20893 31585 20927
rect 31619 20893 31631 20927
rect 31573 20887 31631 20893
rect 31846 20884 31852 20936
rect 31904 20924 31910 20936
rect 32033 20927 32091 20933
rect 32033 20924 32045 20927
rect 31904 20896 32045 20924
rect 31904 20884 31910 20896
rect 32033 20893 32045 20896
rect 32079 20893 32091 20927
rect 32033 20887 32091 20893
rect 28828 20828 29408 20856
rect 28828 20788 28856 20828
rect 29546 20816 29552 20868
rect 29604 20816 29610 20868
rect 29733 20859 29791 20865
rect 29733 20825 29745 20859
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 29917 20859 29975 20865
rect 29917 20825 29929 20859
rect 29963 20856 29975 20859
rect 30009 20859 30067 20865
rect 30009 20856 30021 20859
rect 29963 20828 30021 20856
rect 29963 20825 29975 20828
rect 29917 20819 29975 20825
rect 30009 20825 30021 20828
rect 30055 20825 30067 20859
rect 31128 20856 31156 20884
rect 30009 20819 30067 20825
rect 30576 20828 31156 20856
rect 32048 20856 32076 20887
rect 32214 20884 32220 20936
rect 32272 20924 32278 20936
rect 32784 20933 32812 20964
rect 33060 20964 33339 20992
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 32272 20896 32505 20924
rect 32272 20884 32278 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 32769 20927 32827 20933
rect 32769 20893 32781 20927
rect 32815 20893 32827 20927
rect 32769 20887 32827 20893
rect 32585 20859 32643 20865
rect 32585 20856 32597 20859
rect 32048 20828 32597 20856
rect 28184 20760 28856 20788
rect 29748 20788 29776 20819
rect 30576 20800 30604 20828
rect 32585 20825 32597 20828
rect 32631 20825 32643 20859
rect 32585 20819 32643 20825
rect 29822 20788 29828 20800
rect 29748 20760 29828 20788
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 30558 20748 30564 20800
rect 30616 20748 30622 20800
rect 32950 20748 32956 20800
rect 33008 20748 33014 20800
rect 33060 20788 33088 20964
rect 33311 20933 33339 20964
rect 33520 20964 33732 20992
rect 33137 20927 33195 20933
rect 33137 20893 33149 20927
rect 33183 20924 33195 20927
rect 33311 20927 33379 20933
rect 33183 20896 33272 20924
rect 33311 20896 33333 20927
rect 33183 20893 33195 20896
rect 33137 20887 33195 20893
rect 33244 20868 33272 20896
rect 33321 20893 33333 20896
rect 33367 20893 33379 20927
rect 33321 20887 33379 20893
rect 33413 20927 33471 20933
rect 33413 20893 33425 20927
rect 33459 20926 33471 20927
rect 33520 20926 33548 20964
rect 33704 20933 33732 20964
rect 33459 20898 33548 20926
rect 33597 20927 33655 20933
rect 33459 20893 33471 20898
rect 33413 20887 33471 20893
rect 33597 20893 33609 20927
rect 33643 20893 33655 20927
rect 33597 20887 33655 20893
rect 33689 20927 33747 20933
rect 33689 20893 33701 20927
rect 33735 20893 33747 20927
rect 33689 20887 33747 20893
rect 33873 20927 33931 20933
rect 33873 20893 33885 20927
rect 33919 20924 33931 20927
rect 34164 20924 34192 21088
rect 34348 20992 34376 21088
rect 38473 21063 38531 21069
rect 38473 21029 38485 21063
rect 38519 21060 38531 21063
rect 39022 21060 39028 21072
rect 38519 21032 39028 21060
rect 38519 21029 38531 21032
rect 38473 21023 38531 21029
rect 39022 21020 39028 21032
rect 39080 21020 39086 21072
rect 39592 21060 39620 21088
rect 40770 21060 40776 21072
rect 39132 21032 39528 21060
rect 39592 21032 40776 21060
rect 34348 20964 35020 20992
rect 33919 20896 34192 20924
rect 34517 20927 34575 20933
rect 33919 20893 33931 20896
rect 33873 20887 33931 20893
rect 34517 20893 34529 20927
rect 34563 20924 34575 20927
rect 34606 20924 34612 20936
rect 34563 20896 34612 20924
rect 34563 20893 34575 20896
rect 34517 20887 34575 20893
rect 33226 20816 33232 20868
rect 33284 20816 33290 20868
rect 33502 20816 33508 20868
rect 33560 20816 33566 20868
rect 33612 20856 33640 20887
rect 33888 20856 33916 20887
rect 34606 20884 34612 20896
rect 34664 20924 34670 20936
rect 34992 20933 35020 20964
rect 35618 20952 35624 21004
rect 35676 20992 35682 21004
rect 38562 20992 38568 21004
rect 35676 20964 38568 20992
rect 35676 20952 35682 20964
rect 38562 20952 38568 20964
rect 38620 20952 38626 21004
rect 39132 20992 39160 21032
rect 38672 20964 39160 20992
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 34664 20896 34897 20924
rect 34664 20884 34670 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 34977 20927 35035 20933
rect 34977 20893 34989 20927
rect 35023 20893 35035 20927
rect 34977 20887 35035 20893
rect 35345 20927 35403 20933
rect 35345 20893 35357 20927
rect 35391 20924 35403 20927
rect 35989 20927 36047 20933
rect 35989 20924 36001 20927
rect 35391 20896 36001 20924
rect 35391 20893 35403 20896
rect 35345 20887 35403 20893
rect 35989 20893 36001 20896
rect 36035 20893 36047 20927
rect 35989 20887 36047 20893
rect 36630 20884 36636 20936
rect 36688 20884 36694 20936
rect 38197 20927 38255 20933
rect 38197 20893 38209 20927
rect 38243 20893 38255 20927
rect 38197 20887 38255 20893
rect 33612 20828 33916 20856
rect 33962 20816 33968 20868
rect 34020 20856 34026 20868
rect 34149 20859 34207 20865
rect 34149 20856 34161 20859
rect 34020 20828 34161 20856
rect 34020 20816 34026 20828
rect 34149 20825 34161 20828
rect 34195 20825 34207 20859
rect 34149 20819 34207 20825
rect 34333 20859 34391 20865
rect 34333 20825 34345 20859
rect 34379 20825 34391 20859
rect 34333 20819 34391 20825
rect 33686 20788 33692 20800
rect 33060 20760 33692 20788
rect 33686 20748 33692 20760
rect 33744 20788 33750 20800
rect 34057 20791 34115 20797
rect 34057 20788 34069 20791
rect 33744 20760 34069 20788
rect 33744 20748 33750 20760
rect 34057 20757 34069 20760
rect 34103 20757 34115 20791
rect 34348 20788 34376 20819
rect 34422 20816 34428 20868
rect 34480 20856 34486 20868
rect 35069 20859 35127 20865
rect 35069 20856 35081 20859
rect 34480 20828 35081 20856
rect 34480 20816 34486 20828
rect 35069 20825 35081 20828
rect 35115 20825 35127 20859
rect 35069 20819 35127 20825
rect 35187 20859 35245 20865
rect 35187 20825 35199 20859
rect 35233 20825 35245 20859
rect 35187 20819 35245 20825
rect 34514 20788 34520 20800
rect 34348 20760 34520 20788
rect 34057 20751 34115 20757
rect 34514 20748 34520 20760
rect 34572 20748 34578 20800
rect 34698 20748 34704 20800
rect 34756 20748 34762 20800
rect 34790 20748 34796 20800
rect 34848 20788 34854 20800
rect 35202 20788 35230 20819
rect 34848 20760 35230 20788
rect 38212 20788 38240 20887
rect 38286 20884 38292 20936
rect 38344 20924 38350 20936
rect 38672 20924 38700 20964
rect 39390 20952 39396 21004
rect 39448 20952 39454 21004
rect 39500 20992 39528 21032
rect 40770 21020 40776 21032
rect 40828 21060 40834 21072
rect 41414 21060 41420 21072
rect 40828 21032 41420 21060
rect 40828 21020 40834 21032
rect 41414 21020 41420 21032
rect 41472 21060 41478 21072
rect 41524 21060 41552 21100
rect 42150 21088 42156 21100
rect 42208 21088 42214 21140
rect 43162 21088 43168 21140
rect 43220 21088 43226 21140
rect 43254 21088 43260 21140
rect 43312 21088 43318 21140
rect 42610 21060 42616 21072
rect 41472 21032 41552 21060
rect 41616 21032 42616 21060
rect 41472 21020 41478 21032
rect 39500 20964 39896 20992
rect 38344 20896 38700 20924
rect 38749 20927 38807 20933
rect 38344 20884 38350 20896
rect 38749 20893 38761 20927
rect 38795 20924 38807 20927
rect 38838 20924 38844 20936
rect 38795 20896 38844 20924
rect 38795 20893 38807 20896
rect 38749 20887 38807 20893
rect 38838 20884 38844 20896
rect 38896 20884 38902 20936
rect 38930 20884 38936 20936
rect 38988 20884 38994 20936
rect 38473 20859 38531 20865
rect 38473 20825 38485 20859
rect 38519 20856 38531 20859
rect 39408 20856 39436 20952
rect 39868 20933 39896 20964
rect 39485 20927 39543 20933
rect 39485 20893 39497 20927
rect 39531 20924 39543 20927
rect 39853 20927 39911 20933
rect 39531 20896 39620 20924
rect 39531 20893 39543 20896
rect 39485 20887 39543 20893
rect 38519 20828 39436 20856
rect 38519 20825 38531 20828
rect 38473 20819 38531 20825
rect 39390 20788 39396 20800
rect 38212 20760 39396 20788
rect 34848 20748 34854 20760
rect 39390 20748 39396 20760
rect 39448 20748 39454 20800
rect 39592 20788 39620 20896
rect 39853 20893 39865 20927
rect 39899 20893 39911 20927
rect 39853 20887 39911 20893
rect 39942 20884 39948 20936
rect 40000 20924 40006 20936
rect 40221 20927 40279 20933
rect 40221 20924 40233 20927
rect 40000 20896 40233 20924
rect 40000 20884 40006 20896
rect 40221 20893 40233 20896
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 40310 20884 40316 20936
rect 40368 20924 40374 20936
rect 40405 20927 40463 20933
rect 40405 20924 40417 20927
rect 40368 20896 40417 20924
rect 40368 20884 40374 20896
rect 40405 20893 40417 20896
rect 40451 20893 40463 20927
rect 40405 20887 40463 20893
rect 41417 20927 41475 20933
rect 41417 20893 41429 20927
rect 41463 20924 41475 20927
rect 41616 20924 41644 21032
rect 42610 21020 42616 21032
rect 42668 21020 42674 21072
rect 43272 21060 43300 21088
rect 42996 21032 43300 21060
rect 43349 21063 43407 21069
rect 42245 20995 42303 21001
rect 42245 20961 42257 20995
rect 42291 20992 42303 20995
rect 42886 20992 42892 21004
rect 42291 20964 42892 20992
rect 42291 20961 42303 20964
rect 42245 20955 42303 20961
rect 42886 20952 42892 20964
rect 42944 20952 42950 21004
rect 41463 20896 41644 20924
rect 41463 20893 41475 20896
rect 41417 20887 41475 20893
rect 41230 20816 41236 20868
rect 41288 20856 41294 20868
rect 41432 20856 41460 20887
rect 41690 20884 41696 20936
rect 41748 20884 41754 20936
rect 42150 20884 42156 20936
rect 42208 20884 42214 20936
rect 42518 20884 42524 20936
rect 42576 20884 42582 20936
rect 42610 20884 42616 20936
rect 42668 20884 42674 20936
rect 42996 20933 43024 21032
rect 43349 21029 43361 21063
rect 43395 21029 43407 21063
rect 43349 21023 43407 21029
rect 43257 20995 43315 21001
rect 43257 20961 43269 20995
rect 43303 20992 43315 20995
rect 43364 20992 43392 21023
rect 43303 20964 43392 20992
rect 43303 20961 43315 20964
rect 43257 20955 43315 20961
rect 42981 20927 43039 20933
rect 42981 20893 42993 20927
rect 43027 20893 43039 20927
rect 42981 20887 43039 20893
rect 43070 20884 43076 20936
rect 43128 20884 43134 20936
rect 43346 20884 43352 20936
rect 43404 20884 43410 20936
rect 43622 20884 43628 20936
rect 43680 20884 43686 20936
rect 41288 20828 41460 20856
rect 41288 20816 41294 20828
rect 40037 20791 40095 20797
rect 40037 20788 40049 20791
rect 39592 20760 40049 20788
rect 40037 20757 40049 20760
rect 40083 20757 40095 20791
rect 40037 20751 40095 20757
rect 40218 20748 40224 20800
rect 40276 20788 40282 20800
rect 41708 20788 41736 20884
rect 41877 20859 41935 20865
rect 41877 20825 41889 20859
rect 41923 20856 41935 20859
rect 43088 20856 43116 20884
rect 43533 20859 43591 20865
rect 43533 20856 43545 20859
rect 41923 20828 43024 20856
rect 43088 20828 43545 20856
rect 41923 20825 41935 20828
rect 41877 20819 41935 20825
rect 42996 20800 43024 20828
rect 43533 20825 43545 20828
rect 43579 20825 43591 20859
rect 43533 20819 43591 20825
rect 42242 20788 42248 20800
rect 40276 20760 42248 20788
rect 40276 20748 40282 20760
rect 42242 20748 42248 20760
rect 42300 20748 42306 20800
rect 42797 20791 42855 20797
rect 42797 20757 42809 20791
rect 42843 20788 42855 20791
rect 42886 20788 42892 20800
rect 42843 20760 42892 20788
rect 42843 20757 42855 20760
rect 42797 20751 42855 20757
rect 42886 20748 42892 20760
rect 42944 20748 42950 20800
rect 42978 20748 42984 20800
rect 43036 20748 43042 20800
rect 1104 20698 44620 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 44620 20698
rect 1104 20624 44620 20646
rect 11517 20587 11575 20593
rect 11517 20553 11529 20587
rect 11563 20553 11575 20587
rect 11517 20547 11575 20553
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 11974 20584 11980 20596
rect 11931 20556 11980 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 11532 20448 11560 20547
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 14608 20556 14933 20584
rect 14608 20544 14614 20556
rect 14921 20553 14933 20556
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20553 15623 20587
rect 15565 20547 15623 20553
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16206 20584 16212 20596
rect 15979 20556 16212 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 14642 20516 14648 20528
rect 10919 20420 11560 20448
rect 11900 20488 14648 20516
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 8110 20340 8116 20392
rect 8168 20380 8174 20392
rect 11900 20380 11928 20488
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 11977 20451 12035 20457
rect 11977 20417 11989 20451
rect 12023 20448 12035 20451
rect 12342 20448 12348 20460
rect 12023 20420 12348 20448
rect 12023 20417 12035 20420
rect 11977 20411 12035 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13722 20448 13728 20460
rect 13311 20420 13728 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15580 20448 15608 20547
rect 16206 20544 16212 20556
rect 16264 20544 16270 20596
rect 19702 20544 19708 20596
rect 19760 20584 19766 20596
rect 20622 20584 20628 20596
rect 19760 20556 20628 20584
rect 19760 20544 19766 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 23109 20587 23167 20593
rect 23109 20553 23121 20587
rect 23155 20584 23167 20587
rect 23290 20584 23296 20596
rect 23155 20556 23296 20584
rect 23155 20553 23167 20556
rect 23109 20547 23167 20553
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23474 20544 23480 20596
rect 23532 20544 23538 20596
rect 28534 20544 28540 20596
rect 28592 20584 28598 20596
rect 28813 20587 28871 20593
rect 28813 20584 28825 20587
rect 28592 20556 28825 20584
rect 28592 20544 28598 20556
rect 28813 20553 28825 20556
rect 28859 20584 28871 20587
rect 29822 20584 29828 20596
rect 28859 20556 29828 20584
rect 28859 20553 28871 20556
rect 28813 20547 28871 20553
rect 29822 20544 29828 20556
rect 29880 20584 29886 20596
rect 29880 20556 30880 20584
rect 29880 20544 29886 20556
rect 18233 20519 18291 20525
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 18322 20516 18328 20528
rect 18279 20488 18328 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 20346 20516 20352 20528
rect 19458 20488 20352 20516
rect 20346 20476 20352 20488
rect 20404 20516 20410 20528
rect 22554 20516 22560 20528
rect 20404 20488 22560 20516
rect 20404 20476 20410 20488
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 30561 20519 30619 20525
rect 28184 20488 28764 20516
rect 28184 20460 28212 20488
rect 15335 20420 15608 20448
rect 15664 20420 16252 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 8168 20352 11928 20380
rect 8168 20340 8174 20352
rect 12066 20340 12072 20392
rect 12124 20340 12130 20392
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15664 20380 15692 20420
rect 14792 20352 15692 20380
rect 14792 20340 14798 20352
rect 16022 20340 16028 20392
rect 16080 20340 16086 20392
rect 16224 20389 16252 20420
rect 17862 20408 17868 20460
rect 17920 20448 17926 20460
rect 17957 20451 18015 20457
rect 17957 20448 17969 20451
rect 17920 20420 17969 20448
rect 17920 20408 17926 20420
rect 17957 20417 17969 20420
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 20990 20408 20996 20460
rect 21048 20408 21054 20460
rect 28166 20408 28172 20460
rect 28224 20408 28230 20460
rect 28350 20408 28356 20460
rect 28408 20448 28414 20460
rect 28736 20457 28764 20488
rect 28920 20488 30328 20516
rect 28920 20457 28948 20488
rect 30300 20460 30328 20488
rect 30561 20485 30573 20519
rect 30607 20485 30619 20519
rect 30561 20479 30619 20485
rect 28445 20451 28503 20457
rect 28445 20448 28457 20451
rect 28408 20420 28457 20448
rect 28408 20408 28414 20420
rect 28445 20417 28457 20420
rect 28491 20417 28503 20451
rect 28445 20411 28503 20417
rect 28721 20451 28779 20457
rect 28721 20417 28733 20451
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 28905 20451 28963 20457
rect 28905 20417 28917 20451
rect 28951 20417 28963 20451
rect 28905 20411 28963 20417
rect 28994 20408 29000 20460
rect 29052 20408 29058 20460
rect 29546 20408 29552 20460
rect 29604 20408 29610 20460
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 30190 20408 30196 20460
rect 30248 20408 30254 20460
rect 30282 20408 30288 20460
rect 30340 20408 30346 20460
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20448 30435 20451
rect 30576 20448 30604 20479
rect 30852 20457 30880 20556
rect 33962 20544 33968 20596
rect 34020 20544 34026 20596
rect 34606 20544 34612 20596
rect 34664 20544 34670 20596
rect 36630 20544 36636 20596
rect 36688 20544 36694 20596
rect 37277 20587 37335 20593
rect 37277 20553 37289 20587
rect 37323 20553 37335 20587
rect 37277 20547 37335 20553
rect 33505 20519 33563 20525
rect 33505 20485 33517 20519
rect 33551 20516 33563 20519
rect 33551 20488 33916 20516
rect 33551 20485 33563 20488
rect 33505 20479 33563 20485
rect 30423 20420 30604 20448
rect 30837 20451 30895 20457
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 30837 20417 30849 20451
rect 30883 20417 30895 20451
rect 30837 20411 30895 20417
rect 31294 20408 31300 20460
rect 31352 20408 31358 20460
rect 33413 20451 33471 20457
rect 33413 20417 33425 20451
rect 33459 20417 33471 20451
rect 33413 20411 33471 20417
rect 33597 20451 33655 20457
rect 33597 20417 33609 20451
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20380 16267 20383
rect 19242 20380 19248 20392
rect 16255 20352 19248 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 23566 20340 23572 20392
rect 23624 20340 23630 20392
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20380 23811 20383
rect 23934 20380 23940 20392
rect 23799 20352 23940 20380
rect 23799 20349 23811 20352
rect 23753 20343 23811 20349
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 28261 20383 28319 20389
rect 28261 20349 28273 20383
rect 28307 20380 28319 20383
rect 29086 20380 29092 20392
rect 28307 20352 29092 20380
rect 28307 20349 28319 20352
rect 28261 20343 28319 20349
rect 29086 20340 29092 20352
rect 29144 20340 29150 20392
rect 30561 20383 30619 20389
rect 30561 20380 30573 20383
rect 30484 20352 30573 20380
rect 11238 20272 11244 20324
rect 11296 20312 11302 20324
rect 24854 20312 24860 20324
rect 11296 20284 17080 20312
rect 11296 20272 11302 20284
rect 10594 20204 10600 20256
rect 10652 20244 10658 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 10652 20216 10701 20244
rect 10652 20204 10658 20216
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 10689 20207 10747 20213
rect 13078 20204 13084 20256
rect 13136 20204 13142 20256
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 17052 20244 17080 20284
rect 19260 20284 24860 20312
rect 19260 20244 19288 20284
rect 24854 20272 24860 20284
rect 24912 20272 24918 20324
rect 28629 20315 28687 20321
rect 28629 20281 28641 20315
rect 28675 20312 28687 20315
rect 28902 20312 28908 20324
rect 28675 20284 28908 20312
rect 28675 20281 28687 20284
rect 28629 20275 28687 20281
rect 28902 20272 28908 20284
rect 28960 20272 28966 20324
rect 29822 20312 29828 20324
rect 29656 20284 29828 20312
rect 17052 20216 19288 20244
rect 20806 20204 20812 20256
rect 20864 20204 20870 20256
rect 26142 20204 26148 20256
rect 26200 20244 26206 20256
rect 29656 20244 29684 20284
rect 29822 20272 29828 20284
rect 29880 20272 29886 20324
rect 29914 20272 29920 20324
rect 29972 20312 29978 20324
rect 30484 20312 30512 20352
rect 30561 20349 30573 20352
rect 30607 20349 30619 20383
rect 30561 20343 30619 20349
rect 31389 20383 31447 20389
rect 31389 20349 31401 20383
rect 31435 20380 31447 20383
rect 32950 20380 32956 20392
rect 31435 20352 32956 20380
rect 31435 20349 31447 20352
rect 31389 20343 31447 20349
rect 32950 20340 32956 20352
rect 33008 20340 33014 20392
rect 33428 20324 33456 20411
rect 29972 20284 30512 20312
rect 31665 20315 31723 20321
rect 29972 20272 29978 20284
rect 31665 20281 31677 20315
rect 31711 20312 31723 20315
rect 33410 20312 33416 20324
rect 31711 20284 33416 20312
rect 31711 20281 31723 20284
rect 31665 20275 31723 20281
rect 33410 20272 33416 20284
rect 33468 20272 33474 20324
rect 33612 20256 33640 20411
rect 33686 20408 33692 20460
rect 33744 20408 33750 20460
rect 33888 20457 33916 20488
rect 33980 20457 34008 20544
rect 34072 20488 34560 20516
rect 34072 20457 34100 20488
rect 34532 20460 34560 20488
rect 33873 20451 33931 20457
rect 33873 20417 33885 20451
rect 33919 20417 33931 20451
rect 33873 20411 33931 20417
rect 33965 20451 34023 20457
rect 33965 20417 33977 20451
rect 34011 20417 34023 20451
rect 33965 20411 34023 20417
rect 34057 20451 34115 20457
rect 34057 20417 34069 20451
rect 34103 20417 34115 20451
rect 34057 20411 34115 20417
rect 34425 20451 34483 20457
rect 34425 20417 34437 20451
rect 34471 20417 34483 20451
rect 34425 20411 34483 20417
rect 33704 20380 33732 20408
rect 34440 20380 34468 20411
rect 34514 20408 34520 20460
rect 34572 20408 34578 20460
rect 34624 20457 34652 20544
rect 34698 20476 34704 20528
rect 34756 20516 34762 20528
rect 35161 20519 35219 20525
rect 35161 20516 35173 20519
rect 34756 20488 35173 20516
rect 34756 20476 34762 20488
rect 35161 20485 35173 20488
rect 35207 20485 35219 20519
rect 35161 20479 35219 20485
rect 34609 20451 34667 20457
rect 34609 20417 34621 20451
rect 34655 20417 34667 20451
rect 34609 20411 34667 20417
rect 36262 20408 36268 20460
rect 36320 20408 36326 20460
rect 36909 20451 36967 20457
rect 36909 20417 36921 20451
rect 36955 20448 36967 20451
rect 37292 20448 37320 20547
rect 37642 20544 37648 20596
rect 37700 20584 37706 20596
rect 37737 20587 37795 20593
rect 37737 20584 37749 20587
rect 37700 20556 37749 20584
rect 37700 20544 37706 20556
rect 37737 20553 37749 20556
rect 37783 20553 37795 20587
rect 37737 20547 37795 20553
rect 39577 20587 39635 20593
rect 39577 20553 39589 20587
rect 39623 20584 39635 20587
rect 39850 20584 39856 20596
rect 39623 20556 39856 20584
rect 39623 20553 39635 20556
rect 39577 20547 39635 20553
rect 39850 20544 39856 20556
rect 39908 20544 39914 20596
rect 40310 20544 40316 20596
rect 40368 20544 40374 20596
rect 42150 20544 42156 20596
rect 42208 20544 42214 20596
rect 42518 20544 42524 20596
rect 42576 20584 42582 20596
rect 42613 20587 42671 20593
rect 42613 20584 42625 20587
rect 42576 20556 42625 20584
rect 42576 20544 42582 20556
rect 42613 20553 42625 20556
rect 42659 20553 42671 20587
rect 42613 20547 42671 20553
rect 39393 20519 39451 20525
rect 39393 20485 39405 20519
rect 39439 20516 39451 20519
rect 39758 20516 39764 20528
rect 39439 20488 39764 20516
rect 39439 20485 39451 20488
rect 39393 20479 39451 20485
rect 39758 20476 39764 20488
rect 39816 20476 39822 20528
rect 36955 20420 37320 20448
rect 36955 20417 36967 20420
rect 36909 20411 36967 20417
rect 37458 20408 37464 20460
rect 37516 20408 37522 20460
rect 37645 20451 37703 20457
rect 37645 20417 37657 20451
rect 37691 20448 37703 20451
rect 38105 20451 38163 20457
rect 38105 20448 38117 20451
rect 37691 20420 38117 20448
rect 37691 20417 37703 20420
rect 37645 20411 37703 20417
rect 38105 20417 38117 20420
rect 38151 20417 38163 20451
rect 38105 20411 38163 20417
rect 38286 20408 38292 20460
rect 38344 20448 38350 20460
rect 38657 20451 38715 20457
rect 38657 20448 38669 20451
rect 38344 20420 38669 20448
rect 38344 20408 38350 20420
rect 38657 20417 38669 20420
rect 38703 20417 38715 20451
rect 38657 20411 38715 20417
rect 39022 20408 39028 20460
rect 39080 20408 39086 20460
rect 39114 20408 39120 20460
rect 39172 20448 39178 20460
rect 39209 20451 39267 20457
rect 39209 20448 39221 20451
rect 39172 20420 39221 20448
rect 39172 20408 39178 20420
rect 39209 20417 39221 20420
rect 39255 20417 39267 20451
rect 39209 20411 39267 20417
rect 39669 20451 39727 20457
rect 39669 20417 39681 20451
rect 39715 20448 39727 20451
rect 40328 20448 40356 20544
rect 39715 20420 40356 20448
rect 42168 20448 42196 20544
rect 42242 20476 42248 20528
rect 42300 20516 42306 20528
rect 42797 20519 42855 20525
rect 42797 20516 42809 20519
rect 42300 20488 42809 20516
rect 42300 20476 42306 20488
rect 42797 20485 42809 20488
rect 42843 20516 42855 20519
rect 43438 20516 43444 20528
rect 42843 20488 43444 20516
rect 42843 20485 42855 20488
rect 42797 20479 42855 20485
rect 43438 20476 43444 20488
rect 43496 20476 43502 20528
rect 42521 20451 42579 20457
rect 42521 20448 42533 20451
rect 42168 20420 42533 20448
rect 39715 20417 39727 20420
rect 39669 20411 39727 20417
rect 42521 20417 42533 20420
rect 42567 20417 42579 20451
rect 42521 20411 42579 20417
rect 33704 20352 34468 20380
rect 34885 20383 34943 20389
rect 34885 20349 34897 20383
rect 34931 20349 34943 20383
rect 36280 20380 36308 20408
rect 37476 20380 37504 20408
rect 36280 20352 37504 20380
rect 34885 20343 34943 20349
rect 34054 20272 34060 20324
rect 34112 20312 34118 20324
rect 34790 20312 34796 20324
rect 34112 20284 34796 20312
rect 34112 20272 34118 20284
rect 34790 20272 34796 20284
rect 34848 20272 34854 20324
rect 26200 20216 29684 20244
rect 26200 20204 26206 20216
rect 29730 20204 29736 20256
rect 29788 20244 29794 20256
rect 30745 20247 30803 20253
rect 30745 20244 30757 20247
rect 29788 20216 30757 20244
rect 29788 20204 29794 20216
rect 30745 20213 30757 20216
rect 30791 20213 30803 20247
rect 30745 20207 30803 20213
rect 33594 20204 33600 20256
rect 33652 20204 33658 20256
rect 34330 20204 34336 20256
rect 34388 20204 34394 20256
rect 34514 20204 34520 20256
rect 34572 20204 34578 20256
rect 34900 20244 34928 20343
rect 37550 20340 37556 20392
rect 37608 20380 37614 20392
rect 37829 20383 37887 20389
rect 37829 20380 37841 20383
rect 37608 20352 37841 20380
rect 37608 20340 37614 20352
rect 37829 20349 37841 20352
rect 37875 20349 37887 20383
rect 37829 20343 37887 20349
rect 39301 20383 39359 20389
rect 39301 20349 39313 20383
rect 39347 20380 39359 20383
rect 39347 20352 39436 20380
rect 39347 20349 39359 20352
rect 39301 20343 39359 20349
rect 36538 20272 36544 20324
rect 36596 20312 36602 20324
rect 39408 20321 39436 20352
rect 36725 20315 36783 20321
rect 36725 20312 36737 20315
rect 36596 20284 36737 20312
rect 36596 20272 36602 20284
rect 36725 20281 36737 20284
rect 36771 20281 36783 20315
rect 36725 20275 36783 20281
rect 39393 20315 39451 20321
rect 39393 20281 39405 20315
rect 39439 20281 39451 20315
rect 39393 20275 39451 20281
rect 35894 20244 35900 20256
rect 34900 20216 35900 20244
rect 35894 20204 35900 20216
rect 35952 20204 35958 20256
rect 38838 20204 38844 20256
rect 38896 20204 38902 20256
rect 42794 20204 42800 20256
rect 42852 20204 42858 20256
rect 1104 20154 44620 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 44620 20154
rect 1104 20080 44620 20102
rect 10400 20043 10458 20049
rect 10400 20009 10412 20043
rect 10446 20040 10458 20043
rect 10594 20040 10600 20052
rect 10446 20012 10600 20040
rect 10446 20009 10458 20012
rect 10400 20003 10458 20009
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 11974 20040 11980 20052
rect 11931 20012 11980 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 13722 20000 13728 20052
rect 13780 20000 13786 20052
rect 13909 20043 13967 20049
rect 13909 20009 13921 20043
rect 13955 20040 13967 20043
rect 14274 20040 14280 20052
rect 13955 20012 14280 20040
rect 13955 20009 13967 20012
rect 13909 20003 13967 20009
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 15470 20049 15476 20052
rect 15460 20043 15476 20049
rect 15460 20009 15472 20043
rect 15460 20003 15476 20009
rect 15470 20000 15476 20003
rect 15528 20000 15534 20052
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 17310 20040 17316 20052
rect 15896 20012 17316 20040
rect 15896 20000 15902 20012
rect 17310 20000 17316 20012
rect 17368 20040 17374 20052
rect 17497 20043 17555 20049
rect 17497 20040 17509 20043
rect 17368 20012 17509 20040
rect 17368 20000 17374 20012
rect 17497 20009 17509 20012
rect 17543 20009 17555 20043
rect 17497 20003 17555 20009
rect 6181 19975 6239 19981
rect 6181 19941 6193 19975
rect 6227 19972 6239 19975
rect 7190 19972 7196 19984
rect 6227 19944 7196 19972
rect 6227 19941 6239 19944
rect 6181 19935 6239 19941
rect 6288 19768 6316 19944
rect 7190 19932 7196 19944
rect 7248 19972 7254 19984
rect 8110 19972 8116 19984
rect 7248 19944 8116 19972
rect 7248 19932 7254 19944
rect 8110 19932 8116 19944
rect 8168 19932 8174 19984
rect 13740 19972 13768 20000
rect 14093 19975 14151 19981
rect 14093 19972 14105 19975
rect 13740 19944 14105 19972
rect 14093 19941 14105 19944
rect 14139 19941 14151 19975
rect 14093 19935 14151 19941
rect 9490 19864 9496 19916
rect 9548 19904 9554 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9548 19876 10149 19904
rect 9548 19864 9554 19876
rect 10137 19873 10149 19876
rect 10183 19904 10195 19907
rect 11146 19904 11152 19916
rect 10183 19876 11152 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 11146 19864 11152 19876
rect 11204 19904 11210 19916
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 11204 19876 12173 19904
rect 11204 19864 11210 19876
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19904 12495 19907
rect 13078 19904 13084 19916
rect 12483 19876 13084 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 14737 19907 14795 19913
rect 14737 19873 14749 19907
rect 14783 19904 14795 19907
rect 15010 19904 15016 19916
rect 14783 19876 15016 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 17512 19904 17540 20003
rect 18138 20000 18144 20052
rect 18196 20000 18202 20052
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 18564 20012 19257 20040
rect 18564 20000 18570 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 20530 20040 20536 20052
rect 19245 20003 19303 20009
rect 19812 20012 20536 20040
rect 19812 19913 19840 20012
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 22646 20040 22652 20052
rect 20640 20012 22652 20040
rect 20640 19972 20668 20012
rect 22646 20000 22652 20012
rect 22704 20000 22710 20052
rect 25501 20043 25559 20049
rect 25501 20009 25513 20043
rect 25547 20040 25559 20043
rect 28350 20040 28356 20052
rect 25547 20012 28356 20040
rect 25547 20009 25559 20012
rect 25501 20003 25559 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 28626 20000 28632 20052
rect 28684 20000 28690 20052
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 28960 20012 29592 20040
rect 28960 20000 28966 20012
rect 19904 19944 20668 19972
rect 19797 19907 19855 19913
rect 19797 19904 19809 19907
rect 15252 19876 17356 19904
rect 17512 19876 19809 19904
rect 15252 19864 15258 19876
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 7006 19836 7012 19848
rect 6411 19808 7012 19836
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14516 19808 14565 19836
rect 14516 19796 14522 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 6549 19771 6607 19777
rect 6549 19768 6561 19771
rect 6288 19740 6561 19768
rect 6549 19737 6561 19740
rect 6595 19737 6607 19771
rect 6549 19731 6607 19737
rect 6917 19771 6975 19777
rect 6917 19737 6929 19771
rect 6963 19768 6975 19771
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 6963 19740 7389 19768
rect 6963 19737 6975 19740
rect 6917 19731 6975 19737
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 7064 19672 7113 19700
rect 7064 19660 7070 19672
rect 7101 19669 7113 19672
rect 7147 19669 7159 19703
rect 7392 19700 7420 19731
rect 10962 19728 10968 19780
rect 11020 19728 11026 19780
rect 15028 19768 15056 19864
rect 17328 19848 17356 19876
rect 19797 19873 19809 19876
rect 19843 19873 19855 19907
rect 19797 19867 19855 19873
rect 17310 19796 17316 19848
rect 17368 19796 17374 19848
rect 18598 19796 18604 19848
rect 18656 19796 18662 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 19702 19836 19708 19848
rect 19659 19808 19708 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 15746 19768 15752 19780
rect 12544 19740 12926 19768
rect 15028 19740 15752 19768
rect 7834 19700 7840 19712
rect 7392 19672 7840 19700
rect 7101 19663 7159 19669
rect 7834 19660 7840 19672
rect 7892 19700 7898 19712
rect 11146 19700 11152 19712
rect 7892 19672 11152 19700
rect 7892 19660 7898 19672
rect 11146 19660 11152 19672
rect 11204 19700 11210 19712
rect 12544 19700 12572 19740
rect 15746 19728 15752 19740
rect 15804 19728 15810 19780
rect 16758 19768 16764 19780
rect 16698 19740 16764 19768
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 17221 19771 17279 19777
rect 17221 19737 17233 19771
rect 17267 19737 17279 19771
rect 17221 19731 17279 19737
rect 11204 19672 12572 19700
rect 14461 19703 14519 19709
rect 11204 19660 11210 19672
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 14550 19700 14556 19712
rect 14507 19672 14556 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 16206 19660 16212 19712
rect 16264 19700 16270 19712
rect 17236 19700 17264 19731
rect 17402 19728 17408 19780
rect 17460 19768 17466 19780
rect 18233 19771 18291 19777
rect 18233 19768 18245 19771
rect 17460 19740 18245 19768
rect 17460 19728 17466 19740
rect 18233 19737 18245 19740
rect 18279 19768 18291 19771
rect 18506 19768 18512 19780
rect 18279 19740 18512 19768
rect 18279 19737 18291 19740
rect 18233 19731 18291 19737
rect 18506 19728 18512 19740
rect 18564 19728 18570 19780
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 19904 19768 19932 19944
rect 21910 19932 21916 19984
rect 21968 19972 21974 19984
rect 25774 19972 25780 19984
rect 21968 19944 25780 19972
rect 21968 19932 21974 19944
rect 25774 19932 25780 19944
rect 25832 19932 25838 19984
rect 26326 19972 26332 19984
rect 25884 19944 26332 19972
rect 22462 19904 22468 19916
rect 20548 19876 22468 19904
rect 20548 19845 20576 19876
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 25225 19907 25283 19913
rect 25225 19873 25237 19907
rect 25271 19873 25283 19907
rect 25884 19904 25912 19944
rect 26326 19932 26332 19944
rect 26384 19932 26390 19984
rect 28644 19972 28672 20000
rect 29181 19975 29239 19981
rect 29181 19972 29193 19975
rect 27908 19944 29193 19972
rect 25225 19867 25283 19873
rect 25792 19876 25912 19904
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 19300 19740 19932 19768
rect 20548 19768 20576 19799
rect 24854 19796 24860 19848
rect 24912 19836 24918 19848
rect 25133 19839 25191 19845
rect 25133 19836 25145 19839
rect 24912 19808 25145 19836
rect 24912 19796 24918 19808
rect 25133 19805 25145 19808
rect 25179 19805 25191 19839
rect 25240 19836 25268 19867
rect 25593 19839 25651 19845
rect 25593 19836 25605 19839
rect 25240 19808 25605 19836
rect 25133 19799 25191 19805
rect 25593 19805 25605 19808
rect 25639 19805 25651 19839
rect 25593 19799 25651 19805
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 25792 19845 25820 19876
rect 26050 19864 26056 19916
rect 26108 19864 26114 19916
rect 27908 19913 27936 19944
rect 29181 19941 29193 19944
rect 29227 19941 29239 19975
rect 29181 19935 29239 19941
rect 29362 19932 29368 19984
rect 29420 19932 29426 19984
rect 27893 19907 27951 19913
rect 27893 19873 27905 19907
rect 27939 19873 27951 19907
rect 27893 19867 27951 19873
rect 28258 19864 28264 19916
rect 28316 19864 28322 19916
rect 28629 19907 28687 19913
rect 28629 19873 28641 19907
rect 28675 19904 28687 19907
rect 29380 19904 29408 19932
rect 29564 19913 29592 20012
rect 30006 20000 30012 20052
rect 30064 20000 30070 20052
rect 30098 20000 30104 20052
rect 30156 20040 30162 20052
rect 30193 20043 30251 20049
rect 30193 20040 30205 20043
rect 30156 20012 30205 20040
rect 30156 20000 30162 20012
rect 30193 20009 30205 20012
rect 30239 20009 30251 20043
rect 30193 20003 30251 20009
rect 31018 20000 31024 20052
rect 31076 20000 31082 20052
rect 33410 20000 33416 20052
rect 33468 20000 33474 20052
rect 36630 20040 36636 20052
rect 34164 20012 36636 20040
rect 29914 19932 29920 19984
rect 29972 19932 29978 19984
rect 28675 19876 29408 19904
rect 29549 19907 29607 19913
rect 28675 19873 28687 19876
rect 28629 19867 28687 19873
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25740 19808 25789 19836
rect 25740 19796 25746 19808
rect 25777 19805 25789 19808
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 25866 19796 25872 19848
rect 25924 19836 25930 19848
rect 25961 19839 26019 19845
rect 25961 19836 25973 19839
rect 25924 19808 25973 19836
rect 25924 19796 25930 19808
rect 25961 19805 25973 19808
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19836 28043 19839
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28031 19808 28457 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28721 19839 28779 19845
rect 28721 19805 28733 19839
rect 28767 19836 28779 19839
rect 28994 19836 29000 19848
rect 28767 19808 29000 19836
rect 28767 19805 28779 19808
rect 28721 19799 28779 19805
rect 28994 19796 29000 19808
rect 29052 19836 29058 19848
rect 29196 19845 29224 19876
rect 29549 19873 29561 19907
rect 29595 19904 29607 19907
rect 29730 19904 29736 19916
rect 29595 19876 29736 19904
rect 29595 19873 29607 19876
rect 29549 19867 29607 19873
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 29181 19839 29239 19845
rect 29052 19808 29132 19836
rect 29052 19796 29058 19808
rect 20548 19740 20668 19768
rect 19300 19728 19306 19740
rect 20640 19712 20668 19740
rect 20806 19728 20812 19780
rect 20864 19728 20870 19780
rect 22370 19768 22376 19780
rect 22034 19740 22376 19768
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 26142 19728 26148 19780
rect 26200 19728 26206 19780
rect 28353 19771 28411 19777
rect 28353 19737 28365 19771
rect 28399 19768 28411 19771
rect 28810 19768 28816 19780
rect 28399 19740 28816 19768
rect 28399 19737 28411 19740
rect 28353 19731 28411 19737
rect 28810 19728 28816 19740
rect 28868 19728 28874 19780
rect 29104 19768 29132 19808
rect 29181 19805 29193 19839
rect 29227 19805 29239 19839
rect 29181 19799 29239 19805
rect 29365 19839 29423 19845
rect 29365 19805 29377 19839
rect 29411 19805 29423 19839
rect 30024 19836 30052 20000
rect 31570 19864 31576 19916
rect 31628 19904 31634 19916
rect 32306 19904 32312 19916
rect 31628 19876 32312 19904
rect 31628 19864 31634 19876
rect 32306 19864 32312 19876
rect 32364 19864 32370 19916
rect 33428 19904 33456 20000
rect 33428 19876 33732 19904
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 30024 19808 30113 19836
rect 29365 19799 29423 19805
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 31113 19839 31171 19845
rect 31113 19805 31125 19839
rect 31159 19836 31171 19839
rect 31754 19836 31760 19848
rect 31159 19808 31760 19836
rect 31159 19805 31171 19808
rect 31113 19799 31171 19805
rect 31726 19802 31760 19808
rect 29380 19768 29408 19799
rect 31754 19796 31760 19802
rect 31812 19796 31818 19848
rect 31864 19808 32076 19836
rect 30006 19768 30012 19780
rect 29104 19740 30012 19768
rect 30006 19728 30012 19740
rect 30064 19728 30070 19780
rect 31864 19768 31892 19808
rect 32048 19777 32076 19808
rect 33594 19796 33600 19848
rect 33652 19796 33658 19848
rect 33704 19845 33732 19876
rect 34164 19845 34192 20012
rect 36630 20000 36636 20012
rect 36688 20000 36694 20052
rect 37921 20043 37979 20049
rect 37921 20009 37933 20043
rect 37967 20040 37979 20043
rect 38286 20040 38292 20052
rect 37967 20012 38292 20040
rect 37967 20009 37979 20012
rect 37921 20003 37979 20009
rect 38286 20000 38292 20012
rect 38344 20000 38350 20052
rect 38841 20043 38899 20049
rect 38841 20009 38853 20043
rect 38887 20040 38899 20043
rect 38930 20040 38936 20052
rect 38887 20012 38936 20040
rect 38887 20009 38899 20012
rect 38841 20003 38899 20009
rect 38930 20000 38936 20012
rect 38988 20000 38994 20052
rect 39390 19932 39396 19984
rect 39448 19932 39454 19984
rect 36449 19907 36507 19913
rect 36449 19873 36461 19907
rect 36495 19904 36507 19907
rect 36538 19904 36544 19916
rect 36495 19876 36544 19904
rect 36495 19873 36507 19876
rect 36449 19867 36507 19873
rect 36538 19864 36544 19876
rect 36596 19864 36602 19916
rect 38562 19864 38568 19916
rect 38620 19864 38626 19916
rect 33689 19839 33747 19845
rect 33689 19805 33701 19839
rect 33735 19836 33747 19839
rect 33965 19839 34023 19845
rect 33965 19836 33977 19839
rect 33735 19808 33977 19836
rect 33735 19805 33747 19808
rect 33689 19799 33747 19805
rect 33965 19805 33977 19808
rect 34011 19805 34023 19839
rect 33965 19799 34023 19805
rect 34149 19839 34207 19845
rect 34149 19805 34161 19839
rect 34195 19805 34207 19839
rect 34149 19799 34207 19805
rect 31496 19740 31892 19768
rect 32033 19771 32091 19777
rect 16264 19672 17264 19700
rect 16264 19660 16270 19672
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 20438 19700 20444 19712
rect 19751 19672 20444 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 22281 19703 22339 19709
rect 22281 19700 22293 19703
rect 21232 19672 22293 19700
rect 21232 19660 21238 19672
rect 22281 19669 22293 19672
rect 22327 19700 22339 19703
rect 26160 19700 26188 19728
rect 22327 19672 26188 19700
rect 22327 19669 22339 19672
rect 22281 19663 22339 19669
rect 27706 19660 27712 19712
rect 27764 19660 27770 19712
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 28994 19700 29000 19712
rect 27856 19672 29000 19700
rect 27856 19660 27862 19672
rect 28994 19660 29000 19672
rect 29052 19660 29058 19712
rect 29089 19703 29147 19709
rect 29089 19669 29101 19703
rect 29135 19700 29147 19703
rect 29178 19700 29184 19712
rect 29135 19672 29184 19700
rect 29135 19669 29147 19672
rect 29089 19663 29147 19669
rect 29178 19660 29184 19672
rect 29236 19700 29242 19712
rect 31496 19700 31524 19740
rect 32033 19737 32045 19771
rect 32079 19737 32091 19771
rect 33612 19768 33640 19796
rect 34164 19768 34192 19799
rect 35986 19796 35992 19848
rect 36044 19836 36050 19848
rect 36173 19839 36231 19845
rect 36173 19836 36185 19839
rect 36044 19808 36185 19836
rect 36044 19796 36050 19808
rect 36173 19805 36185 19808
rect 36219 19805 36231 19839
rect 36173 19799 36231 19805
rect 38749 19839 38807 19845
rect 38749 19805 38761 19839
rect 38795 19805 38807 19839
rect 38749 19799 38807 19805
rect 38933 19839 38991 19845
rect 38933 19805 38945 19839
rect 38979 19836 38991 19839
rect 39408 19836 39436 19932
rect 39945 19839 40003 19845
rect 39945 19836 39957 19839
rect 38979 19808 39957 19836
rect 38979 19805 38991 19808
rect 38933 19799 38991 19805
rect 39945 19805 39957 19808
rect 39991 19805 40003 19839
rect 39945 19799 40003 19805
rect 33612 19740 34192 19768
rect 32033 19731 32091 19737
rect 29236 19672 31524 19700
rect 32048 19700 32076 19731
rect 37458 19728 37464 19780
rect 37516 19728 37522 19780
rect 38764 19768 38792 19799
rect 40126 19796 40132 19848
rect 40184 19796 40190 19848
rect 40405 19839 40463 19845
rect 40405 19805 40417 19839
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 42889 19839 42947 19845
rect 42889 19805 42901 19839
rect 42935 19836 42947 19839
rect 42978 19836 42984 19848
rect 42935 19808 42984 19836
rect 42935 19805 42947 19808
rect 42889 19799 42947 19805
rect 39025 19771 39083 19777
rect 39025 19768 39037 19771
rect 38764 19740 39037 19768
rect 39025 19737 39037 19740
rect 39071 19768 39083 19771
rect 39758 19768 39764 19780
rect 39071 19740 39764 19768
rect 39071 19737 39083 19740
rect 39025 19731 39083 19737
rect 39758 19728 39764 19740
rect 39816 19768 39822 19780
rect 40420 19768 40448 19799
rect 42978 19796 42984 19808
rect 43036 19796 43042 19848
rect 39816 19740 40448 19768
rect 42705 19771 42763 19777
rect 39816 19728 39822 19740
rect 42705 19737 42717 19771
rect 42751 19768 42763 19771
rect 43438 19768 43444 19780
rect 42751 19740 43444 19768
rect 42751 19737 42763 19740
rect 42705 19731 42763 19737
rect 43438 19728 43444 19740
rect 43496 19728 43502 19780
rect 33778 19700 33784 19712
rect 32048 19672 33784 19700
rect 29236 19660 29242 19672
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 33870 19660 33876 19712
rect 33928 19660 33934 19712
rect 34057 19703 34115 19709
rect 34057 19669 34069 19703
rect 34103 19700 34115 19703
rect 34422 19700 34428 19712
rect 34103 19672 34428 19700
rect 34103 19669 34115 19672
rect 34057 19663 34115 19669
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 38010 19660 38016 19712
rect 38068 19660 38074 19712
rect 39482 19660 39488 19712
rect 39540 19660 39546 19712
rect 42518 19660 42524 19712
rect 42576 19660 42582 19712
rect 1104 19610 44620 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 44620 19610
rect 1104 19536 44620 19558
rect 6914 19496 6920 19508
rect 2884 19468 6920 19496
rect 2884 19369 2912 19468
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 11238 19456 11244 19508
rect 11296 19456 11302 19508
rect 14734 19496 14740 19508
rect 13464 19468 14740 19496
rect 13464 19440 13492 19468
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 15194 19456 15200 19508
rect 15252 19456 15258 19508
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 16080 19468 16681 19496
rect 16080 19456 16086 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 20901 19499 20959 19505
rect 16816 19468 19288 19496
rect 16816 19456 16822 19468
rect 7006 19428 7012 19440
rect 4370 19400 7012 19428
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 11606 19388 11612 19440
rect 11664 19428 11670 19440
rect 12066 19428 12072 19440
rect 11664 19400 12072 19428
rect 11664 19388 11670 19400
rect 12066 19388 12072 19400
rect 12124 19428 12130 19440
rect 13446 19428 13452 19440
rect 12124 19400 13452 19428
rect 12124 19388 12130 19400
rect 13446 19388 13452 19400
rect 13504 19388 13510 19440
rect 15212 19428 15240 19456
rect 16776 19428 16804 19456
rect 14752 19400 15240 19428
rect 16238 19400 16804 19428
rect 18141 19431 18199 19437
rect 2869 19363 2927 19369
rect 2869 19329 2881 19363
rect 2915 19329 2927 19363
rect 7285 19363 7343 19369
rect 2869 19323 2927 19329
rect 4632 19332 6684 19360
rect 3142 19252 3148 19304
rect 3200 19252 3206 19304
rect 4632 19301 4660 19332
rect 6656 19301 6684 19332
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 8478 19360 8484 19372
rect 7331 19332 8484 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 11054 19360 11060 19372
rect 10902 19332 11060 19360
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 14642 19360 14648 19372
rect 13219 19332 14648 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 14752 19369 14780 19400
rect 18141 19397 18153 19431
rect 18187 19428 18199 19431
rect 18414 19428 18420 19440
rect 18187 19400 18420 19428
rect 18187 19397 18199 19400
rect 18141 19391 18199 19397
rect 18414 19388 18420 19400
rect 18472 19388 18478 19440
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 17310 19320 17316 19372
rect 17368 19360 17374 19372
rect 17862 19360 17868 19372
rect 17368 19332 17868 19360
rect 17368 19320 17374 19332
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 19260 19360 19288 19468
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20990 19496 20996 19508
rect 20947 19468 20996 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 21232 19468 21281 19496
rect 21232 19456 21238 19468
rect 21269 19465 21281 19468
rect 21315 19465 21327 19499
rect 21269 19459 21327 19465
rect 22462 19456 22468 19508
rect 22520 19496 22526 19508
rect 23750 19496 23756 19508
rect 22520 19468 23756 19496
rect 22520 19456 22526 19468
rect 23750 19456 23756 19468
rect 23808 19456 23814 19508
rect 26142 19456 26148 19508
rect 26200 19456 26206 19508
rect 28258 19456 28264 19508
rect 28316 19496 28322 19508
rect 28721 19499 28779 19505
rect 28316 19468 28580 19496
rect 28316 19456 28322 19468
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 19886 19428 19892 19440
rect 19484 19400 19892 19428
rect 19484 19388 19490 19400
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 22370 19428 22376 19440
rect 19996 19400 22376 19428
rect 19996 19360 20024 19400
rect 22370 19388 22376 19400
rect 22428 19428 22434 19440
rect 24581 19431 24639 19437
rect 22428 19400 23322 19428
rect 22428 19388 22434 19400
rect 24581 19397 24593 19431
rect 24627 19428 24639 19431
rect 25685 19431 25743 19437
rect 25685 19428 25697 19431
rect 24627 19400 25697 19428
rect 24627 19397 24639 19400
rect 24581 19391 24639 19397
rect 25685 19397 25697 19400
rect 25731 19428 25743 19431
rect 25774 19428 25780 19440
rect 25731 19400 25780 19428
rect 25731 19397 25743 19400
rect 25685 19391 25743 19397
rect 25774 19388 25780 19400
rect 25832 19388 25838 19440
rect 19260 19346 20024 19360
rect 19274 19332 20024 19346
rect 21358 19320 21364 19372
rect 21416 19320 21422 19372
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 22520 19332 22569 19360
rect 22520 19320 22526 19332
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 25498 19320 25504 19372
rect 25556 19360 25562 19372
rect 25869 19363 25927 19369
rect 25869 19360 25881 19363
rect 25556 19332 25881 19360
rect 25556 19320 25562 19332
rect 25869 19329 25881 19332
rect 25915 19329 25927 19363
rect 25869 19323 25927 19329
rect 25961 19363 26019 19369
rect 25961 19329 25973 19363
rect 26007 19360 26019 19363
rect 26160 19360 26188 19456
rect 27798 19388 27804 19440
rect 27856 19388 27862 19440
rect 26007 19332 26188 19360
rect 26007 19329 26019 19332
rect 25961 19323 26019 19329
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26292 19332 26985 19360
rect 26292 19320 26298 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 28552 19360 28580 19468
rect 28721 19465 28733 19499
rect 28767 19465 28779 19499
rect 28721 19459 28779 19465
rect 28736 19428 28764 19459
rect 28810 19456 28816 19508
rect 28868 19456 28874 19508
rect 29086 19456 29092 19508
rect 29144 19456 29150 19508
rect 29914 19456 29920 19508
rect 29972 19456 29978 19508
rect 32030 19496 32036 19508
rect 31312 19468 32036 19496
rect 29104 19428 29132 19456
rect 29733 19431 29791 19437
rect 29733 19428 29745 19431
rect 28736 19400 29745 19428
rect 29380 19369 29408 19400
rect 29733 19397 29745 19400
rect 29779 19397 29791 19431
rect 29733 19391 29791 19397
rect 29365 19363 29423 19369
rect 28552 19332 29316 19360
rect 26973 19323 27031 19329
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 7926 19252 7932 19304
rect 7984 19252 7990 19304
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19292 9827 19295
rect 10134 19292 10140 19304
rect 9815 19264 10140 19292
rect 9815 19261 9827 19264
rect 9769 19255 9827 19261
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 15010 19252 15016 19304
rect 15068 19252 15074 19304
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16531 19264 17233 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 21545 19295 21603 19301
rect 21545 19292 21557 19295
rect 17221 19255 17279 19261
rect 21468 19264 21557 19292
rect 21468 19236 21496 19264
rect 21545 19261 21557 19264
rect 21591 19261 21603 19295
rect 22833 19295 22891 19301
rect 22833 19292 22845 19295
rect 21545 19255 21603 19261
rect 22388 19264 22845 19292
rect 21450 19184 21456 19236
rect 21508 19184 21514 19236
rect 22388 19233 22416 19264
rect 22833 19261 22845 19264
rect 22879 19261 22891 19295
rect 22833 19255 22891 19261
rect 27249 19295 27307 19301
rect 27249 19261 27261 19295
rect 27295 19292 27307 19295
rect 27706 19292 27712 19304
rect 27295 19264 27712 19292
rect 27295 19261 27307 19264
rect 27249 19255 27307 19261
rect 27706 19252 27712 19264
rect 27764 19252 27770 19304
rect 29288 19292 29316 19332
rect 29365 19329 29377 19363
rect 29411 19329 29423 19363
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 29365 19323 29423 19329
rect 29472 19332 29561 19360
rect 29472 19292 29500 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 30374 19320 30380 19372
rect 30432 19360 30438 19372
rect 31312 19369 31340 19468
rect 32030 19456 32036 19468
rect 32088 19456 32094 19508
rect 33870 19456 33876 19508
rect 33928 19456 33934 19508
rect 34514 19456 34520 19508
rect 34572 19456 34578 19508
rect 39482 19456 39488 19508
rect 39540 19456 39546 19508
rect 39574 19456 39580 19508
rect 39632 19496 39638 19508
rect 39669 19499 39727 19505
rect 39669 19496 39681 19499
rect 39632 19468 39681 19496
rect 39632 19456 39638 19468
rect 39669 19465 39681 19468
rect 39715 19465 39727 19499
rect 39669 19459 39727 19465
rect 42518 19456 42524 19508
rect 42576 19496 42582 19508
rect 42576 19468 42656 19496
rect 42576 19456 42582 19468
rect 31389 19431 31447 19437
rect 31389 19397 31401 19431
rect 31435 19428 31447 19431
rect 32125 19431 32183 19437
rect 32125 19428 32137 19431
rect 31435 19400 32137 19428
rect 31435 19397 31447 19400
rect 31389 19391 31447 19397
rect 32125 19397 32137 19400
rect 32171 19397 32183 19431
rect 33888 19428 33916 19456
rect 34532 19428 34560 19456
rect 33888 19400 34284 19428
rect 32125 19391 32183 19397
rect 31297 19363 31355 19369
rect 31297 19360 31309 19363
rect 30432 19332 31309 19360
rect 30432 19320 30438 19332
rect 31297 19329 31309 19332
rect 31343 19329 31355 19363
rect 31297 19323 31355 19329
rect 31481 19363 31539 19369
rect 31481 19329 31493 19363
rect 31527 19360 31539 19363
rect 31570 19360 31576 19372
rect 31527 19332 31576 19360
rect 31527 19329 31539 19332
rect 31481 19323 31539 19329
rect 31570 19320 31576 19332
rect 31628 19320 31634 19372
rect 31662 19320 31668 19372
rect 31720 19320 31726 19372
rect 31754 19320 31760 19372
rect 31812 19360 31818 19372
rect 32582 19360 32588 19372
rect 31812 19332 32588 19360
rect 31812 19320 31818 19332
rect 32582 19320 32588 19332
rect 32640 19360 32646 19372
rect 32677 19363 32735 19369
rect 32677 19360 32689 19363
rect 32640 19332 32689 19360
rect 32640 19320 32646 19332
rect 32677 19329 32689 19332
rect 32723 19329 32735 19363
rect 32677 19323 32735 19329
rect 33778 19320 33784 19372
rect 33836 19360 33842 19372
rect 34256 19369 34284 19400
rect 34348 19400 34744 19428
rect 33873 19363 33931 19369
rect 33873 19360 33885 19363
rect 33836 19332 33885 19360
rect 33836 19320 33842 19332
rect 33873 19329 33885 19332
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19329 34299 19363
rect 34241 19323 34299 19329
rect 29288 19264 29500 19292
rect 34149 19295 34207 19301
rect 34149 19261 34161 19295
rect 34195 19292 34207 19295
rect 34348 19292 34376 19400
rect 34422 19320 34428 19372
rect 34480 19320 34486 19372
rect 34716 19369 34744 19400
rect 39500 19369 39528 19456
rect 42628 19437 42656 19468
rect 42794 19456 42800 19508
rect 42852 19456 42858 19508
rect 42613 19431 42671 19437
rect 42613 19397 42625 19431
rect 42659 19397 42671 19431
rect 42812 19428 42840 19456
rect 42812 19400 43576 19428
rect 42613 19391 42671 19397
rect 34517 19363 34575 19369
rect 34517 19329 34529 19363
rect 34563 19329 34575 19363
rect 34517 19323 34575 19329
rect 34701 19363 34759 19369
rect 34701 19329 34713 19363
rect 34747 19329 34759 19363
rect 34701 19323 34759 19329
rect 39485 19363 39543 19369
rect 39485 19329 39497 19363
rect 39531 19329 39543 19363
rect 39485 19323 39543 19329
rect 42429 19363 42487 19369
rect 42429 19329 42441 19363
rect 42475 19360 42487 19363
rect 42475 19332 42656 19360
rect 42475 19329 42487 19332
rect 42429 19323 42487 19329
rect 34532 19292 34560 19323
rect 34195 19264 34376 19292
rect 34440 19264 34560 19292
rect 42628 19292 42656 19332
rect 42702 19320 42708 19372
rect 42760 19320 42766 19372
rect 42797 19363 42855 19369
rect 42797 19329 42809 19363
rect 42843 19360 42855 19363
rect 42886 19360 42892 19372
rect 42843 19332 42892 19360
rect 42843 19329 42855 19332
rect 42797 19323 42855 19329
rect 42886 19320 42892 19332
rect 42944 19320 42950 19372
rect 42978 19320 42984 19372
rect 43036 19360 43042 19372
rect 43257 19363 43315 19369
rect 43257 19360 43269 19363
rect 43036 19332 43269 19360
rect 43036 19320 43042 19332
rect 43257 19329 43269 19332
rect 43303 19329 43315 19363
rect 43257 19323 43315 19329
rect 43349 19363 43407 19369
rect 43349 19329 43361 19363
rect 43395 19360 43407 19363
rect 43438 19360 43444 19372
rect 43395 19332 43444 19360
rect 43395 19329 43407 19332
rect 43349 19323 43407 19329
rect 43438 19320 43444 19332
rect 43496 19320 43502 19372
rect 43548 19369 43576 19400
rect 43533 19363 43591 19369
rect 43533 19329 43545 19363
rect 43579 19329 43591 19363
rect 43533 19323 43591 19329
rect 43622 19320 43628 19372
rect 43680 19320 43686 19372
rect 43073 19295 43131 19301
rect 43073 19292 43085 19295
rect 42628 19264 43085 19292
rect 34195 19261 34207 19264
rect 34149 19255 34207 19261
rect 22373 19227 22431 19233
rect 22373 19193 22385 19227
rect 22419 19193 22431 19227
rect 31846 19224 31852 19236
rect 22373 19187 22431 19193
rect 25976 19196 26280 19224
rect 7374 19116 7380 19168
rect 7432 19116 7438 19168
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17862 19156 17868 19168
rect 17184 19128 17868 19156
rect 17184 19116 17190 19128
rect 17862 19116 17868 19128
rect 17920 19156 17926 19168
rect 25976 19165 26004 19196
rect 25961 19159 26019 19165
rect 25961 19156 25973 19159
rect 17920 19128 25973 19156
rect 17920 19116 17926 19128
rect 25961 19125 25973 19128
rect 26007 19125 26019 19159
rect 25961 19119 26019 19125
rect 26142 19116 26148 19168
rect 26200 19116 26206 19168
rect 26252 19156 26280 19196
rect 28276 19196 31852 19224
rect 28276 19156 28304 19196
rect 31846 19184 31852 19196
rect 31904 19184 31910 19236
rect 34440 19233 34468 19264
rect 43073 19261 43085 19264
rect 43119 19261 43131 19295
rect 43073 19255 43131 19261
rect 34057 19227 34115 19233
rect 34057 19193 34069 19227
rect 34103 19224 34115 19227
rect 34425 19227 34483 19233
rect 34425 19224 34437 19227
rect 34103 19196 34437 19224
rect 34103 19193 34115 19196
rect 34057 19187 34115 19193
rect 34425 19193 34437 19196
rect 34471 19193 34483 19227
rect 34425 19187 34483 19193
rect 26252 19128 28304 19156
rect 31110 19116 31116 19168
rect 31168 19116 31174 19168
rect 33686 19116 33692 19168
rect 33744 19116 33750 19168
rect 34609 19159 34667 19165
rect 34609 19125 34621 19159
rect 34655 19156 34667 19159
rect 35802 19156 35808 19168
rect 34655 19128 35808 19156
rect 34655 19125 34667 19128
rect 34609 19119 34667 19125
rect 35802 19116 35808 19128
rect 35860 19116 35866 19168
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 38194 19156 38200 19168
rect 37884 19128 38200 19156
rect 37884 19116 37890 19128
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 42978 19116 42984 19168
rect 43036 19116 43042 19168
rect 1104 19066 44620 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 44620 19066
rect 1104 18992 44620 19014
rect 6503 18955 6561 18961
rect 6503 18921 6515 18955
rect 6549 18952 6561 18955
rect 7926 18952 7932 18964
rect 6549 18924 7932 18952
rect 6549 18921 6561 18924
rect 6503 18915 6561 18921
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 9490 18912 9496 18964
rect 9548 18912 9554 18964
rect 10870 18912 10876 18964
rect 10928 18912 10934 18964
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 15068 18924 15301 18952
rect 15068 18912 15074 18924
rect 15289 18921 15301 18924
rect 15335 18921 15347 18955
rect 15289 18915 15347 18921
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 18656 18924 19257 18952
rect 18656 18912 18662 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 19245 18915 19303 18921
rect 22186 18912 22192 18964
rect 22244 18952 22250 18964
rect 22373 18955 22431 18961
rect 22373 18952 22385 18955
rect 22244 18924 22385 18952
rect 22244 18912 22250 18924
rect 22373 18921 22385 18924
rect 22419 18921 22431 18955
rect 22373 18915 22431 18921
rect 23750 18912 23756 18964
rect 23808 18912 23814 18964
rect 25866 18912 25872 18964
rect 25924 18912 25930 18964
rect 26326 18912 26332 18964
rect 26384 18912 26390 18964
rect 28966 18924 32536 18952
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 2041 18887 2099 18893
rect 2041 18884 2053 18887
rect 1627 18856 2053 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 2041 18853 2053 18856
rect 2087 18853 2099 18887
rect 2041 18847 2099 18853
rect 1762 18776 1768 18828
rect 1820 18776 1826 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 8352 18788 8493 18816
rect 8352 18776 8358 18788
rect 8481 18785 8493 18788
rect 8527 18816 8539 18819
rect 9508 18816 9536 18912
rect 10778 18844 10784 18896
rect 10836 18884 10842 18896
rect 28966 18884 28994 18924
rect 10836 18856 17448 18884
rect 10836 18844 10842 18856
rect 8527 18788 9536 18816
rect 10321 18819 10379 18825
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 10321 18785 10333 18819
rect 10367 18816 10379 18819
rect 11606 18816 11612 18828
rect 10367 18788 11612 18816
rect 10367 18785 10379 18788
rect 10321 18779 10379 18785
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 14700 18788 15692 18816
rect 14700 18776 14706 18788
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4672 18720 4721 18748
rect 4672 18708 4678 18720
rect 4709 18717 4721 18720
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5074 18708 5080 18760
rect 5132 18708 5138 18760
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8159 18720 8953 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 9272 18720 9505 18748
rect 9272 18708 9278 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10744 18720 10977 18748
rect 10744 18708 10750 18720
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 12986 18708 12992 18760
rect 13044 18708 13050 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 15519 18720 15608 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 10413 18683 10471 18689
rect 5368 18652 5474 18680
rect 7774 18652 7880 18680
rect 2222 18572 2228 18624
rect 2280 18572 2286 18624
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 5368 18612 5396 18652
rect 7852 18624 7880 18652
rect 10413 18649 10425 18683
rect 10459 18680 10471 18683
rect 11882 18680 11888 18692
rect 10459 18652 11888 18680
rect 10459 18649 10471 18652
rect 10413 18643 10471 18649
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 4764 18584 5396 18612
rect 6687 18615 6745 18621
rect 4764 18572 4770 18584
rect 6687 18581 6699 18615
rect 6733 18612 6745 18615
rect 7650 18612 7656 18624
rect 6733 18584 7656 18612
rect 6733 18581 6745 18584
rect 6687 18575 6745 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 11238 18612 11244 18624
rect 10551 18584 11244 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 12434 18572 12440 18624
rect 12492 18572 12498 18624
rect 12802 18572 12808 18624
rect 12860 18572 12866 18624
rect 15580 18621 15608 18720
rect 15664 18680 15692 18788
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16117 18819 16175 18825
rect 16117 18816 16129 18819
rect 15804 18788 16129 18816
rect 15804 18776 15810 18788
rect 16117 18785 16129 18788
rect 16163 18785 16175 18819
rect 16117 18779 16175 18785
rect 17310 18776 17316 18828
rect 17368 18776 17374 18828
rect 17420 18816 17448 18856
rect 18616 18856 28994 18884
rect 32508 18884 32536 18924
rect 32582 18912 32588 18964
rect 32640 18912 32646 18964
rect 33686 18912 33692 18964
rect 33744 18912 33750 18964
rect 42334 18912 42340 18964
rect 42392 18912 42398 18964
rect 42886 18912 42892 18964
rect 42944 18912 42950 18964
rect 43346 18912 43352 18964
rect 43404 18912 43410 18964
rect 32858 18884 32864 18896
rect 32508 18856 32864 18884
rect 18616 18816 18644 18856
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 17420 18788 18644 18816
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16022 18748 16028 18760
rect 15979 18720 16028 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18717 16451 18751
rect 19076 18748 19104 18779
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19392 18788 19809 18816
rect 19392 18776 19398 18788
rect 19797 18785 19809 18788
rect 19843 18816 19855 18819
rect 21450 18816 21456 18828
rect 19843 18788 21456 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 21450 18776 21456 18788
rect 21508 18816 21514 18828
rect 21729 18819 21787 18825
rect 21729 18816 21741 18819
rect 21508 18788 21741 18816
rect 21508 18776 21514 18788
rect 21729 18785 21741 18788
rect 21775 18816 21787 18819
rect 23474 18816 23480 18828
rect 21775 18788 23480 18816
rect 21775 18785 21787 18788
rect 21729 18779 21787 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 25792 18788 26096 18816
rect 25792 18760 25820 18788
rect 20717 18751 20775 18757
rect 20717 18748 20729 18751
rect 19076 18720 20729 18748
rect 16393 18711 16451 18717
rect 20717 18717 20729 18720
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 16408 18680 16436 18711
rect 21910 18708 21916 18760
rect 21968 18748 21974 18760
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21968 18720 22017 18748
rect 21968 18708 21974 18720
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 23106 18708 23112 18760
rect 23164 18748 23170 18760
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23164 18720 24409 18748
rect 23164 18708 23170 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 25774 18708 25780 18760
rect 25832 18708 25838 18760
rect 25866 18708 25872 18760
rect 25924 18708 25930 18760
rect 26068 18757 26096 18788
rect 30834 18776 30840 18828
rect 30892 18776 30898 18828
rect 31110 18776 31116 18828
rect 31168 18776 31174 18828
rect 33704 18816 33732 18912
rect 35437 18887 35495 18893
rect 35437 18853 35449 18887
rect 35483 18884 35495 18887
rect 35710 18884 35716 18896
rect 35483 18856 35716 18884
rect 35483 18853 35495 18856
rect 35437 18847 35495 18853
rect 35710 18844 35716 18856
rect 35768 18844 35774 18896
rect 38194 18844 38200 18896
rect 38252 18884 38258 18896
rect 38930 18884 38936 18896
rect 38252 18856 38936 18884
rect 38252 18844 38258 18856
rect 38930 18844 38936 18856
rect 38988 18844 38994 18896
rect 37461 18819 37519 18825
rect 33704 18788 36032 18816
rect 26053 18751 26111 18757
rect 26053 18717 26065 18751
rect 26099 18717 26111 18751
rect 26053 18711 26111 18717
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 34698 18708 34704 18760
rect 34756 18708 34762 18760
rect 35434 18708 35440 18760
rect 35492 18748 35498 18760
rect 35621 18751 35679 18757
rect 35621 18748 35633 18751
rect 35492 18720 35633 18748
rect 35492 18708 35498 18720
rect 35621 18717 35633 18720
rect 35667 18717 35679 18751
rect 35621 18711 35679 18717
rect 35802 18708 35808 18760
rect 35860 18708 35866 18760
rect 36004 18757 36032 18788
rect 37461 18785 37473 18819
rect 37507 18816 37519 18819
rect 37507 18788 37872 18816
rect 37507 18785 37519 18788
rect 37461 18779 37519 18785
rect 35989 18751 36047 18757
rect 35989 18717 36001 18751
rect 36035 18717 36047 18751
rect 37844 18748 37872 18788
rect 37918 18776 37924 18828
rect 37976 18776 37982 18828
rect 38286 18776 38292 18828
rect 38344 18816 38350 18828
rect 38344 18788 39252 18816
rect 38344 18776 38350 18788
rect 39224 18760 39252 18788
rect 40402 18776 40408 18828
rect 40460 18816 40466 18828
rect 41141 18819 41199 18825
rect 41141 18816 41153 18819
rect 40460 18788 41153 18816
rect 40460 18776 40466 18788
rect 41141 18785 41153 18788
rect 41187 18785 41199 18819
rect 42153 18819 42211 18825
rect 42153 18816 42165 18819
rect 41141 18779 41199 18785
rect 41340 18788 42165 18816
rect 38105 18751 38163 18757
rect 38105 18748 38117 18751
rect 37844 18720 38117 18748
rect 35989 18711 36047 18717
rect 38105 18717 38117 18720
rect 38151 18717 38163 18751
rect 39117 18751 39175 18757
rect 39117 18748 39129 18751
rect 38105 18711 38163 18717
rect 38856 18720 39129 18748
rect 15664 18652 16436 18680
rect 15565 18615 15623 18621
rect 15565 18581 15577 18615
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 16022 18572 16028 18624
rect 16080 18572 16086 18624
rect 16408 18612 16436 18652
rect 16669 18683 16727 18689
rect 16669 18649 16681 18683
rect 16715 18680 16727 18683
rect 17218 18680 17224 18692
rect 16715 18652 17224 18680
rect 16715 18649 16727 18652
rect 16669 18643 16727 18649
rect 17218 18640 17224 18652
rect 17276 18640 17282 18692
rect 17586 18640 17592 18692
rect 17644 18640 17650 18692
rect 18874 18680 18880 18692
rect 18814 18652 18880 18680
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 19426 18640 19432 18692
rect 19484 18680 19490 18692
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 19484 18652 19625 18680
rect 19484 18640 19490 18652
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 19613 18643 19671 18649
rect 22094 18640 22100 18692
rect 22152 18680 22158 18692
rect 22465 18683 22523 18689
rect 22465 18680 22477 18683
rect 22152 18652 22477 18680
rect 22152 18640 22158 18652
rect 22465 18649 22477 18652
rect 22511 18649 22523 18683
rect 25884 18680 25912 18708
rect 26329 18683 26387 18689
rect 26329 18680 26341 18683
rect 25884 18652 26341 18680
rect 22465 18643 22523 18649
rect 26329 18649 26341 18652
rect 26375 18649 26387 18683
rect 26329 18643 26387 18649
rect 28994 18640 29000 18692
rect 29052 18680 29058 18692
rect 29362 18680 29368 18692
rect 29052 18652 29368 18680
rect 29052 18640 29058 18652
rect 29362 18640 29368 18652
rect 29420 18680 29426 18692
rect 35345 18683 35403 18689
rect 29420 18652 31602 18680
rect 29420 18640 29426 18652
rect 35345 18649 35357 18683
rect 35391 18680 35403 18683
rect 35713 18683 35771 18689
rect 35713 18680 35725 18683
rect 35391 18652 35725 18680
rect 35391 18649 35403 18652
rect 35345 18643 35403 18649
rect 35713 18649 35725 18652
rect 35759 18649 35771 18683
rect 35713 18643 35771 18649
rect 37645 18683 37703 18689
rect 37645 18649 37657 18683
rect 37691 18649 37703 18683
rect 37645 18643 37703 18649
rect 17954 18612 17960 18624
rect 16408 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 19705 18615 19763 18621
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 19978 18612 19984 18624
rect 19751 18584 19984 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 19978 18572 19984 18584
rect 20036 18612 20042 18624
rect 20073 18615 20131 18621
rect 20073 18612 20085 18615
rect 20036 18584 20085 18612
rect 20036 18572 20042 18584
rect 20073 18581 20085 18584
rect 20119 18581 20131 18615
rect 20073 18575 20131 18581
rect 21910 18572 21916 18624
rect 21968 18572 21974 18624
rect 24581 18615 24639 18621
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 24670 18612 24676 18624
rect 24627 18584 24676 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 26602 18572 26608 18624
rect 26660 18612 26666 18624
rect 37550 18612 37556 18624
rect 26660 18584 37556 18612
rect 26660 18572 26666 18584
rect 37550 18572 37556 18584
rect 37608 18572 37614 18624
rect 37660 18612 37688 18643
rect 37826 18640 37832 18692
rect 37884 18640 37890 18692
rect 38746 18680 38752 18692
rect 37936 18652 38752 18680
rect 37936 18612 37964 18652
rect 38746 18640 38752 18652
rect 38804 18680 38810 18692
rect 38856 18689 38884 18720
rect 39117 18717 39129 18720
rect 39163 18717 39175 18751
rect 39117 18711 39175 18717
rect 39206 18708 39212 18760
rect 39264 18708 39270 18760
rect 39298 18708 39304 18760
rect 39356 18708 39362 18760
rect 39485 18751 39543 18757
rect 39485 18717 39497 18751
rect 39531 18748 39543 18751
rect 40420 18748 40448 18776
rect 39531 18720 40448 18748
rect 40957 18751 41015 18757
rect 39531 18717 39543 18720
rect 39485 18711 39543 18717
rect 40957 18717 40969 18751
rect 41003 18717 41015 18751
rect 40957 18711 41015 18717
rect 38841 18683 38899 18689
rect 38841 18680 38853 18683
rect 38804 18652 38853 18680
rect 38804 18640 38810 18652
rect 38841 18649 38853 18652
rect 38887 18649 38899 18683
rect 38841 18643 38899 18649
rect 39025 18683 39083 18689
rect 39025 18649 39037 18683
rect 39071 18680 39083 18683
rect 39316 18680 39344 18708
rect 39071 18652 39344 18680
rect 39393 18683 39451 18689
rect 39071 18649 39083 18652
rect 39025 18643 39083 18649
rect 39393 18649 39405 18683
rect 39439 18680 39451 18683
rect 40218 18680 40224 18692
rect 39439 18652 40224 18680
rect 39439 18649 39451 18652
rect 39393 18643 39451 18649
rect 40218 18640 40224 18652
rect 40276 18680 40282 18692
rect 40972 18680 41000 18711
rect 41230 18708 41236 18760
rect 41288 18708 41294 18760
rect 41340 18757 41368 18788
rect 42153 18785 42165 18788
rect 42199 18785 42211 18819
rect 42352 18816 42380 18912
rect 42702 18884 42708 18896
rect 42628 18856 42708 18884
rect 42628 18825 42656 18856
rect 42702 18844 42708 18856
rect 42760 18844 42766 18896
rect 42521 18819 42579 18825
rect 42521 18816 42533 18819
rect 42352 18788 42533 18816
rect 42153 18779 42211 18785
rect 42521 18785 42533 18788
rect 42567 18785 42579 18819
rect 42521 18779 42579 18785
rect 42613 18819 42671 18825
rect 42613 18785 42625 18819
rect 42659 18785 42671 18819
rect 42904 18816 42932 18912
rect 42613 18779 42671 18785
rect 42720 18788 42932 18816
rect 41325 18751 41383 18757
rect 41325 18717 41337 18751
rect 41371 18717 41383 18751
rect 41325 18711 41383 18717
rect 41509 18751 41567 18757
rect 41509 18717 41521 18751
rect 41555 18748 41567 18751
rect 41601 18751 41659 18757
rect 41601 18748 41613 18751
rect 41555 18720 41613 18748
rect 41555 18717 41567 18720
rect 41509 18711 41567 18717
rect 41601 18717 41613 18720
rect 41647 18717 41659 18751
rect 41601 18711 41659 18717
rect 41874 18708 41880 18760
rect 41932 18708 41938 18760
rect 41966 18708 41972 18760
rect 42024 18708 42030 18760
rect 42720 18757 42748 18788
rect 42337 18751 42395 18757
rect 42337 18717 42349 18751
rect 42383 18717 42395 18751
rect 42337 18711 42395 18717
rect 42705 18751 42763 18757
rect 42705 18717 42717 18751
rect 42751 18717 42763 18751
rect 42705 18711 42763 18717
rect 42889 18751 42947 18757
rect 42889 18717 42901 18751
rect 42935 18748 42947 18751
rect 42978 18748 42984 18760
rect 42935 18720 42984 18748
rect 42935 18717 42947 18720
rect 42889 18711 42947 18717
rect 41785 18683 41843 18689
rect 41785 18680 41797 18683
rect 40276 18652 41000 18680
rect 41616 18652 41797 18680
rect 40276 18640 40282 18652
rect 41616 18624 41644 18652
rect 41785 18649 41797 18652
rect 41831 18649 41843 18683
rect 41892 18680 41920 18708
rect 42352 18680 42380 18711
rect 42978 18708 42984 18720
rect 43036 18708 43042 18760
rect 43070 18708 43076 18760
rect 43128 18708 43134 18760
rect 41892 18652 42380 18680
rect 43349 18683 43407 18689
rect 41785 18643 41843 18649
rect 43349 18649 43361 18683
rect 43395 18680 43407 18683
rect 43622 18680 43628 18692
rect 43395 18652 43628 18680
rect 43395 18649 43407 18652
rect 43349 18643 43407 18649
rect 43622 18640 43628 18652
rect 43680 18640 43686 18692
rect 37660 18584 37964 18612
rect 38654 18572 38660 18624
rect 38712 18572 38718 18624
rect 39666 18572 39672 18624
rect 39724 18572 39730 18624
rect 40770 18572 40776 18624
rect 40828 18572 40834 18624
rect 41598 18572 41604 18624
rect 41656 18572 41662 18624
rect 43165 18615 43223 18621
rect 43165 18581 43177 18615
rect 43211 18612 43223 18615
rect 43438 18612 43444 18624
rect 43211 18584 43444 18612
rect 43211 18581 43223 18584
rect 43165 18575 43223 18581
rect 43438 18572 43444 18584
rect 43496 18572 43502 18624
rect 1104 18522 44620 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 44620 18522
rect 1104 18448 44620 18470
rect 2222 18368 2228 18420
rect 2280 18368 2286 18420
rect 2777 18411 2835 18417
rect 2777 18377 2789 18411
rect 2823 18408 2835 18411
rect 3142 18408 3148 18420
rect 2823 18380 3148 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 7374 18408 7380 18420
rect 6656 18380 7380 18408
rect 2240 18272 2268 18368
rect 4706 18300 4712 18352
rect 4764 18300 4770 18352
rect 6656 18349 6684 18380
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 8113 18411 8171 18417
rect 8113 18377 8125 18411
rect 8159 18408 8171 18411
rect 9214 18408 9220 18420
rect 8159 18380 9220 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 10192 18380 10517 18408
rect 10192 18368 10198 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 10778 18368 10784 18420
rect 10836 18368 10842 18420
rect 10870 18368 10876 18420
rect 10928 18368 10934 18420
rect 12342 18368 12348 18420
rect 12400 18368 12406 18420
rect 12802 18368 12808 18420
rect 12860 18368 12866 18420
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 18325 18411 18383 18417
rect 18325 18408 18337 18411
rect 17644 18380 18337 18408
rect 17644 18368 17650 18380
rect 18325 18377 18337 18380
rect 18371 18377 18383 18411
rect 18325 18371 18383 18377
rect 18877 18411 18935 18417
rect 18877 18377 18889 18411
rect 18923 18377 18935 18411
rect 18877 18371 18935 18377
rect 19245 18411 19303 18417
rect 19245 18377 19257 18411
rect 19291 18408 19303 18411
rect 19978 18408 19984 18420
rect 19291 18380 19984 18408
rect 19291 18377 19303 18380
rect 19245 18371 19303 18377
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18309 6699 18343
rect 6641 18303 6699 18309
rect 8478 18300 8484 18352
rect 8536 18340 8542 18352
rect 8573 18343 8631 18349
rect 8573 18340 8585 18343
rect 8536 18312 8585 18340
rect 8536 18300 8542 18312
rect 8573 18309 8585 18312
rect 8619 18309 8631 18343
rect 8573 18303 8631 18309
rect 9030 18300 9036 18352
rect 9088 18300 9094 18352
rect 10321 18343 10379 18349
rect 10321 18309 10333 18343
rect 10367 18340 10379 18343
rect 10796 18340 10824 18368
rect 10367 18312 10824 18340
rect 10367 18309 10379 18312
rect 10321 18303 10379 18309
rect 2593 18275 2651 18281
rect 2593 18272 2605 18275
rect 2240 18244 2605 18272
rect 2593 18241 2605 18244
rect 2639 18241 2651 18275
rect 7774 18244 7880 18272
rect 2593 18235 2651 18241
rect 7852 18216 7880 18244
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18272 10747 18275
rect 10888 18272 10916 18368
rect 12713 18343 12771 18349
rect 12713 18309 12725 18343
rect 12759 18340 12771 18343
rect 12820 18340 12848 18368
rect 12759 18312 12848 18340
rect 12759 18309 12771 18312
rect 12713 18303 12771 18309
rect 14366 18300 14372 18352
rect 14424 18340 14430 18352
rect 14461 18343 14519 18349
rect 14461 18340 14473 18343
rect 14424 18312 14473 18340
rect 14424 18300 14430 18312
rect 14461 18309 14473 18312
rect 14507 18309 14519 18343
rect 14461 18303 14519 18309
rect 10735 18244 10916 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 16485 18275 16543 18281
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18173 3387 18207
rect 3329 18167 3387 18173
rect 3344 18080 3372 18167
rect 3694 18164 3700 18216
rect 3752 18164 3758 18216
rect 5123 18207 5181 18213
rect 5123 18173 5135 18207
rect 5169 18204 5181 18207
rect 5537 18207 5595 18213
rect 5537 18204 5549 18207
rect 5169 18176 5549 18204
rect 5169 18173 5181 18176
rect 5123 18167 5181 18173
rect 5537 18173 5549 18176
rect 5583 18173 5595 18207
rect 5537 18167 5595 18173
rect 6365 18207 6423 18213
rect 6365 18173 6377 18207
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 6086 18136 6092 18148
rect 4632 18108 6092 18136
rect 4632 18080 4660 18108
rect 6086 18096 6092 18108
rect 6144 18136 6150 18148
rect 6380 18136 6408 18167
rect 7834 18164 7840 18216
rect 7892 18164 7898 18216
rect 11790 18164 11796 18216
rect 11848 18164 11854 18216
rect 6144 18108 6408 18136
rect 6144 18096 6150 18108
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 4614 18068 4620 18080
rect 3384 18040 4620 18068
rect 3384 18028 3390 18040
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 6178 18028 6184 18080
rect 6236 18028 6242 18080
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 13832 18068 13860 18258
rect 16485 18241 16497 18275
rect 16531 18272 16543 18275
rect 16574 18272 16580 18284
rect 16531 18244 16580 18272
rect 16531 18241 16543 18244
rect 16485 18235 16543 18241
rect 16574 18232 16580 18244
rect 16632 18232 16638 18284
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18272 18567 18275
rect 18892 18272 18920 18371
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20456 18380 22094 18408
rect 20456 18352 20484 18380
rect 20438 18300 20444 18352
rect 20496 18300 20502 18352
rect 20806 18300 20812 18352
rect 20864 18300 20870 18352
rect 18555 18244 18920 18272
rect 18555 18241 18567 18244
rect 18509 18235 18567 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 22066 18272 22094 18380
rect 23106 18368 23112 18420
rect 23164 18368 23170 18420
rect 23293 18411 23351 18417
rect 23293 18377 23305 18411
rect 23339 18408 23351 18411
rect 23382 18408 23388 18420
rect 23339 18380 23388 18408
rect 23339 18377 23351 18380
rect 23293 18371 23351 18377
rect 22741 18343 22799 18349
rect 22741 18309 22753 18343
rect 22787 18340 22799 18343
rect 23308 18340 23336 18371
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 26234 18408 26240 18420
rect 23808 18380 26240 18408
rect 23808 18368 23814 18380
rect 22787 18312 23336 18340
rect 22787 18309 22799 18312
rect 22741 18303 22799 18309
rect 24026 18300 24032 18352
rect 24084 18300 24090 18352
rect 24670 18300 24676 18352
rect 24728 18340 24734 18352
rect 24765 18343 24823 18349
rect 24765 18340 24777 18343
rect 24728 18312 24777 18340
rect 24728 18300 24734 18312
rect 24765 18309 24777 18312
rect 24811 18309 24823 18343
rect 24765 18303 24823 18309
rect 25056 18281 25084 18380
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 37918 18368 37924 18420
rect 37976 18368 37982 18420
rect 38286 18368 38292 18420
rect 38344 18368 38350 18420
rect 38654 18368 38660 18420
rect 38712 18368 38718 18420
rect 38838 18368 38844 18420
rect 38896 18408 38902 18420
rect 39574 18408 39580 18420
rect 38896 18380 39580 18408
rect 38896 18368 38902 18380
rect 39574 18368 39580 18380
rect 39632 18368 39638 18420
rect 39666 18368 39672 18420
rect 39724 18368 39730 18420
rect 40770 18368 40776 18420
rect 40828 18368 40834 18420
rect 41230 18368 41236 18420
rect 41288 18408 41294 18420
rect 41325 18411 41383 18417
rect 41325 18408 41337 18411
rect 41288 18380 41337 18408
rect 41288 18368 41294 18380
rect 41325 18377 41337 18380
rect 41371 18377 41383 18411
rect 41325 18371 41383 18377
rect 43622 18368 43628 18420
rect 43680 18368 43686 18420
rect 25130 18300 25136 18352
rect 25188 18340 25194 18352
rect 25682 18340 25688 18352
rect 25188 18312 25688 18340
rect 25188 18300 25194 18312
rect 25682 18300 25688 18312
rect 25740 18300 25746 18352
rect 37936 18340 37964 18368
rect 29196 18312 29868 18340
rect 35374 18312 36216 18340
rect 29196 18284 29224 18312
rect 25041 18275 25099 18281
rect 19300 18244 19472 18272
rect 22066 18244 23612 18272
rect 19300 18232 19306 18244
rect 19058 18164 19064 18216
rect 19116 18204 19122 18216
rect 19444 18213 19472 18244
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 19116 18176 19349 18204
rect 19116 18164 19122 18176
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18204 20223 18207
rect 20714 18204 20720 18216
rect 20211 18176 20720 18204
rect 20211 18173 20223 18176
rect 20165 18167 20223 18173
rect 10836 18040 13860 18068
rect 10836 18028 10842 18040
rect 16298 18028 16304 18080
rect 16356 18028 16362 18080
rect 19904 18068 19932 18167
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 22557 18207 22615 18213
rect 22557 18173 22569 18207
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18204 22707 18207
rect 22830 18204 22836 18216
rect 22695 18176 22836 18204
rect 22695 18173 22707 18176
rect 22649 18167 22707 18173
rect 22572 18136 22600 18167
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 23474 18164 23480 18216
rect 23532 18164 23538 18216
rect 23584 18204 23612 18244
rect 25041 18241 25053 18275
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 25516 18204 25544 18235
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 25648 18244 26157 18272
rect 25648 18232 25654 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 26145 18235 26203 18241
rect 29178 18232 29184 18284
rect 29236 18232 29242 18284
rect 29638 18232 29644 18284
rect 29696 18232 29702 18284
rect 29840 18281 29868 18312
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18241 29883 18275
rect 29825 18235 29883 18241
rect 30098 18232 30104 18284
rect 30156 18232 30162 18284
rect 26421 18207 26479 18213
rect 26421 18204 26433 18207
rect 23584 18176 26433 18204
rect 26421 18173 26433 18176
rect 26467 18204 26479 18207
rect 27062 18204 27068 18216
rect 26467 18176 27068 18204
rect 26467 18173 26479 18176
rect 26421 18167 26479 18173
rect 27062 18164 27068 18176
rect 27120 18164 27126 18216
rect 30190 18164 30196 18216
rect 30248 18164 30254 18216
rect 30469 18207 30527 18213
rect 30469 18173 30481 18207
rect 30515 18204 30527 18207
rect 31662 18204 31668 18216
rect 30515 18176 31668 18204
rect 30515 18173 30527 18176
rect 30469 18167 30527 18173
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 35710 18164 35716 18216
rect 35768 18204 35774 18216
rect 35805 18207 35863 18213
rect 35805 18204 35817 18207
rect 35768 18176 35817 18204
rect 35768 18164 35774 18176
rect 35805 18173 35817 18176
rect 35851 18173 35863 18207
rect 36081 18207 36139 18213
rect 36081 18204 36093 18207
rect 35805 18167 35863 18173
rect 36004 18176 36093 18204
rect 23492 18136 23520 18164
rect 22572 18108 23520 18136
rect 36004 18080 36032 18176
rect 36081 18173 36093 18176
rect 36127 18173 36139 18207
rect 36081 18167 36139 18173
rect 36188 18136 36216 18312
rect 36832 18312 37964 18340
rect 36832 18281 36860 18312
rect 36265 18275 36323 18281
rect 36265 18241 36277 18275
rect 36311 18241 36323 18275
rect 36265 18235 36323 18241
rect 36817 18275 36875 18281
rect 36817 18241 36829 18275
rect 36863 18241 36875 18275
rect 36817 18235 36875 18241
rect 37645 18275 37703 18281
rect 37645 18241 37657 18275
rect 37691 18272 37703 18275
rect 38013 18275 38071 18281
rect 38013 18272 38025 18275
rect 37691 18244 38025 18272
rect 37691 18241 37703 18244
rect 37645 18235 37703 18241
rect 38013 18241 38025 18244
rect 38059 18241 38071 18275
rect 38013 18235 38071 18241
rect 36280 18204 36308 18235
rect 37458 18204 37464 18216
rect 36280 18176 37464 18204
rect 37458 18164 37464 18176
rect 37516 18164 37522 18216
rect 37737 18207 37795 18213
rect 37737 18173 37749 18207
rect 37783 18204 37795 18207
rect 38304 18204 38332 18368
rect 38672 18272 38700 18368
rect 38749 18275 38807 18281
rect 38749 18272 38761 18275
rect 38672 18244 38761 18272
rect 38749 18241 38761 18244
rect 38795 18241 38807 18275
rect 38856 18272 38884 18368
rect 39684 18340 39712 18368
rect 39132 18312 39712 18340
rect 39132 18281 39160 18312
rect 38933 18275 38991 18281
rect 38933 18272 38945 18275
rect 38856 18244 38945 18272
rect 38749 18235 38807 18241
rect 38933 18241 38945 18244
rect 38979 18241 38991 18275
rect 38933 18235 38991 18241
rect 39117 18275 39175 18281
rect 39117 18241 39129 18275
rect 39163 18241 39175 18275
rect 39117 18235 39175 18241
rect 39301 18275 39359 18281
rect 39301 18241 39313 18275
rect 39347 18241 39359 18275
rect 39301 18235 39359 18241
rect 37783 18176 38332 18204
rect 38657 18207 38715 18213
rect 37783 18173 37795 18176
rect 37737 18167 37795 18173
rect 38657 18173 38669 18207
rect 38703 18204 38715 18207
rect 39025 18207 39083 18213
rect 39025 18204 39037 18207
rect 38703 18176 39037 18204
rect 38703 18173 38715 18176
rect 38657 18167 38715 18173
rect 39025 18173 39037 18176
rect 39071 18173 39083 18207
rect 39316 18204 39344 18235
rect 39390 18232 39396 18284
rect 39448 18272 39454 18284
rect 39577 18275 39635 18281
rect 39577 18272 39589 18275
rect 39448 18244 39589 18272
rect 39448 18232 39454 18244
rect 39577 18241 39589 18244
rect 39623 18241 39635 18275
rect 39577 18235 39635 18241
rect 39666 18232 39672 18284
rect 39724 18272 39730 18284
rect 39761 18275 39819 18281
rect 39761 18272 39773 18275
rect 39724 18244 39773 18272
rect 39724 18232 39730 18244
rect 39761 18241 39773 18244
rect 39807 18241 39819 18275
rect 39761 18235 39819 18241
rect 40788 18204 40816 18368
rect 41693 18343 41751 18349
rect 41693 18309 41705 18343
rect 41739 18340 41751 18343
rect 42334 18340 42340 18352
rect 41739 18312 42340 18340
rect 41739 18309 41751 18312
rect 41693 18303 41751 18309
rect 42334 18300 42340 18312
rect 42392 18300 42398 18352
rect 41509 18275 41567 18281
rect 41509 18241 41521 18275
rect 41555 18241 41567 18275
rect 41509 18235 41567 18241
rect 39316 18176 40816 18204
rect 41524 18204 41552 18235
rect 41598 18232 41604 18284
rect 41656 18232 41662 18284
rect 41874 18232 41880 18284
rect 41932 18232 41938 18284
rect 41966 18232 41972 18284
rect 42024 18232 42030 18284
rect 43346 18232 43352 18284
rect 43404 18232 43410 18284
rect 41984 18204 42012 18232
rect 41524 18176 42012 18204
rect 39025 18167 39083 18173
rect 36541 18139 36599 18145
rect 36541 18136 36553 18139
rect 36188 18108 36553 18136
rect 36541 18105 36553 18108
rect 36587 18136 36599 18139
rect 37182 18136 37188 18148
rect 36587 18108 37188 18136
rect 36587 18105 36599 18108
rect 36541 18099 36599 18105
rect 37182 18096 37188 18108
rect 37240 18096 37246 18148
rect 39040 18136 39068 18167
rect 44174 18164 44180 18216
rect 44232 18164 44238 18216
rect 39114 18136 39120 18148
rect 39040 18108 39120 18136
rect 39114 18096 39120 18108
rect 39172 18136 39178 18148
rect 39390 18136 39396 18148
rect 39172 18108 39396 18136
rect 39172 18096 39178 18108
rect 39390 18096 39396 18108
rect 39448 18096 39454 18148
rect 20622 18068 20628 18080
rect 19904 18040 20628 18068
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 21634 18028 21640 18080
rect 21692 18028 21698 18080
rect 25866 18028 25872 18080
rect 25924 18028 25930 18080
rect 25961 18071 26019 18077
rect 25961 18037 25973 18071
rect 26007 18068 26019 18071
rect 26050 18068 26056 18080
rect 26007 18040 26056 18068
rect 26007 18037 26019 18040
rect 25961 18031 26019 18037
rect 26050 18028 26056 18040
rect 26108 18028 26114 18080
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 26329 18071 26387 18077
rect 26329 18068 26341 18071
rect 26292 18040 26341 18068
rect 26292 18028 26298 18040
rect 26329 18037 26341 18040
rect 26375 18037 26387 18071
rect 26329 18031 26387 18037
rect 29825 18071 29883 18077
rect 29825 18037 29837 18071
rect 29871 18068 29883 18071
rect 30374 18068 30380 18080
rect 29871 18040 30380 18068
rect 29871 18037 29883 18040
rect 29825 18031 29883 18037
rect 30374 18028 30380 18040
rect 30432 18028 30438 18080
rect 34333 18071 34391 18077
rect 34333 18037 34345 18071
rect 34379 18068 34391 18071
rect 34698 18068 34704 18080
rect 34379 18040 34704 18068
rect 34379 18037 34391 18040
rect 34333 18031 34391 18037
rect 34698 18028 34704 18040
rect 34756 18028 34762 18080
rect 35986 18028 35992 18080
rect 36044 18028 36050 18080
rect 37001 18071 37059 18077
rect 37001 18037 37013 18071
rect 37047 18068 37059 18071
rect 37274 18068 37280 18080
rect 37047 18040 37280 18068
rect 37047 18037 37059 18040
rect 37001 18031 37059 18037
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 37366 18028 37372 18080
rect 37424 18028 37430 18080
rect 38930 18028 38936 18080
rect 38988 18068 38994 18080
rect 39485 18071 39543 18077
rect 39485 18068 39497 18071
rect 38988 18040 39497 18068
rect 38988 18028 38994 18040
rect 39485 18037 39497 18040
rect 39531 18037 39543 18071
rect 39485 18031 39543 18037
rect 39574 18028 39580 18080
rect 39632 18068 39638 18080
rect 39669 18071 39727 18077
rect 39669 18068 39681 18071
rect 39632 18040 39681 18068
rect 39632 18028 39638 18040
rect 39669 18037 39681 18040
rect 39715 18037 39727 18071
rect 39669 18031 39727 18037
rect 42794 18028 42800 18080
rect 42852 18028 42858 18080
rect 1104 17978 44620 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 44620 17978
rect 1104 17904 44620 17926
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 3694 17864 3700 17876
rect 3651 17836 3700 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 9548 17836 10088 17864
rect 9548 17824 9554 17836
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 6144 17700 6193 17728
rect 6144 17688 6150 17700
rect 6181 17697 6193 17700
rect 6227 17728 6239 17731
rect 7006 17728 7012 17740
rect 6227 17700 7012 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 7650 17688 7656 17740
rect 7708 17688 7714 17740
rect 10060 17737 10088 17836
rect 11882 17824 11888 17876
rect 11940 17824 11946 17876
rect 12621 17867 12679 17873
rect 12621 17833 12633 17867
rect 12667 17864 12679 17867
rect 12986 17864 12992 17876
rect 12667 17836 12992 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 14936 17836 20668 17864
rect 14936 17808 14964 17836
rect 12434 17796 12440 17808
rect 12406 17756 12440 17796
rect 12492 17756 12498 17808
rect 14918 17756 14924 17808
rect 14976 17756 14982 17808
rect 17310 17756 17316 17808
rect 17368 17756 17374 17808
rect 20640 17796 20668 17836
rect 20714 17824 20720 17876
rect 20772 17824 20778 17876
rect 21910 17864 21916 17876
rect 21376 17836 21916 17864
rect 20640 17768 21312 17796
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 7975 17700 9505 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 12406 17728 12434 17756
rect 10091 17700 12434 17728
rect 13265 17731 13323 17737
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 13265 17697 13277 17731
rect 13311 17728 13323 17731
rect 13446 17728 13452 17740
rect 13311 17700 13452 17728
rect 13311 17697 13323 17700
rect 13265 17691 13323 17697
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 17328 17728 17356 17756
rect 15979 17700 17356 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17920 17700 17969 17728
rect 17920 17688 17926 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2832 17632 2973 17660
rect 2832 17620 2838 17632
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 7668 17660 7696 17688
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 7668 17632 8585 17660
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 12437 17663 12495 17669
rect 12437 17660 12449 17663
rect 8573 17623 8631 17629
rect 11808 17632 12449 17660
rect 5813 17595 5871 17601
rect 5813 17561 5825 17595
rect 5859 17592 5871 17595
rect 6178 17592 6184 17604
rect 5859 17564 6184 17592
rect 5859 17561 5871 17564
rect 5813 17555 5871 17561
rect 6178 17552 6184 17564
rect 6236 17552 6242 17604
rect 6454 17552 6460 17604
rect 6512 17552 6518 17604
rect 6546 17552 6552 17604
rect 6604 17592 6610 17604
rect 6604 17564 6946 17592
rect 6604 17552 6610 17564
rect 9030 17552 9036 17604
rect 9088 17552 9094 17604
rect 10318 17552 10324 17604
rect 10376 17552 10382 17604
rect 10778 17592 10784 17604
rect 10612 17564 10784 17592
rect 4338 17484 4344 17536
rect 4396 17484 4402 17536
rect 8018 17484 8024 17536
rect 8076 17484 8082 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 8720 17496 8953 17524
rect 8720 17484 8726 17496
rect 8941 17493 8953 17496
rect 8987 17493 8999 17527
rect 9048 17524 9076 17552
rect 10612 17524 10640 17564
rect 10778 17552 10784 17564
rect 10836 17552 10842 17604
rect 11808 17533 11836 17632
rect 12437 17629 12449 17632
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 14366 17660 14372 17672
rect 13035 17632 14372 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 14366 17620 14372 17632
rect 14424 17620 14430 17672
rect 14550 17620 14556 17672
rect 14608 17620 14614 17672
rect 14642 17620 14648 17672
rect 14700 17620 14706 17672
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17660 20959 17663
rect 20947 17632 21036 17660
rect 20947 17629 20959 17632
rect 20901 17623 20959 17629
rect 13817 17595 13875 17601
rect 13817 17561 13829 17595
rect 13863 17592 13875 17595
rect 14660 17592 14688 17620
rect 13863 17564 14688 17592
rect 16209 17595 16267 17601
rect 13863 17561 13875 17564
rect 13817 17555 13875 17561
rect 16209 17561 16221 17595
rect 16255 17592 16267 17595
rect 16298 17592 16304 17604
rect 16255 17564 16304 17592
rect 16255 17561 16267 17564
rect 16209 17555 16267 17561
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 17586 17592 17592 17604
rect 17434 17564 17592 17592
rect 17586 17552 17592 17564
rect 17644 17592 17650 17604
rect 17644 17564 18920 17592
rect 17644 17552 17650 17564
rect 18892 17536 18920 17564
rect 9048 17496 10640 17524
rect 11793 17527 11851 17533
rect 8941 17487 8999 17493
rect 11793 17493 11805 17527
rect 11839 17493 11851 17527
rect 11793 17487 11851 17493
rect 13078 17484 13084 17536
rect 13136 17484 13142 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 13504 17496 13553 17524
rect 13504 17484 13510 17496
rect 13541 17493 13553 17496
rect 13587 17493 13599 17527
rect 13541 17487 13599 17493
rect 14366 17484 14372 17536
rect 14424 17484 14430 17536
rect 18874 17484 18880 17536
rect 18932 17484 18938 17536
rect 21008 17533 21036 17632
rect 21284 17592 21312 17768
rect 21376 17669 21404 17836
rect 21910 17824 21916 17836
rect 21968 17864 21974 17876
rect 22465 17867 22523 17873
rect 22465 17864 22477 17867
rect 21968 17836 22477 17864
rect 21968 17824 21974 17836
rect 22465 17833 22477 17836
rect 22511 17833 22523 17867
rect 22465 17827 22523 17833
rect 25866 17824 25872 17876
rect 25924 17864 25930 17876
rect 27249 17867 27307 17873
rect 27249 17864 27261 17867
rect 25924 17836 27261 17864
rect 25924 17824 25930 17836
rect 26068 17805 26096 17836
rect 27249 17833 27261 17836
rect 27295 17833 27307 17867
rect 27249 17827 27307 17833
rect 27338 17824 27344 17876
rect 27396 17864 27402 17876
rect 30098 17864 30104 17876
rect 27396 17836 28028 17864
rect 27396 17824 27402 17836
rect 22557 17799 22615 17805
rect 22557 17796 22569 17799
rect 21468 17768 22569 17796
rect 21468 17672 21496 17768
rect 22557 17765 22569 17768
rect 22603 17765 22615 17799
rect 22557 17759 22615 17765
rect 26053 17799 26111 17805
rect 26053 17765 26065 17799
rect 26099 17765 26111 17799
rect 26053 17759 26111 17765
rect 26145 17799 26203 17805
rect 26145 17765 26157 17799
rect 26191 17796 26203 17799
rect 26234 17796 26240 17808
rect 26191 17768 26240 17796
rect 26191 17765 26203 17768
rect 26145 17759 26203 17765
rect 26234 17756 26240 17768
rect 26292 17796 26298 17808
rect 27430 17796 27436 17808
rect 26292 17768 27436 17796
rect 26292 17756 26298 17768
rect 21545 17731 21603 17737
rect 21545 17697 21557 17731
rect 21591 17697 21603 17731
rect 21545 17691 21603 17697
rect 21361 17663 21419 17669
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 21560 17660 21588 17691
rect 21634 17688 21640 17740
rect 21692 17728 21698 17740
rect 21821 17731 21879 17737
rect 21821 17728 21833 17731
rect 21692 17700 21833 17728
rect 21692 17688 21698 17700
rect 21821 17697 21833 17700
rect 21867 17697 21879 17731
rect 25774 17728 25780 17740
rect 21821 17691 21879 17697
rect 22066 17700 25780 17728
rect 21726 17660 21732 17672
rect 21560 17632 21732 17660
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 22066 17592 22094 17700
rect 25774 17688 25780 17700
rect 25832 17728 25838 17740
rect 27172 17737 27200 17768
rect 27430 17756 27436 17768
rect 27488 17756 27494 17808
rect 27614 17756 27620 17808
rect 27672 17756 27678 17808
rect 26421 17731 26479 17737
rect 25832 17700 26188 17728
rect 25832 17688 25838 17700
rect 23106 17620 23112 17672
rect 23164 17620 23170 17672
rect 25590 17620 25596 17672
rect 25648 17660 25654 17672
rect 25961 17663 26019 17669
rect 25961 17660 25973 17663
rect 25648 17632 25973 17660
rect 25648 17620 25654 17632
rect 25961 17629 25973 17632
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 21284 17564 22094 17592
rect 20993 17527 21051 17533
rect 20993 17493 21005 17527
rect 21039 17493 21051 17527
rect 20993 17487 21051 17493
rect 21450 17484 21456 17536
rect 21508 17484 21514 17536
rect 25976 17524 26004 17623
rect 26160 17592 26188 17700
rect 26421 17697 26433 17731
rect 26467 17728 26479 17731
rect 26605 17731 26663 17737
rect 26605 17728 26617 17731
rect 26467 17700 26617 17728
rect 26467 17697 26479 17700
rect 26421 17691 26479 17697
rect 26605 17697 26617 17700
rect 26651 17697 26663 17731
rect 26605 17691 26663 17697
rect 27157 17731 27215 17737
rect 27157 17697 27169 17731
rect 27203 17697 27215 17731
rect 27157 17691 27215 17697
rect 26237 17663 26295 17669
rect 26237 17629 26249 17663
rect 26283 17660 26295 17663
rect 26326 17660 26332 17672
rect 26283 17632 26332 17660
rect 26283 17629 26295 17632
rect 26237 17623 26295 17629
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 26697 17663 26755 17669
rect 26697 17629 26709 17663
rect 26743 17629 26755 17663
rect 27433 17663 27491 17669
rect 27433 17660 27445 17663
rect 26697 17623 26755 17629
rect 26804 17632 27445 17660
rect 26712 17592 26740 17623
rect 26160 17564 26740 17592
rect 26804 17524 26832 17632
rect 27433 17629 27445 17632
rect 27479 17660 27491 17663
rect 27522 17660 27528 17672
rect 27479 17632 27528 17660
rect 27479 17629 27491 17632
rect 27433 17623 27491 17629
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 27632 17660 27660 17756
rect 27699 17663 27757 17669
rect 27699 17660 27711 17663
rect 27632 17632 27711 17660
rect 27699 17629 27711 17632
rect 27745 17629 27757 17663
rect 27699 17623 27757 17629
rect 27890 17620 27896 17672
rect 27948 17620 27954 17672
rect 28000 17592 28028 17836
rect 29840 17836 30104 17864
rect 29840 17737 29868 17836
rect 30098 17824 30104 17836
rect 30156 17864 30162 17876
rect 30745 17867 30803 17873
rect 30745 17864 30757 17867
rect 30156 17836 30757 17864
rect 30156 17824 30162 17836
rect 30745 17833 30757 17836
rect 30791 17833 30803 17867
rect 30745 17827 30803 17833
rect 38746 17824 38752 17876
rect 38804 17824 38810 17876
rect 40218 17824 40224 17876
rect 40276 17864 40282 17876
rect 41601 17867 41659 17873
rect 41601 17864 41613 17867
rect 40276 17836 41613 17864
rect 40276 17824 40282 17836
rect 41601 17833 41613 17836
rect 41647 17833 41659 17867
rect 42794 17864 42800 17876
rect 41601 17827 41659 17833
rect 42444 17836 42800 17864
rect 30006 17756 30012 17808
rect 30064 17796 30070 17808
rect 30193 17799 30251 17805
rect 30193 17796 30205 17799
rect 30064 17768 30205 17796
rect 30064 17756 30070 17768
rect 30193 17765 30205 17768
rect 30239 17765 30251 17799
rect 30193 17759 30251 17765
rect 30374 17756 30380 17808
rect 30432 17756 30438 17808
rect 33045 17799 33103 17805
rect 33045 17796 33057 17799
rect 31588 17768 33057 17796
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17728 29055 17731
rect 29365 17731 29423 17737
rect 29043 17700 29316 17728
rect 29043 17697 29055 17700
rect 28997 17691 29055 17697
rect 29178 17620 29184 17672
rect 29236 17620 29242 17672
rect 29288 17660 29316 17700
rect 29365 17697 29377 17731
rect 29411 17728 29423 17731
rect 29733 17731 29791 17737
rect 29733 17728 29745 17731
rect 29411 17700 29745 17728
rect 29411 17697 29423 17700
rect 29365 17691 29423 17697
rect 29733 17697 29745 17700
rect 29779 17697 29791 17731
rect 29733 17691 29791 17697
rect 29825 17731 29883 17737
rect 29825 17697 29837 17731
rect 29871 17697 29883 17731
rect 29825 17691 29883 17697
rect 29917 17731 29975 17737
rect 29917 17697 29929 17731
rect 29963 17728 29975 17731
rect 30282 17728 30288 17740
rect 29963 17700 30288 17728
rect 29963 17697 29975 17700
rect 29917 17691 29975 17697
rect 29288 17632 29500 17660
rect 29196 17592 29224 17620
rect 28000 17564 29224 17592
rect 25976 17496 26832 17524
rect 27065 17527 27123 17533
rect 27065 17493 27077 17527
rect 27111 17524 27123 17527
rect 27338 17524 27344 17536
rect 27111 17496 27344 17524
rect 27111 17493 27123 17496
rect 27065 17487 27123 17493
rect 27338 17484 27344 17496
rect 27396 17484 27402 17536
rect 27614 17484 27620 17536
rect 27672 17484 27678 17536
rect 27798 17484 27804 17536
rect 27856 17484 27862 17536
rect 29472 17524 29500 17632
rect 29546 17620 29552 17672
rect 29604 17620 29610 17672
rect 29748 17592 29776 17691
rect 30282 17688 30288 17700
rect 30340 17688 30346 17740
rect 30009 17663 30067 17669
rect 30009 17629 30021 17663
rect 30055 17660 30067 17663
rect 30098 17660 30104 17672
rect 30055 17632 30104 17660
rect 30055 17629 30067 17632
rect 30009 17623 30067 17629
rect 30098 17620 30104 17632
rect 30156 17620 30162 17672
rect 30392 17660 30420 17756
rect 31588 17740 31616 17768
rect 33045 17765 33057 17768
rect 33091 17796 33103 17799
rect 33502 17796 33508 17808
rect 33091 17768 33508 17796
rect 33091 17765 33103 17768
rect 33045 17759 33103 17765
rect 33502 17756 33508 17768
rect 33560 17756 33566 17808
rect 31570 17688 31576 17740
rect 31628 17688 31634 17740
rect 32232 17700 32904 17728
rect 32232 17672 32260 17700
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 30392 17632 30573 17660
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 31938 17620 31944 17672
rect 31996 17620 32002 17672
rect 32214 17620 32220 17672
rect 32272 17620 32278 17672
rect 32306 17620 32312 17672
rect 32364 17660 32370 17672
rect 32876 17669 32904 17700
rect 37274 17688 37280 17740
rect 37332 17688 37338 17740
rect 42334 17728 42340 17740
rect 41432 17700 42340 17728
rect 32769 17663 32827 17669
rect 32769 17660 32781 17663
rect 32364 17632 32781 17660
rect 32364 17620 32370 17632
rect 32769 17629 32781 17632
rect 32815 17629 32827 17663
rect 32769 17623 32827 17629
rect 32861 17663 32919 17669
rect 32861 17629 32873 17663
rect 32907 17629 32919 17663
rect 32861 17623 32919 17629
rect 33137 17663 33195 17669
rect 33137 17629 33149 17663
rect 33183 17660 33195 17663
rect 33594 17660 33600 17672
rect 33183 17632 33600 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 33594 17620 33600 17632
rect 33652 17620 33658 17672
rect 36998 17660 37004 17672
rect 36464 17632 37004 17660
rect 30377 17595 30435 17601
rect 30377 17592 30389 17595
rect 29748 17564 30389 17592
rect 30377 17561 30389 17564
rect 30423 17561 30435 17595
rect 30377 17555 30435 17561
rect 31110 17552 31116 17604
rect 31168 17592 31174 17604
rect 31956 17592 31984 17620
rect 35161 17595 35219 17601
rect 35161 17592 35173 17595
rect 31168 17564 35173 17592
rect 31168 17552 31174 17564
rect 35161 17561 35173 17564
rect 35207 17561 35219 17595
rect 35161 17555 35219 17561
rect 29638 17524 29644 17536
rect 29472 17496 29644 17524
rect 29638 17484 29644 17496
rect 29696 17524 29702 17536
rect 30006 17524 30012 17536
rect 29696 17496 30012 17524
rect 29696 17484 29702 17496
rect 30006 17484 30012 17496
rect 30064 17484 30070 17536
rect 32398 17484 32404 17536
rect 32456 17524 32462 17536
rect 32585 17527 32643 17533
rect 32585 17524 32597 17527
rect 32456 17496 32597 17524
rect 32456 17484 32462 17496
rect 32585 17493 32597 17496
rect 32631 17493 32643 17527
rect 32585 17487 32643 17493
rect 35986 17484 35992 17536
rect 36044 17524 36050 17536
rect 36464 17533 36492 17632
rect 36998 17620 37004 17632
rect 37056 17620 37062 17672
rect 39390 17620 39396 17672
rect 39448 17660 39454 17672
rect 39577 17663 39635 17669
rect 39577 17660 39589 17663
rect 39448 17632 39589 17660
rect 39448 17620 39454 17632
rect 39577 17629 39589 17632
rect 39623 17629 39635 17663
rect 39577 17623 39635 17629
rect 39853 17663 39911 17669
rect 39853 17629 39865 17663
rect 39899 17629 39911 17663
rect 39853 17623 39911 17629
rect 39868 17592 39896 17623
rect 37200 17564 37766 17592
rect 39868 17564 39988 17592
rect 37200 17536 37228 17564
rect 39960 17536 39988 17564
rect 40126 17552 40132 17604
rect 40184 17552 40190 17604
rect 41432 17592 41460 17700
rect 42334 17688 42340 17700
rect 42392 17688 42398 17740
rect 42444 17669 42472 17836
rect 42794 17824 42800 17836
rect 42852 17824 42858 17876
rect 42794 17688 42800 17740
rect 42852 17728 42858 17740
rect 44174 17728 44180 17740
rect 42852 17700 44180 17728
rect 42852 17688 42858 17700
rect 44174 17688 44180 17700
rect 44232 17728 44238 17740
rect 44269 17731 44327 17737
rect 44269 17728 44281 17731
rect 44232 17700 44281 17728
rect 44232 17688 44238 17700
rect 44269 17697 44281 17700
rect 44315 17697 44327 17731
rect 44269 17691 44327 17697
rect 42245 17663 42303 17669
rect 42245 17660 42257 17663
rect 41354 17564 41460 17592
rect 36449 17527 36507 17533
rect 36449 17524 36461 17527
rect 36044 17496 36461 17524
rect 36044 17484 36050 17496
rect 36449 17493 36461 17496
rect 36495 17493 36507 17527
rect 36449 17487 36507 17493
rect 37182 17484 37188 17536
rect 37240 17484 37246 17536
rect 39022 17484 39028 17536
rect 39080 17484 39086 17536
rect 39942 17484 39948 17536
rect 40000 17484 40006 17536
rect 40862 17484 40868 17536
rect 40920 17524 40926 17536
rect 41432 17524 41460 17564
rect 42168 17632 42257 17660
rect 42168 17536 42196 17632
rect 42245 17629 42257 17632
rect 42291 17629 42303 17663
rect 42245 17623 42303 17629
rect 42429 17663 42487 17669
rect 42429 17629 42441 17663
rect 42475 17629 42487 17663
rect 42429 17623 42487 17629
rect 42518 17620 42524 17672
rect 42576 17620 42582 17672
rect 42337 17595 42395 17601
rect 42337 17561 42349 17595
rect 42383 17592 42395 17595
rect 42797 17595 42855 17601
rect 42797 17592 42809 17595
rect 42383 17564 42809 17592
rect 42383 17561 42395 17564
rect 42337 17555 42395 17561
rect 42797 17561 42809 17564
rect 42843 17561 42855 17595
rect 42797 17555 42855 17561
rect 42904 17564 43286 17592
rect 40920 17496 41460 17524
rect 40920 17484 40926 17496
rect 42150 17484 42156 17536
rect 42208 17484 42214 17536
rect 42426 17484 42432 17536
rect 42484 17524 42490 17536
rect 42904 17524 42932 17564
rect 42484 17496 42932 17524
rect 42484 17484 42490 17496
rect 1104 17434 44620 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 44620 17434
rect 1104 17360 44620 17382
rect 4338 17280 4344 17332
rect 4396 17280 4402 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5353 17323 5411 17329
rect 5353 17320 5365 17323
rect 5132 17292 5365 17320
rect 5132 17280 5138 17292
rect 5353 17289 5365 17292
rect 5399 17289 5411 17323
rect 5353 17283 5411 17289
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 6512 17292 6929 17320
rect 6512 17280 6518 17292
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 8938 17320 8944 17332
rect 6917 17283 6975 17289
rect 7852 17292 8944 17320
rect 4356 17184 4384 17280
rect 7852 17252 7880 17292
rect 6932 17224 7880 17252
rect 7929 17255 7987 17261
rect 6932 17196 6960 17224
rect 7929 17221 7941 17255
rect 7975 17252 7987 17255
rect 8018 17252 8024 17264
rect 7975 17224 8024 17252
rect 7975 17221 7987 17224
rect 7929 17215 7987 17221
rect 8018 17212 8024 17224
rect 8076 17212 8082 17264
rect 8312 17252 8340 17292
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10376 17292 10701 17320
rect 10376 17280 10382 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 8312 17224 8418 17252
rect 4709 17187 4767 17193
rect 4709 17184 4721 17187
rect 4356 17156 4721 17184
rect 4709 17153 4721 17156
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6914 17184 6920 17196
rect 5859 17156 6920 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7653 17187 7711 17193
rect 7653 17184 7665 17187
rect 7024 17156 7665 17184
rect 7024 17128 7052 17156
rect 7653 17153 7665 17156
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11532 17184 11560 17283
rect 11882 17280 11888 17332
rect 11940 17280 11946 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16632 17292 16681 17320
rect 16632 17280 16638 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 16669 17283 16727 17289
rect 17037 17323 17095 17329
rect 17037 17289 17049 17323
rect 17083 17320 17095 17323
rect 17862 17320 17868 17332
rect 17083 17292 17868 17320
rect 17083 17289 17095 17292
rect 17037 17283 17095 17289
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 18932 17292 19840 17320
rect 18932 17280 18938 17292
rect 16390 17212 16396 17264
rect 16448 17212 16454 17264
rect 12894 17184 12900 17196
rect 10919 17156 11560 17184
rect 12176 17156 12900 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17116 7619 17119
rect 8938 17116 8944 17128
rect 7607 17088 8944 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9447 17088 9965 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 11974 17076 11980 17128
rect 12032 17076 12038 17128
rect 12176 17125 12204 17156
rect 12894 17144 12900 17156
rect 12952 17184 12958 17196
rect 13446 17184 13452 17196
rect 12952 17156 13452 17184
rect 12952 17144 12958 17156
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 17129 17187 17187 17193
rect 15528 17156 16344 17184
rect 15528 17144 15534 17156
rect 12161 17119 12219 17125
rect 12161 17085 12173 17119
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 12492 17088 14105 17116
rect 12492 17076 12498 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 14918 17076 14924 17128
rect 14976 17116 14982 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 14976 17088 15853 17116
rect 14976 17076 14982 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 4764 16952 5917 16980
rect 4764 16940 4770 16952
rect 5905 16949 5917 16952
rect 5951 16980 5963 16983
rect 6546 16980 6552 16992
rect 5951 16952 6552 16980
rect 5951 16949 5963 16952
rect 5905 16943 5963 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 10594 16940 10600 16992
rect 10652 16940 10658 16992
rect 16316 16989 16344 17156
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17494 17184 17500 17196
rect 17175 17156 17500 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 19812 17184 19840 17292
rect 27798 17280 27804 17332
rect 27856 17280 27862 17332
rect 29546 17280 29552 17332
rect 29604 17280 29610 17332
rect 30101 17323 30159 17329
rect 30101 17289 30113 17323
rect 30147 17320 30159 17323
rect 30190 17320 30196 17332
rect 30147 17292 30196 17320
rect 30147 17289 30159 17292
rect 30101 17283 30159 17289
rect 30190 17280 30196 17292
rect 30248 17280 30254 17332
rect 34146 17320 34152 17332
rect 33244 17292 34152 17320
rect 20438 17212 20444 17264
rect 20496 17212 20502 17264
rect 20806 17252 20812 17264
rect 20548 17224 20812 17252
rect 20548 17196 20576 17224
rect 20806 17212 20812 17224
rect 20864 17212 20870 17264
rect 22554 17212 22560 17264
rect 22612 17212 22618 17264
rect 20530 17184 20536 17196
rect 19812 17170 20536 17184
rect 19826 17156 20536 17170
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 20680 17156 21833 17184
rect 20680 17144 20686 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 25682 17144 25688 17196
rect 25740 17184 25746 17196
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25740 17156 25973 17184
rect 25740 17144 25746 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 27062 17144 27068 17196
rect 27120 17144 27126 17196
rect 27816 17184 27844 17280
rect 28077 17255 28135 17261
rect 28077 17221 28089 17255
rect 28123 17252 28135 17255
rect 31570 17252 31576 17264
rect 28123 17224 31576 17252
rect 28123 17221 28135 17224
rect 28077 17215 28135 17221
rect 31570 17212 31576 17224
rect 31628 17212 31634 17264
rect 27738 17156 27844 17184
rect 29178 17144 29184 17196
rect 29236 17144 29242 17196
rect 29733 17187 29791 17193
rect 29733 17153 29745 17187
rect 29779 17184 29791 17187
rect 30285 17187 30343 17193
rect 30285 17184 30297 17187
rect 29779 17156 30297 17184
rect 29779 17153 29791 17156
rect 29733 17147 29791 17153
rect 30285 17153 30297 17156
rect 30331 17184 30343 17187
rect 30466 17184 30472 17196
rect 30331 17156 30472 17184
rect 30331 17153 30343 17156
rect 30285 17147 30343 17153
rect 30466 17144 30472 17156
rect 30524 17144 30530 17196
rect 32125 17187 32183 17193
rect 32125 17153 32137 17187
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 17218 17076 17224 17128
rect 17276 17076 17282 17128
rect 18046 17076 18052 17128
rect 18104 17076 18110 17128
rect 18322 17076 18328 17128
rect 18380 17116 18386 17128
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 18380 17088 18429 17116
rect 18380 17076 18386 17088
rect 18417 17085 18429 17088
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 22186 17116 22192 17128
rect 22143 17088 22192 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 23569 17119 23627 17125
rect 23569 17085 23581 17119
rect 23615 17116 23627 17119
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 23615 17088 24225 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 26050 17076 26056 17128
rect 26108 17076 26114 17128
rect 26789 17119 26847 17125
rect 26789 17085 26801 17119
rect 26835 17085 26847 17119
rect 29196 17116 29224 17144
rect 29917 17119 29975 17125
rect 29917 17116 29929 17119
rect 29196 17088 29929 17116
rect 26789 17079 26847 17085
rect 29917 17085 29929 17088
rect 29963 17085 29975 17119
rect 29917 17079 29975 17085
rect 30009 17119 30067 17125
rect 30009 17085 30021 17119
rect 30055 17116 30067 17119
rect 30098 17116 30104 17128
rect 30055 17088 30104 17116
rect 30055 17085 30067 17088
rect 30009 17079 30067 17085
rect 26804 17048 26832 17079
rect 30098 17076 30104 17088
rect 30156 17076 30162 17128
rect 30190 17076 30196 17128
rect 30248 17116 30254 17128
rect 30558 17116 30564 17128
rect 30248 17088 30564 17116
rect 30248 17076 30254 17088
rect 30558 17076 30564 17088
rect 30616 17076 30622 17128
rect 32140 17116 32168 17147
rect 32214 17144 32220 17196
rect 32272 17144 32278 17196
rect 32398 17144 32404 17196
rect 32456 17144 32462 17196
rect 33244 17193 33272 17292
rect 34146 17280 34152 17292
rect 34204 17280 34210 17332
rect 34422 17320 34428 17332
rect 34256 17292 34428 17320
rect 34256 17252 34284 17292
rect 34422 17280 34428 17292
rect 34480 17280 34486 17332
rect 37366 17280 37372 17332
rect 37424 17280 37430 17332
rect 38838 17280 38844 17332
rect 38896 17280 38902 17332
rect 39025 17323 39083 17329
rect 39025 17289 39037 17323
rect 39071 17320 39083 17323
rect 39114 17320 39120 17332
rect 39071 17292 39120 17320
rect 39071 17289 39083 17292
rect 39025 17283 39083 17289
rect 39114 17280 39120 17292
rect 39172 17280 39178 17332
rect 39206 17280 39212 17332
rect 39264 17280 39270 17332
rect 39390 17280 39396 17332
rect 39448 17320 39454 17332
rect 39491 17323 39549 17329
rect 39491 17320 39503 17323
rect 39448 17292 39503 17320
rect 39448 17280 39454 17292
rect 39491 17289 39503 17292
rect 39537 17289 39549 17323
rect 39491 17283 39549 17289
rect 39577 17323 39635 17329
rect 39577 17289 39589 17323
rect 39623 17320 39635 17323
rect 41598 17320 41604 17332
rect 39623 17292 41604 17320
rect 39623 17289 39635 17292
rect 39577 17283 39635 17289
rect 33428 17224 34284 17252
rect 37384 17252 37412 17280
rect 37553 17255 37611 17261
rect 37553 17252 37565 17255
rect 37384 17224 37565 17252
rect 33428 17193 33456 17224
rect 32953 17187 33011 17193
rect 32953 17153 32965 17187
rect 32999 17153 33011 17187
rect 32953 17147 33011 17153
rect 33229 17187 33287 17193
rect 33229 17153 33241 17187
rect 33275 17153 33287 17187
rect 33229 17147 33287 17153
rect 33413 17187 33471 17193
rect 33413 17153 33425 17187
rect 33459 17153 33471 17187
rect 33413 17147 33471 17153
rect 32306 17116 32312 17128
rect 32140 17088 32312 17116
rect 32140 17060 32168 17088
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 32585 17119 32643 17125
rect 32585 17085 32597 17119
rect 32631 17116 32643 17119
rect 32968 17116 32996 17147
rect 33502 17144 33508 17196
rect 33560 17144 33566 17196
rect 33594 17144 33600 17196
rect 33652 17184 33658 17196
rect 33689 17187 33747 17193
rect 33689 17184 33701 17187
rect 33652 17156 33701 17184
rect 33652 17144 33658 17156
rect 33689 17153 33701 17156
rect 33735 17153 33747 17187
rect 33689 17147 33747 17153
rect 32631 17088 32996 17116
rect 33704 17116 33732 17147
rect 33778 17144 33784 17196
rect 33836 17184 33842 17196
rect 33965 17187 34023 17193
rect 33965 17184 33977 17187
rect 33836 17156 33977 17184
rect 33836 17144 33842 17156
rect 33965 17153 33977 17156
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34146 17144 34152 17196
rect 34204 17144 34210 17196
rect 34256 17193 34284 17224
rect 37553 17221 37565 17224
rect 37599 17221 37611 17255
rect 38856 17252 38884 17280
rect 40005 17255 40063 17261
rect 40005 17252 40017 17255
rect 38856 17224 39344 17252
rect 37553 17215 37611 17221
rect 34241 17187 34299 17193
rect 34241 17153 34253 17187
rect 34287 17153 34299 17187
rect 34241 17147 34299 17153
rect 34330 17144 34336 17196
rect 34388 17184 34394 17196
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34388 17156 34437 17184
rect 34388 17144 34394 17156
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34425 17147 34483 17153
rect 34698 17144 34704 17196
rect 34756 17144 34762 17196
rect 36998 17144 37004 17196
rect 37056 17184 37062 17196
rect 39316 17193 39344 17224
rect 39776 17224 40017 17252
rect 39776 17196 39804 17224
rect 40005 17221 40017 17224
rect 40051 17221 40063 17255
rect 40005 17215 40063 17221
rect 40218 17212 40224 17264
rect 40276 17212 40282 17264
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 37056 17156 37289 17184
rect 37056 17144 37062 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 39117 17187 39175 17193
rect 37277 17147 37335 17153
rect 34609 17119 34667 17125
rect 34609 17116 34621 17119
rect 33704 17088 34621 17116
rect 32631 17085 32643 17088
rect 32585 17079 32643 17085
rect 34609 17085 34621 17088
rect 34655 17085 34667 17119
rect 34609 17079 34667 17085
rect 37182 17076 37188 17128
rect 37240 17116 37246 17128
rect 38672 17116 38700 17170
rect 39117 17153 39129 17187
rect 39163 17153 39175 17187
rect 39117 17147 39175 17153
rect 39301 17187 39359 17193
rect 39301 17153 39313 17187
rect 39347 17153 39359 17187
rect 39301 17147 39359 17153
rect 39393 17187 39451 17193
rect 39393 17153 39405 17187
rect 39439 17153 39451 17187
rect 39393 17147 39451 17153
rect 39669 17187 39727 17193
rect 39669 17153 39681 17187
rect 39715 17184 39727 17187
rect 39758 17184 39764 17196
rect 39715 17156 39764 17184
rect 39715 17153 39727 17156
rect 39669 17147 39727 17153
rect 37240 17088 38700 17116
rect 37240 17076 37246 17088
rect 38746 17076 38752 17128
rect 38804 17116 38810 17128
rect 39132 17116 39160 17147
rect 38804 17088 39160 17116
rect 38804 17076 38810 17088
rect 32122 17048 32128 17060
rect 26804 17020 32128 17048
rect 32122 17008 32128 17020
rect 32180 17008 32186 17060
rect 33137 17051 33195 17057
rect 32232 17020 32720 17048
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 17586 16980 17592 16992
rect 16347 16952 17592 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 22646 16980 22652 16992
rect 18564 16952 22652 16980
rect 18564 16940 18570 16952
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 22830 16940 22836 16992
rect 22888 16980 22894 16992
rect 23661 16983 23719 16989
rect 23661 16980 23673 16983
rect 22888 16952 23673 16980
rect 22888 16940 22894 16952
rect 23661 16949 23673 16952
rect 23707 16949 23719 16983
rect 23661 16943 23719 16949
rect 30374 16940 30380 16992
rect 30432 16980 30438 16992
rect 30469 16983 30527 16989
rect 30469 16980 30481 16983
rect 30432 16952 30481 16980
rect 30432 16940 30438 16952
rect 30469 16949 30481 16952
rect 30515 16980 30527 16983
rect 31386 16980 31392 16992
rect 30515 16952 31392 16980
rect 30515 16949 30527 16952
rect 30469 16943 30527 16949
rect 31386 16940 31392 16952
rect 31444 16980 31450 16992
rect 32232 16980 32260 17020
rect 32692 16989 32720 17020
rect 33137 17017 33149 17051
rect 33183 17048 33195 17051
rect 34057 17051 34115 17057
rect 34057 17048 34069 17051
rect 33183 17020 34069 17048
rect 33183 17017 33195 17020
rect 33137 17011 33195 17017
rect 34057 17017 34069 17020
rect 34103 17017 34115 17051
rect 39316 17048 39344 17147
rect 39408 17116 39436 17147
rect 39758 17144 39764 17156
rect 39816 17144 39822 17196
rect 40236 17184 40264 17212
rect 40236 17156 40724 17184
rect 40589 17119 40647 17125
rect 40589 17116 40601 17119
rect 39408 17088 40601 17116
rect 40589 17085 40601 17088
rect 40635 17085 40647 17119
rect 40696 17116 40724 17156
rect 41141 17119 41199 17125
rect 41141 17116 41153 17119
rect 40696 17088 41153 17116
rect 40589 17079 40647 17085
rect 41141 17085 41153 17088
rect 41187 17085 41199 17119
rect 41141 17079 41199 17085
rect 39853 17051 39911 17057
rect 39853 17048 39865 17051
rect 39316 17020 39865 17048
rect 34057 17011 34115 17017
rect 39853 17017 39865 17020
rect 39899 17017 39911 17051
rect 39853 17011 39911 17017
rect 41386 17048 41414 17292
rect 41598 17280 41604 17292
rect 41656 17280 41662 17332
rect 43257 17323 43315 17329
rect 43257 17289 43269 17323
rect 43303 17289 43315 17323
rect 43257 17283 43315 17289
rect 43425 17323 43483 17329
rect 43425 17289 43437 17323
rect 43471 17320 43483 17323
rect 43530 17320 43536 17332
rect 43471 17292 43536 17320
rect 43471 17289 43483 17292
rect 43425 17283 43483 17289
rect 42150 17252 42156 17264
rect 42076 17224 42156 17252
rect 42076 17193 42104 17224
rect 42150 17212 42156 17224
rect 42208 17252 42214 17264
rect 43272 17252 43300 17283
rect 43530 17280 43536 17292
rect 43588 17280 43594 17332
rect 42208 17224 43300 17252
rect 43625 17255 43683 17261
rect 42208 17212 42214 17224
rect 43625 17221 43637 17255
rect 43671 17252 43683 17255
rect 44174 17252 44180 17264
rect 43671 17224 44180 17252
rect 43671 17221 43683 17224
rect 43625 17215 43683 17221
rect 44174 17212 44180 17224
rect 44232 17212 44238 17264
rect 41785 17187 41843 17193
rect 41785 17153 41797 17187
rect 41831 17184 41843 17187
rect 42061 17187 42119 17193
rect 42061 17184 42073 17187
rect 41831 17156 42073 17184
rect 41831 17153 41843 17156
rect 41785 17147 41843 17153
rect 42061 17153 42073 17156
rect 42107 17153 42119 17187
rect 42061 17147 42119 17153
rect 42245 17187 42303 17193
rect 42245 17153 42257 17187
rect 42291 17184 42303 17187
rect 42521 17187 42579 17193
rect 42521 17184 42533 17187
rect 42291 17156 42533 17184
rect 42291 17153 42303 17156
rect 42245 17147 42303 17153
rect 42521 17153 42533 17156
rect 42567 17153 42579 17187
rect 42521 17147 42579 17153
rect 41874 17076 41880 17128
rect 41932 17116 41938 17128
rect 41969 17119 42027 17125
rect 41969 17116 41981 17119
rect 41932 17088 41981 17116
rect 41932 17076 41938 17088
rect 41969 17085 41981 17088
rect 42015 17116 42027 17119
rect 42702 17116 42708 17128
rect 42015 17088 42708 17116
rect 42015 17085 42027 17088
rect 41969 17079 42027 17085
rect 42702 17076 42708 17088
rect 42760 17116 42766 17128
rect 43073 17119 43131 17125
rect 43073 17116 43085 17119
rect 42760 17088 43085 17116
rect 42760 17076 42766 17088
rect 43073 17085 43085 17088
rect 43119 17085 43131 17119
rect 43073 17079 43131 17085
rect 41386 17020 42196 17048
rect 31444 16952 32260 16980
rect 32677 16983 32735 16989
rect 31444 16940 31450 16952
rect 32677 16949 32689 16983
rect 32723 16949 32735 16983
rect 32677 16943 32735 16949
rect 33042 16940 33048 16992
rect 33100 16940 33106 16992
rect 33686 16940 33692 16992
rect 33744 16980 33750 16992
rect 33873 16983 33931 16989
rect 33873 16980 33885 16983
rect 33744 16952 33885 16980
rect 33744 16940 33750 16952
rect 33873 16949 33885 16952
rect 33919 16949 33931 16983
rect 33873 16943 33931 16949
rect 34425 16983 34483 16989
rect 34425 16949 34437 16983
rect 34471 16980 34483 16983
rect 34514 16980 34520 16992
rect 34471 16952 34520 16980
rect 34471 16949 34483 16952
rect 34425 16943 34483 16949
rect 34514 16940 34520 16952
rect 34572 16940 34578 16992
rect 40037 16983 40095 16989
rect 40037 16949 40049 16983
rect 40083 16980 40095 16983
rect 41386 16980 41414 17020
rect 42168 16992 42196 17020
rect 40083 16952 41414 16980
rect 40083 16949 40095 16952
rect 40037 16943 40095 16949
rect 41598 16940 41604 16992
rect 41656 16940 41662 16992
rect 42058 16940 42064 16992
rect 42116 16940 42122 16992
rect 42150 16940 42156 16992
rect 42208 16940 42214 16992
rect 43438 16940 43444 16992
rect 43496 16980 43502 16992
rect 44266 16980 44272 16992
rect 43496 16952 44272 16980
rect 43496 16940 43502 16952
rect 44266 16940 44272 16952
rect 44324 16940 44330 16992
rect 1104 16890 44620 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 44620 16890
rect 1104 16816 44620 16838
rect 8938 16736 8944 16788
rect 8996 16736 9002 16788
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 10594 16736 10600 16788
rect 10652 16736 10658 16788
rect 12434 16776 12440 16788
rect 11440 16748 12440 16776
rect 9048 16572 9076 16736
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 10612 16640 10640 16736
rect 11440 16649 11468 16748
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 13136 16748 13277 16776
rect 13136 16736 13142 16748
rect 13265 16745 13277 16748
rect 13311 16745 13323 16779
rect 13265 16739 13323 16745
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 17218 16776 17224 16788
rect 15212 16748 17224 16776
rect 15212 16649 15240 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17681 16779 17739 16785
rect 17681 16745 17693 16779
rect 17727 16776 17739 16779
rect 18046 16776 18052 16788
rect 17727 16748 18052 16776
rect 17727 16745 17739 16748
rect 17681 16739 17739 16745
rect 18046 16736 18052 16748
rect 18104 16736 18110 16788
rect 18690 16736 18696 16788
rect 18748 16736 18754 16788
rect 21729 16779 21787 16785
rect 21729 16745 21741 16779
rect 21775 16776 21787 16779
rect 22186 16776 22192 16788
rect 21775 16748 22192 16776
rect 21775 16745 21787 16748
rect 21729 16739 21787 16745
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 27614 16736 27620 16788
rect 27672 16736 27678 16788
rect 30098 16736 30104 16788
rect 30156 16776 30162 16788
rect 30377 16779 30435 16785
rect 30377 16776 30389 16779
rect 30156 16748 30389 16776
rect 30156 16736 30162 16748
rect 30377 16745 30389 16748
rect 30423 16745 30435 16779
rect 30377 16739 30435 16745
rect 32677 16779 32735 16785
rect 32677 16745 32689 16779
rect 32723 16776 32735 16779
rect 33042 16776 33048 16788
rect 32723 16748 33048 16776
rect 32723 16745 32735 16748
rect 32677 16739 32735 16745
rect 33042 16736 33048 16748
rect 33100 16736 33106 16788
rect 33229 16779 33287 16785
rect 33229 16745 33241 16779
rect 33275 16776 33287 16779
rect 34146 16776 34152 16788
rect 33275 16748 34152 16776
rect 33275 16745 33287 16748
rect 33229 16739 33287 16745
rect 34146 16736 34152 16748
rect 34204 16736 34210 16788
rect 38838 16736 38844 16788
rect 38896 16736 38902 16788
rect 39022 16736 39028 16788
rect 39080 16736 39086 16788
rect 39301 16779 39359 16785
rect 39301 16745 39313 16779
rect 39347 16776 39359 16779
rect 40126 16776 40132 16788
rect 39347 16748 40132 16776
rect 39347 16745 39359 16748
rect 39301 16739 39359 16745
rect 40126 16736 40132 16748
rect 40184 16736 40190 16788
rect 40497 16779 40555 16785
rect 40497 16745 40509 16779
rect 40543 16776 40555 16779
rect 40862 16776 40868 16788
rect 40543 16748 40868 16776
rect 40543 16745 40555 16748
rect 40497 16739 40555 16745
rect 40862 16736 40868 16748
rect 40920 16736 40926 16788
rect 42702 16736 42708 16788
rect 42760 16736 42766 16788
rect 17236 16708 17264 16736
rect 19334 16708 19340 16720
rect 17236 16680 19340 16708
rect 19334 16668 19340 16680
rect 19392 16708 19398 16720
rect 19392 16680 19840 16708
rect 19392 16668 19398 16680
rect 10459 16612 10640 16640
rect 10689 16643 10747 16649
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 10735 16612 11437 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16609 13875 16643
rect 13817 16603 13875 16609
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 18322 16640 18328 16652
rect 15979 16612 18328 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 9306 16572 9312 16584
rect 9048 16544 9312 16572
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 13832 16572 13860 16603
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 19812 16649 19840 16680
rect 22646 16668 22652 16720
rect 22704 16708 22710 16720
rect 22704 16680 27200 16708
rect 22704 16668 22710 16680
rect 27172 16652 27200 16680
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20346 16600 20352 16652
rect 20404 16640 20410 16652
rect 21726 16640 21732 16652
rect 20404 16612 21732 16640
rect 20404 16600 20410 16612
rect 21726 16600 21732 16612
rect 21784 16640 21790 16652
rect 22370 16640 22376 16652
rect 21784 16612 22376 16640
rect 21784 16600 21790 16612
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23474 16600 23480 16652
rect 23532 16640 23538 16652
rect 25041 16643 25099 16649
rect 25041 16640 25053 16643
rect 23532 16612 25053 16640
rect 23532 16600 23538 16612
rect 25041 16609 25053 16612
rect 25087 16640 25099 16643
rect 26602 16640 26608 16652
rect 25087 16612 26608 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 26602 16600 26608 16612
rect 26660 16600 26666 16652
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16640 27399 16643
rect 27632 16640 27660 16736
rect 33502 16708 33508 16720
rect 33152 16680 33508 16708
rect 27387 16612 27660 16640
rect 30024 16612 30420 16640
rect 27387 16609 27399 16612
rect 27341 16603 27399 16609
rect 13188 16544 13860 16572
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 6822 16504 6828 16516
rect 6411 16476 6828 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 6822 16464 6828 16476
rect 6880 16464 6886 16516
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7064 16408 7665 16436
rect 7064 16396 7070 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 9324 16436 9352 16532
rect 11698 16464 11704 16516
rect 11756 16464 11762 16516
rect 11808 16476 12190 16504
rect 11808 16436 11836 16476
rect 13188 16445 13216 16544
rect 14918 16532 14924 16584
rect 14976 16532 14982 16584
rect 17586 16572 17592 16584
rect 17342 16544 17592 16572
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19613 16575 19671 16581
rect 18923 16544 19288 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 16255 16476 16620 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 16592 16448 16620 16476
rect 9324 16408 11836 16436
rect 13173 16439 13231 16445
rect 7653 16399 7711 16405
rect 13173 16405 13185 16439
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 15013 16439 15071 16445
rect 15013 16405 15025 16439
rect 15059 16436 15071 16439
rect 15102 16436 15108 16448
rect 15059 16408 15108 16436
rect 15059 16405 15071 16408
rect 15013 16399 15071 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 16574 16396 16580 16448
rect 16632 16396 16638 16448
rect 19260 16445 19288 16544
rect 19613 16541 19625 16575
rect 19659 16572 19671 16575
rect 20438 16572 20444 16584
rect 19659 16544 20444 16572
rect 19659 16541 19671 16544
rect 19613 16535 19671 16541
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16572 21603 16575
rect 22189 16575 22247 16581
rect 21591 16544 21864 16572
rect 21591 16541 21603 16544
rect 21545 16535 21603 16541
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 19705 16439 19763 16445
rect 19705 16405 19717 16439
rect 19751 16436 19763 16439
rect 19978 16436 19984 16448
rect 19751 16408 19984 16436
rect 19751 16405 19763 16408
rect 19705 16399 19763 16405
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 21836 16445 21864 16544
rect 22189 16541 22201 16575
rect 22235 16572 22247 16575
rect 22830 16572 22836 16584
rect 22235 16544 22836 16572
rect 22235 16541 22247 16544
rect 22189 16535 22247 16541
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16572 23903 16575
rect 24765 16575 24823 16581
rect 23891 16544 24440 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 21821 16439 21879 16445
rect 21821 16405 21833 16439
rect 21867 16405 21879 16439
rect 21821 16399 21879 16405
rect 22278 16396 22284 16448
rect 22336 16396 22342 16448
rect 23661 16439 23719 16445
rect 23661 16405 23673 16439
rect 23707 16436 23719 16439
rect 23842 16436 23848 16448
rect 23707 16408 23848 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 24412 16445 24440 16544
rect 24765 16541 24777 16575
rect 24811 16572 24823 16575
rect 25682 16572 25688 16584
rect 24811 16544 25688 16572
rect 24811 16541 24823 16544
rect 24765 16535 24823 16541
rect 25682 16532 25688 16544
rect 25740 16532 25746 16584
rect 26326 16532 26332 16584
rect 26384 16572 26390 16584
rect 27249 16575 27307 16581
rect 27249 16572 27261 16575
rect 26384 16544 27261 16572
rect 26384 16532 26390 16544
rect 27249 16541 27261 16544
rect 27295 16541 27307 16575
rect 27249 16535 27307 16541
rect 29546 16532 29552 16584
rect 29604 16572 29610 16584
rect 30024 16581 30052 16612
rect 29825 16575 29883 16581
rect 29825 16572 29837 16575
rect 29604 16544 29837 16572
rect 29604 16532 29610 16544
rect 29825 16541 29837 16544
rect 29871 16541 29883 16575
rect 29825 16535 29883 16541
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 30285 16575 30343 16581
rect 30285 16541 30297 16575
rect 30331 16541 30343 16575
rect 30285 16535 30343 16541
rect 24857 16507 24915 16513
rect 24857 16504 24869 16507
rect 24688 16476 24869 16504
rect 24688 16448 24716 16476
rect 24857 16473 24869 16476
rect 24903 16473 24915 16507
rect 24857 16467 24915 16473
rect 30190 16464 30196 16516
rect 30248 16464 30254 16516
rect 24397 16439 24455 16445
rect 24397 16405 24409 16439
rect 24443 16405 24455 16439
rect 24397 16399 24455 16405
rect 24670 16396 24676 16448
rect 24728 16396 24734 16448
rect 27617 16439 27675 16445
rect 27617 16405 27629 16439
rect 27663 16436 27675 16439
rect 29638 16436 29644 16448
rect 27663 16408 29644 16436
rect 27663 16405 27675 16408
rect 27617 16399 27675 16405
rect 29638 16396 29644 16408
rect 29696 16396 29702 16448
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 30300 16436 30328 16535
rect 30392 16504 30420 16612
rect 32122 16600 32128 16652
rect 32180 16640 32186 16652
rect 32309 16643 32367 16649
rect 32309 16640 32321 16643
rect 32180 16612 32321 16640
rect 32180 16600 32186 16612
rect 32309 16609 32321 16612
rect 32355 16609 32367 16643
rect 32309 16603 32367 16609
rect 30466 16532 30472 16584
rect 30524 16572 30530 16584
rect 30561 16575 30619 16581
rect 30561 16572 30573 16575
rect 30524 16544 30573 16572
rect 30524 16532 30530 16544
rect 30561 16541 30573 16544
rect 30607 16572 30619 16575
rect 30650 16572 30656 16584
rect 30607 16544 30656 16572
rect 30607 16541 30619 16544
rect 30561 16535 30619 16541
rect 30650 16532 30656 16544
rect 30708 16532 30714 16584
rect 30745 16575 30803 16581
rect 30745 16541 30757 16575
rect 30791 16572 30803 16575
rect 31846 16572 31852 16584
rect 30791 16544 31852 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 31846 16532 31852 16544
rect 31904 16532 31910 16584
rect 32214 16532 32220 16584
rect 32272 16572 32278 16584
rect 33152 16581 33180 16680
rect 33502 16668 33508 16680
rect 33560 16668 33566 16720
rect 33594 16668 33600 16720
rect 33652 16668 33658 16720
rect 34514 16708 34520 16720
rect 34348 16680 34520 16708
rect 33612 16640 33640 16668
rect 33336 16612 33640 16640
rect 33336 16581 33364 16612
rect 34348 16581 34376 16680
rect 34514 16668 34520 16680
rect 34572 16708 34578 16720
rect 34572 16680 35572 16708
rect 34572 16668 34578 16680
rect 34793 16643 34851 16649
rect 34793 16640 34805 16643
rect 34440 16612 34805 16640
rect 32401 16575 32459 16581
rect 32401 16572 32413 16575
rect 32272 16544 32413 16572
rect 32272 16532 32278 16544
rect 32401 16541 32413 16544
rect 32447 16572 32459 16575
rect 33137 16575 33195 16581
rect 32447 16544 33088 16572
rect 32447 16541 32459 16544
rect 32401 16535 32459 16541
rect 30392 16476 30696 16504
rect 30156 16408 30328 16436
rect 30156 16396 30162 16408
rect 30558 16396 30564 16448
rect 30616 16436 30622 16448
rect 30668 16445 30696 16476
rect 30834 16464 30840 16516
rect 30892 16504 30898 16516
rect 32950 16504 32956 16516
rect 30892 16476 32956 16504
rect 30892 16464 30898 16476
rect 32950 16464 32956 16476
rect 33008 16464 33014 16516
rect 30653 16439 30711 16445
rect 30653 16436 30665 16439
rect 30616 16408 30665 16436
rect 30616 16396 30622 16408
rect 30653 16405 30665 16408
rect 30699 16436 30711 16439
rect 31478 16436 31484 16448
rect 30699 16408 31484 16436
rect 30699 16405 30711 16408
rect 30653 16399 30711 16405
rect 31478 16396 31484 16408
rect 31536 16396 31542 16448
rect 33060 16436 33088 16544
rect 33137 16541 33149 16575
rect 33183 16541 33195 16575
rect 33137 16535 33195 16541
rect 33321 16575 33379 16581
rect 33321 16541 33333 16575
rect 33367 16541 33379 16575
rect 33321 16535 33379 16541
rect 34333 16575 34391 16581
rect 34333 16541 34345 16575
rect 34379 16541 34391 16575
rect 34333 16535 34391 16541
rect 33152 16504 33180 16535
rect 34440 16504 34468 16612
rect 34793 16609 34805 16612
rect 34839 16609 34851 16643
rect 34793 16603 34851 16609
rect 34517 16575 34575 16581
rect 34517 16541 34529 16575
rect 34563 16541 34575 16575
rect 34517 16535 34575 16541
rect 33152 16476 34468 16504
rect 34532 16504 34560 16535
rect 34698 16532 34704 16584
rect 34756 16572 34762 16584
rect 35544 16581 35572 16680
rect 38856 16640 38884 16736
rect 39040 16640 39068 16736
rect 38856 16612 38976 16640
rect 39040 16612 39344 16640
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34756 16544 34897 16572
rect 34756 16532 34762 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35529 16575 35587 16581
rect 35529 16541 35541 16575
rect 35575 16541 35587 16575
rect 38948 16572 38976 16612
rect 39316 16581 39344 16612
rect 39942 16600 39948 16652
rect 40000 16640 40006 16652
rect 40957 16643 41015 16649
rect 40957 16640 40969 16643
rect 40000 16612 40969 16640
rect 40000 16600 40006 16612
rect 40957 16609 40969 16612
rect 41003 16640 41015 16643
rect 42518 16640 42524 16652
rect 41003 16612 42524 16640
rect 41003 16609 41015 16612
rect 40957 16603 41015 16609
rect 42518 16600 42524 16612
rect 42576 16600 42582 16652
rect 39117 16575 39175 16581
rect 39117 16572 39129 16575
rect 38948 16544 39129 16572
rect 35529 16535 35587 16541
rect 39117 16541 39129 16544
rect 39163 16541 39175 16575
rect 39117 16535 39175 16541
rect 39301 16575 39359 16581
rect 39301 16541 39313 16575
rect 39347 16541 39359 16575
rect 39301 16535 39359 16541
rect 35345 16507 35403 16513
rect 35345 16504 35357 16507
rect 34532 16476 35357 16504
rect 33778 16436 33784 16448
rect 33060 16408 33784 16436
rect 33778 16396 33784 16408
rect 33836 16396 33842 16448
rect 33870 16396 33876 16448
rect 33928 16436 33934 16448
rect 35268 16445 35296 16476
rect 35345 16473 35357 16476
rect 35391 16473 35403 16507
rect 35345 16467 35403 16473
rect 37458 16464 37464 16516
rect 37516 16504 37522 16516
rect 40405 16507 40463 16513
rect 40405 16504 40417 16507
rect 37516 16476 40417 16504
rect 37516 16464 37522 16476
rect 40405 16473 40417 16476
rect 40451 16473 40463 16507
rect 40405 16467 40463 16473
rect 41233 16507 41291 16513
rect 41233 16473 41245 16507
rect 41279 16504 41291 16507
rect 41506 16504 41512 16516
rect 41279 16476 41512 16504
rect 41279 16473 41291 16476
rect 41233 16467 41291 16473
rect 41506 16464 41512 16476
rect 41564 16464 41570 16516
rect 42242 16464 42248 16516
rect 42300 16464 42306 16516
rect 34333 16439 34391 16445
rect 34333 16436 34345 16439
rect 33928 16408 34345 16436
rect 33928 16396 33934 16408
rect 34333 16405 34345 16408
rect 34379 16405 34391 16439
rect 34333 16399 34391 16405
rect 35253 16439 35311 16445
rect 35253 16405 35265 16439
rect 35299 16436 35311 16439
rect 35299 16408 35333 16436
rect 35299 16405 35311 16408
rect 35253 16399 35311 16405
rect 35710 16396 35716 16448
rect 35768 16396 35774 16448
rect 1104 16346 44620 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 44620 16346
rect 1104 16272 44620 16294
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16232 2651 16235
rect 2774 16232 2780 16244
rect 2639 16204 2780 16232
rect 2639 16201 2651 16204
rect 2593 16195 2651 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 4706 16232 4712 16244
rect 3988 16204 4712 16232
rect 3988 16164 4016 16204
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 9582 16232 9588 16244
rect 9232 16204 9588 16232
rect 3634 16136 4016 16164
rect 4065 16167 4123 16173
rect 4065 16133 4077 16167
rect 4111 16164 4123 16167
rect 4801 16167 4859 16173
rect 4801 16164 4813 16167
rect 4111 16136 4813 16164
rect 4111 16133 4123 16136
rect 4065 16127 4123 16133
rect 4801 16133 4813 16136
rect 4847 16133 4859 16167
rect 4801 16127 4859 16133
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 9232 16173 9260 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11756 16204 11897 16232
rect 11756 16192 11762 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16201 12311 16235
rect 12253 16195 12311 16201
rect 12621 16235 12679 16241
rect 12621 16201 12633 16235
rect 12667 16232 12679 16235
rect 13078 16232 13084 16244
rect 12667 16204 13084 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 9217 16167 9275 16173
rect 6604 16136 7498 16164
rect 6604 16124 6610 16136
rect 9217 16133 9229 16167
rect 9263 16133 9275 16167
rect 9217 16127 9275 16133
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 9674 16164 9680 16176
rect 9364 16136 9680 16164
rect 9364 16124 9370 16136
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5776 16068 5917 16096
rect 5776 16056 5782 16068
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 5905 16059 5963 16065
rect 8404 16068 8861 16096
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 3326 15852 3332 15904
rect 3384 15892 3390 15904
rect 4356 15892 4384 15991
rect 5350 15988 5356 16040
rect 5408 15988 5414 16040
rect 5994 15988 6000 16040
rect 6052 16028 6058 16040
rect 7055 16031 7113 16037
rect 7055 16028 7067 16031
rect 6052 16000 7067 16028
rect 6052 15988 6058 16000
rect 7055 15997 7067 16000
rect 7101 15997 7113 16031
rect 7055 15991 7113 15997
rect 8294 15988 8300 16040
rect 8352 16028 8358 16040
rect 8404 16028 8432 16068
rect 8849 16065 8861 16068
rect 8895 16096 8907 16099
rect 8941 16099 8999 16105
rect 8941 16096 8953 16099
rect 8895 16068 8953 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 8941 16065 8953 16068
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12268 16096 12296 16195
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 16632 16204 16681 16232
rect 16632 16192 16638 16204
rect 16669 16201 16681 16204
rect 16715 16201 16727 16235
rect 16669 16195 16727 16201
rect 17129 16235 17187 16241
rect 17129 16201 17141 16235
rect 17175 16201 17187 16235
rect 17129 16195 17187 16201
rect 15470 16164 15476 16176
rect 12452 16136 13308 16164
rect 14766 16136 15476 16164
rect 12452 16108 12480 16136
rect 12115 16068 12296 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12434 16056 12440 16108
rect 12492 16056 12498 16108
rect 13280 16105 13308 16136
rect 15470 16124 15476 16136
rect 15528 16124 15534 16176
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 17144 16096 17172 16195
rect 17494 16192 17500 16244
rect 17552 16192 17558 16244
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 18380 16204 19441 16232
rect 18380 16192 18386 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 23750 16192 23756 16244
rect 23808 16192 23814 16244
rect 24486 16192 24492 16244
rect 24544 16232 24550 16244
rect 26878 16232 26884 16244
rect 24544 16204 26884 16232
rect 24544 16192 24550 16204
rect 26878 16192 26884 16204
rect 26936 16192 26942 16244
rect 31389 16235 31447 16241
rect 31389 16201 31401 16235
rect 31435 16232 31447 16235
rect 31846 16232 31852 16244
rect 31435 16204 31852 16232
rect 31435 16201 31447 16204
rect 31389 16195 31447 16201
rect 31846 16192 31852 16204
rect 31904 16192 31910 16244
rect 32950 16192 32956 16244
rect 33008 16232 33014 16244
rect 33008 16204 33180 16232
rect 33008 16192 33014 16204
rect 17589 16167 17647 16173
rect 17589 16133 17601 16167
rect 17635 16164 17647 16167
rect 17954 16164 17960 16176
rect 17635 16136 17960 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 17954 16124 17960 16136
rect 18012 16124 18018 16176
rect 23768 16164 23796 16192
rect 23492 16136 23796 16164
rect 25501 16167 25559 16173
rect 23492 16108 23520 16136
rect 25501 16133 25513 16167
rect 25547 16164 25559 16167
rect 25682 16164 25688 16176
rect 25547 16136 25688 16164
rect 25547 16133 25559 16136
rect 25501 16127 25559 16133
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 29270 16124 29276 16176
rect 29328 16164 29334 16176
rect 29641 16167 29699 16173
rect 29641 16164 29653 16167
rect 29328 16136 29653 16164
rect 29328 16124 29334 16136
rect 29641 16133 29653 16136
rect 29687 16164 29699 16167
rect 30834 16164 30840 16176
rect 29687 16136 30840 16164
rect 29687 16133 29699 16136
rect 29641 16127 29699 16133
rect 30834 16124 30840 16136
rect 30892 16124 30898 16176
rect 33152 16173 33180 16204
rect 35710 16192 35716 16244
rect 35768 16192 35774 16244
rect 42518 16192 42524 16244
rect 42576 16192 42582 16244
rect 30929 16167 30987 16173
rect 30929 16133 30941 16167
rect 30975 16133 30987 16167
rect 30929 16127 30987 16133
rect 33137 16167 33195 16173
rect 33137 16133 33149 16167
rect 33183 16164 33195 16167
rect 35728 16164 35756 16192
rect 42245 16167 42303 16173
rect 33183 16136 33456 16164
rect 33183 16133 33195 16136
rect 33137 16127 33195 16133
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 16899 16068 17172 16096
rect 17236 16068 18153 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 8352 16000 8432 16028
rect 8481 16031 8539 16037
rect 8352 15988 8358 16000
rect 8481 15997 8493 16031
rect 8527 16028 8539 16031
rect 8662 16028 8668 16040
rect 8527 16000 8668 16028
rect 8527 15997 8539 16000
rect 8481 15991 8539 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 12710 15988 12716 16040
rect 12768 15988 12774 16040
rect 12894 15988 12900 16040
rect 12952 15988 12958 16040
rect 13538 15988 13544 16040
rect 13596 15988 13602 16040
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15059 16000 15669 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 17236 16028 17264 16068
rect 18141 16065 18153 16068
rect 18187 16096 18199 16099
rect 18782 16096 18788 16108
rect 18187 16068 18788 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 18782 16056 18788 16068
rect 18840 16096 18846 16108
rect 21818 16096 21824 16108
rect 18840 16068 21824 16096
rect 18840 16056 18846 16068
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 26694 16096 26700 16108
rect 24886 16068 26700 16096
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 26970 16056 26976 16108
rect 27028 16056 27034 16108
rect 29457 16099 29515 16105
rect 29457 16065 29469 16099
rect 29503 16065 29515 16099
rect 29457 16059 29515 16065
rect 16356 16000 17264 16028
rect 16356 15988 16362 16000
rect 17678 15988 17684 16040
rect 17736 15988 17742 16040
rect 20070 15988 20076 16040
rect 20128 16028 20134 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20128 16000 20545 16028
rect 20128 15988 20134 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 23842 16028 23848 16040
rect 23799 16000 23848 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 22646 15920 22652 15972
rect 22704 15960 22710 15972
rect 22922 15960 22928 15972
rect 22704 15932 22928 15960
rect 22704 15920 22710 15932
rect 22922 15920 22928 15932
rect 22980 15920 22986 15972
rect 29086 15960 29092 15972
rect 27080 15932 29092 15960
rect 3384 15864 4384 15892
rect 5537 15895 5595 15901
rect 3384 15852 3390 15864
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 5626 15892 5632 15904
rect 5583 15864 5632 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 13630 15892 13636 15904
rect 10735 15864 13636 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 15102 15852 15108 15904
rect 15160 15852 15166 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 27080 15892 27108 15932
rect 29086 15920 29092 15932
rect 29144 15920 29150 15972
rect 22520 15864 27108 15892
rect 27157 15895 27215 15901
rect 22520 15852 22526 15864
rect 27157 15861 27169 15895
rect 27203 15892 27215 15895
rect 27246 15892 27252 15904
rect 27203 15864 27252 15892
rect 27203 15861 27215 15864
rect 27157 15855 27215 15861
rect 27246 15852 27252 15864
rect 27304 15852 27310 15904
rect 29270 15852 29276 15904
rect 29328 15852 29334 15904
rect 29472 15892 29500 16059
rect 29546 16056 29552 16108
rect 29604 16056 29610 16108
rect 29779 16099 29837 16105
rect 29779 16065 29791 16099
rect 29825 16096 29837 16099
rect 30282 16096 30288 16108
rect 29825 16068 30288 16096
rect 29825 16065 29837 16068
rect 29779 16059 29837 16065
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 30944 16096 30972 16127
rect 30852 16068 30972 16096
rect 31094 16099 31152 16105
rect 30852 16040 30880 16068
rect 31094 16065 31106 16099
rect 31140 16096 31152 16099
rect 31195 16099 31253 16105
rect 31140 16086 31156 16096
rect 31195 16086 31207 16099
rect 31140 16065 31207 16086
rect 31241 16065 31253 16099
rect 31094 16059 31253 16065
rect 31128 16058 31248 16059
rect 29638 15988 29644 16040
rect 29696 15988 29702 16040
rect 29917 16031 29975 16037
rect 29917 15997 29929 16031
rect 29963 16028 29975 16031
rect 30009 16031 30067 16037
rect 30009 16028 30021 16031
rect 29963 16000 30021 16028
rect 29963 15997 29975 16000
rect 29917 15991 29975 15997
rect 30009 15997 30021 16000
rect 30055 15997 30067 16031
rect 30009 15991 30067 15997
rect 30098 15988 30104 16040
rect 30156 16028 30162 16040
rect 30561 16031 30619 16037
rect 30561 16028 30573 16031
rect 30156 16000 30573 16028
rect 30156 15988 30162 16000
rect 30561 15997 30573 16000
rect 30607 15997 30619 16031
rect 30561 15991 30619 15997
rect 30650 15988 30656 16040
rect 30708 16028 30714 16040
rect 30745 16031 30803 16037
rect 30745 16028 30757 16031
rect 30708 16000 30757 16028
rect 30708 15988 30714 16000
rect 30745 15997 30757 16000
rect 30791 15997 30803 16031
rect 30745 15991 30803 15997
rect 30834 15988 30840 16040
rect 30892 15988 30898 16040
rect 31128 16028 31156 16058
rect 31294 16056 31300 16108
rect 31352 16096 31358 16108
rect 31389 16099 31447 16105
rect 31389 16096 31401 16099
rect 31352 16068 31401 16096
rect 31352 16056 31358 16068
rect 31389 16065 31401 16068
rect 31435 16065 31447 16099
rect 31389 16059 31447 16065
rect 31478 16056 31484 16108
rect 31536 16056 31542 16108
rect 31665 16099 31723 16105
rect 31665 16096 31677 16099
rect 31588 16068 31677 16096
rect 31588 16040 31616 16068
rect 31665 16065 31677 16068
rect 31711 16065 31723 16099
rect 31665 16059 31723 16065
rect 31941 16099 31999 16105
rect 31941 16065 31953 16099
rect 31987 16096 31999 16099
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 31987 16068 32137 16096
rect 31987 16065 31999 16068
rect 31941 16059 31999 16065
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 30944 16000 31156 16028
rect 29656 15960 29684 15988
rect 30944 15960 30972 16000
rect 31570 15988 31576 16040
rect 31628 15988 31634 16040
rect 31956 16028 31984 16059
rect 32214 16056 32220 16108
rect 32272 16096 32278 16108
rect 33019 16099 33077 16105
rect 33019 16096 33031 16099
rect 32272 16068 33031 16096
rect 32272 16056 32278 16068
rect 33019 16065 33031 16068
rect 33065 16065 33077 16099
rect 33019 16059 33077 16065
rect 31726 16000 31984 16028
rect 32769 16031 32827 16037
rect 29656 15932 30972 15960
rect 31018 15920 31024 15972
rect 31076 15960 31082 15972
rect 31726 15960 31754 16000
rect 32769 15997 32781 16031
rect 32815 16028 32827 16031
rect 32861 16031 32919 16037
rect 32861 16028 32873 16031
rect 32815 16000 32873 16028
rect 32815 15997 32827 16000
rect 32769 15991 32827 15997
rect 32861 15997 32873 16000
rect 32907 15997 32919 16031
rect 32861 15991 32919 15997
rect 31076 15932 31754 15960
rect 31076 15920 31082 15932
rect 31846 15920 31852 15972
rect 31904 15920 31910 15972
rect 33034 15960 33062 16059
rect 33226 16056 33232 16108
rect 33284 16056 33290 16108
rect 33318 16056 33324 16108
rect 33376 16056 33382 16108
rect 33428 16028 33456 16136
rect 33796 16136 35756 16164
rect 39868 16136 41414 16164
rect 33796 16105 33824 16136
rect 33781 16099 33839 16105
rect 33781 16065 33793 16099
rect 33827 16065 33839 16099
rect 33781 16059 33839 16065
rect 33870 16056 33876 16108
rect 33928 16056 33934 16108
rect 33965 16099 34023 16105
rect 33965 16065 33977 16099
rect 34011 16065 34023 16099
rect 33965 16059 34023 16065
rect 33980 16028 34008 16059
rect 34054 16056 34060 16108
rect 34112 16105 34118 16108
rect 39868 16105 39896 16136
rect 34112 16099 34141 16105
rect 34129 16065 34141 16099
rect 34112 16059 34141 16065
rect 39853 16099 39911 16105
rect 39853 16065 39865 16099
rect 39899 16065 39911 16099
rect 39853 16059 39911 16065
rect 34112 16056 34118 16059
rect 40494 16056 40500 16108
rect 40552 16056 40558 16108
rect 41386 16096 41414 16136
rect 42245 16133 42257 16167
rect 42291 16164 42303 16167
rect 42536 16164 42564 16192
rect 42291 16136 42564 16164
rect 42291 16133 42303 16136
rect 42245 16127 42303 16133
rect 42429 16099 42487 16105
rect 42429 16096 42441 16099
rect 41386 16068 42441 16096
rect 42429 16065 42441 16068
rect 42475 16065 42487 16099
rect 42429 16059 42487 16065
rect 43990 16056 43996 16108
rect 44048 16056 44054 16108
rect 33428 16000 34008 16028
rect 34072 15960 34100 16056
rect 34241 16031 34299 16037
rect 34241 15997 34253 16031
rect 34287 16028 34299 16031
rect 34333 16031 34391 16037
rect 34333 16028 34345 16031
rect 34287 16000 34345 16028
rect 34287 15997 34299 16000
rect 34241 15991 34299 15997
rect 34333 15997 34345 16000
rect 34379 15997 34391 16031
rect 34333 15991 34391 15997
rect 34606 15988 34612 16040
rect 34664 16028 34670 16040
rect 34885 16031 34943 16037
rect 34885 16028 34897 16031
rect 34664 16000 34897 16028
rect 34664 15988 34670 16000
rect 34885 15997 34897 16000
rect 34931 15997 34943 16031
rect 34885 15991 34943 15997
rect 39758 15988 39764 16040
rect 39816 16028 39822 16040
rect 39945 16031 40003 16037
rect 39945 16028 39957 16031
rect 39816 16000 39957 16028
rect 39816 15988 39822 16000
rect 39945 15997 39957 16000
rect 39991 16028 40003 16031
rect 41598 16028 41604 16040
rect 39991 16000 41604 16028
rect 39991 15997 40003 16000
rect 39945 15991 40003 15997
rect 41598 15988 41604 16000
rect 41656 15988 41662 16040
rect 42150 15988 42156 16040
rect 42208 16028 42214 16040
rect 42981 16031 43039 16037
rect 42981 16028 42993 16031
rect 42208 16000 42993 16028
rect 42208 15988 42214 16000
rect 42981 15997 42993 16000
rect 43027 15997 43039 16031
rect 42981 15991 43039 15997
rect 33034 15932 34100 15960
rect 31573 15895 31631 15901
rect 31573 15892 31585 15895
rect 29472 15864 31585 15892
rect 31573 15861 31585 15864
rect 31619 15861 31631 15895
rect 31573 15855 31631 15861
rect 33502 15852 33508 15904
rect 33560 15852 33566 15904
rect 33594 15852 33600 15904
rect 33652 15852 33658 15904
rect 40218 15852 40224 15904
rect 40276 15852 40282 15904
rect 44174 15852 44180 15904
rect 44232 15852 44238 15904
rect 1104 15802 44620 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 44620 15802
rect 1104 15728 44620 15750
rect 5350 15648 5356 15700
rect 5408 15697 5414 15700
rect 5408 15691 5457 15697
rect 5408 15657 5411 15691
rect 5445 15657 5457 15691
rect 5408 15651 5457 15657
rect 5408 15648 5414 15651
rect 5994 15648 6000 15700
rect 6052 15648 6058 15700
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11848 15660 11989 15688
rect 11848 15648 11854 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 11977 15651 12035 15657
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13725 15691 13783 15697
rect 13725 15688 13737 15691
rect 13596 15660 13737 15688
rect 13596 15648 13602 15660
rect 13725 15657 13737 15660
rect 13771 15657 13783 15691
rect 22462 15688 22468 15700
rect 13725 15651 13783 15657
rect 13832 15660 22468 15688
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 3326 15552 3332 15564
rect 1903 15524 3332 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15552 3663 15555
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 3651 15524 4353 15552
rect 3651 15521 3663 15524
rect 3605 15515 3663 15521
rect 4341 15521 4353 15524
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15552 5319 15555
rect 6012 15552 6040 15648
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 13832 15620 13860 15660
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23106 15688 23112 15700
rect 22572 15660 23112 15688
rect 21821 15623 21879 15629
rect 13688 15592 13860 15620
rect 17696 15592 18920 15620
rect 13688 15580 13694 15592
rect 17696 15564 17724 15592
rect 5307 15524 6040 15552
rect 5307 15521 5319 15524
rect 5261 15515 5319 15521
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 7193 15555 7251 15561
rect 7193 15552 7205 15555
rect 7064 15524 7205 15552
rect 7064 15512 7070 15524
rect 7193 15521 7205 15524
rect 7239 15552 7251 15555
rect 8294 15552 8300 15564
rect 7239 15524 8300 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 8294 15512 8300 15524
rect 8352 15552 8358 15564
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 8352 15524 10241 15552
rect 8352 15512 8358 15524
rect 10229 15521 10241 15524
rect 10275 15521 10287 15555
rect 10229 15515 10287 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12894 15552 12900 15564
rect 12759 15524 12900 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12894 15512 12900 15524
rect 12952 15552 12958 15564
rect 14645 15555 14703 15561
rect 14645 15552 14657 15555
rect 12952 15524 14657 15552
rect 12952 15512 12958 15524
rect 14645 15521 14657 15524
rect 14691 15552 14703 15555
rect 17678 15552 17684 15564
rect 14691 15524 17684 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 18322 15512 18328 15564
rect 18380 15552 18386 15564
rect 18892 15552 18920 15592
rect 21821 15589 21833 15623
rect 21867 15620 21879 15623
rect 22572 15620 22600 15660
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 26510 15648 26516 15700
rect 26568 15648 26574 15700
rect 26697 15691 26755 15697
rect 26697 15657 26709 15691
rect 26743 15688 26755 15691
rect 26970 15688 26976 15700
rect 26743 15660 26976 15688
rect 26743 15657 26755 15660
rect 26697 15651 26755 15657
rect 26970 15648 26976 15660
rect 27028 15648 27034 15700
rect 29270 15648 29276 15700
rect 29328 15648 29334 15700
rect 29365 15691 29423 15697
rect 29365 15657 29377 15691
rect 29411 15688 29423 15691
rect 30098 15688 30104 15700
rect 29411 15660 30104 15688
rect 29411 15657 29423 15660
rect 29365 15651 29423 15657
rect 30098 15648 30104 15660
rect 30156 15648 30162 15700
rect 30561 15691 30619 15697
rect 30561 15657 30573 15691
rect 30607 15688 30619 15691
rect 31018 15688 31024 15700
rect 30607 15660 31024 15688
rect 30607 15657 30619 15660
rect 30561 15651 30619 15657
rect 31018 15648 31024 15660
rect 31076 15648 31082 15700
rect 31294 15648 31300 15700
rect 31352 15688 31358 15700
rect 32861 15691 32919 15697
rect 31352 15660 32812 15688
rect 31352 15648 31358 15660
rect 21867 15592 22600 15620
rect 26528 15620 26556 15648
rect 26789 15623 26847 15629
rect 26789 15620 26801 15623
rect 26528 15592 26801 15620
rect 21867 15589 21879 15592
rect 21821 15583 21879 15589
rect 26789 15589 26801 15592
rect 26835 15589 26847 15623
rect 26789 15583 26847 15589
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 18380 15524 18828 15552
rect 18892 15524 19901 15552
rect 18380 15512 18386 15524
rect 3266 15456 4752 15484
rect 4724 15428 4752 15456
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6788 15456 6837 15484
rect 6788 15444 6794 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 12400 15456 12449 15484
rect 12400 15444 12406 15456
rect 12437 15453 12449 15456
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 14461 15487 14519 15493
rect 13955 15456 14136 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 2133 15419 2191 15425
rect 2133 15385 2145 15419
rect 2179 15385 2191 15419
rect 2133 15379 2191 15385
rect 3712 15388 4660 15416
rect 2148 15348 2176 15379
rect 3712 15348 3740 15388
rect 2148 15320 3740 15348
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 4632 15357 4660 15388
rect 4706 15376 4712 15428
rect 4764 15416 4770 15428
rect 4764 15388 5842 15416
rect 4764 15376 4770 15388
rect 10502 15376 10508 15428
rect 10560 15376 10566 15428
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15317 4675 15351
rect 4617 15311 4675 15317
rect 12066 15308 12072 15360
rect 12124 15308 12130 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 14108 15357 14136 15456
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 15102 15484 15108 15496
rect 14507 15456 15108 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15453 18751 15487
rect 18800 15484 18828 15524
rect 19889 15521 19901 15524
rect 19935 15552 19947 15555
rect 20346 15552 20352 15564
rect 19935 15524 20352 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 21542 15552 21548 15564
rect 20496 15524 21548 15552
rect 20496 15512 20502 15524
rect 20073 15487 20131 15493
rect 20073 15484 20085 15487
rect 18800 15456 20085 15484
rect 18693 15447 18751 15453
rect 20073 15453 20085 15456
rect 20119 15453 20131 15487
rect 21468 15470 21496 15524
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 22465 15555 22523 15561
rect 22465 15521 22477 15555
rect 22511 15552 22523 15555
rect 23474 15552 23480 15564
rect 22511 15524 23480 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15552 24271 15555
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 24259 15524 24409 15552
rect 24259 15521 24271 15524
rect 24213 15515 24271 15521
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 26145 15555 26203 15561
rect 26145 15521 26157 15555
rect 26191 15552 26203 15555
rect 26602 15552 26608 15564
rect 26191 15524 26608 15552
rect 26191 15521 26203 15524
rect 26145 15515 26203 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 27617 15555 27675 15561
rect 27617 15521 27629 15555
rect 27663 15521 27675 15555
rect 27617 15515 27675 15521
rect 27893 15555 27951 15561
rect 27893 15521 27905 15555
rect 27939 15552 27951 15555
rect 29288 15552 29316 15648
rect 32784 15620 32812 15660
rect 32861 15657 32873 15691
rect 32907 15688 32919 15691
rect 33226 15688 33232 15700
rect 32907 15660 33232 15688
rect 32907 15657 32919 15660
rect 32861 15651 32919 15657
rect 33226 15648 33232 15660
rect 33284 15648 33290 15700
rect 33318 15648 33324 15700
rect 33376 15688 33382 15700
rect 33505 15691 33563 15697
rect 33505 15688 33517 15691
rect 33376 15660 33517 15688
rect 33376 15648 33382 15660
rect 33505 15657 33517 15660
rect 33551 15657 33563 15691
rect 33505 15651 33563 15657
rect 33778 15648 33784 15700
rect 33836 15688 33842 15700
rect 34241 15691 34299 15697
rect 34241 15688 34253 15691
rect 33836 15660 34253 15688
rect 33836 15648 33842 15660
rect 34241 15657 34253 15660
rect 34287 15657 34299 15691
rect 38010 15688 38016 15700
rect 34241 15651 34299 15657
rect 37936 15660 38016 15688
rect 36265 15623 36323 15629
rect 36265 15620 36277 15623
rect 32784 15592 36277 15620
rect 36265 15589 36277 15592
rect 36311 15589 36323 15623
rect 36265 15583 36323 15589
rect 27939 15524 29316 15552
rect 32033 15555 32091 15561
rect 27939 15521 27951 15524
rect 27893 15515 27951 15521
rect 32033 15521 32045 15555
rect 32079 15552 32091 15555
rect 33502 15552 33508 15564
rect 32079 15524 33508 15552
rect 32079 15521 32091 15524
rect 32033 15515 32091 15521
rect 20073 15447 20131 15453
rect 18708 15416 18736 15447
rect 22186 15444 22192 15496
rect 22244 15444 22250 15496
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26510 15484 26516 15496
rect 26384 15456 26516 15484
rect 26384 15444 26390 15456
rect 26510 15444 26516 15456
rect 26568 15484 26574 15496
rect 27341 15487 27399 15493
rect 27341 15484 27353 15487
rect 26568 15456 27353 15484
rect 26568 15444 26574 15456
rect 27341 15453 27353 15456
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 19613 15419 19671 15425
rect 18708 15388 19288 15416
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 12492 15320 12541 15348
rect 12492 15308 12498 15320
rect 12529 15317 12541 15320
rect 12575 15317 12587 15351
rect 12529 15311 12587 15317
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14550 15308 14556 15360
rect 14608 15308 14614 15360
rect 18506 15308 18512 15360
rect 18564 15308 18570 15360
rect 19260 15357 19288 15388
rect 19613 15385 19625 15419
rect 19659 15416 19671 15419
rect 19978 15416 19984 15428
rect 19659 15388 19984 15416
rect 19659 15385 19671 15388
rect 19613 15379 19671 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 20346 15376 20352 15428
rect 20404 15376 20410 15428
rect 22741 15419 22799 15425
rect 22741 15416 22753 15419
rect 22572 15388 22753 15416
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15317 19303 15351
rect 19245 15311 19303 15317
rect 19705 15351 19763 15357
rect 19705 15317 19717 15351
rect 19751 15348 19763 15351
rect 20162 15348 20168 15360
rect 19751 15320 20168 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 22373 15351 22431 15357
rect 22373 15317 22385 15351
rect 22419 15348 22431 15351
rect 22572 15348 22600 15388
rect 22741 15385 22753 15388
rect 22787 15385 22799 15419
rect 22741 15379 22799 15385
rect 23198 15376 23204 15428
rect 23256 15376 23262 15428
rect 27632 15416 27660 15515
rect 33502 15512 33508 15524
rect 33560 15512 33566 15564
rect 33870 15552 33876 15564
rect 33612 15524 33876 15552
rect 29362 15484 29368 15496
rect 29026 15470 29368 15484
rect 29012 15456 29368 15470
rect 27798 15416 27804 15428
rect 27632 15388 27804 15416
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 22419 15320 22600 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 24210 15308 24216 15360
rect 24268 15348 24274 15360
rect 24670 15348 24676 15360
rect 24268 15320 24676 15348
rect 24268 15308 24274 15320
rect 24670 15308 24676 15320
rect 24728 15348 24734 15360
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 24728 15320 25053 15348
rect 24728 15308 24734 15320
rect 25041 15317 25053 15320
rect 25087 15317 25099 15351
rect 25041 15311 25099 15317
rect 26234 15308 26240 15360
rect 26292 15308 26298 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 29012 15348 29040 15456
rect 29362 15444 29368 15456
rect 29420 15484 29426 15496
rect 32309 15487 32367 15493
rect 29420 15456 30958 15484
rect 29420 15444 29426 15456
rect 32309 15453 32321 15487
rect 32355 15484 32367 15487
rect 32766 15484 32772 15496
rect 32355 15456 32772 15484
rect 32355 15453 32367 15456
rect 32309 15447 32367 15453
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 33042 15444 33048 15496
rect 33100 15444 33106 15496
rect 33612 15493 33640 15524
rect 33870 15512 33876 15524
rect 33928 15512 33934 15564
rect 34606 15552 34612 15564
rect 34348 15524 34612 15552
rect 33321 15487 33379 15493
rect 33321 15453 33333 15487
rect 33367 15484 33379 15487
rect 33597 15487 33655 15493
rect 33597 15484 33609 15487
rect 33367 15456 33609 15484
rect 33367 15453 33379 15456
rect 33321 15447 33379 15453
rect 33597 15453 33609 15456
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 33686 15444 33692 15496
rect 33744 15444 33750 15496
rect 34348 15493 34376 15524
rect 34606 15512 34612 15524
rect 34664 15512 34670 15564
rect 37737 15555 37795 15561
rect 37737 15521 37749 15555
rect 37783 15552 37795 15555
rect 37936 15552 37964 15660
rect 38010 15648 38016 15660
rect 38068 15648 38074 15700
rect 41506 15648 41512 15700
rect 41564 15688 41570 15700
rect 41969 15691 42027 15697
rect 41969 15688 41981 15691
rect 41564 15660 41981 15688
rect 41564 15648 41570 15660
rect 41969 15657 41981 15660
rect 42015 15657 42027 15691
rect 41969 15651 42027 15657
rect 42150 15648 42156 15700
rect 42208 15648 42214 15700
rect 41693 15623 41751 15629
rect 38028 15592 39988 15620
rect 38028 15564 38056 15592
rect 39960 15564 39988 15592
rect 41693 15589 41705 15623
rect 41739 15620 41751 15623
rect 42168 15620 42196 15648
rect 41739 15592 42196 15620
rect 41739 15589 41751 15592
rect 41693 15583 41751 15589
rect 37783 15524 37964 15552
rect 37783 15521 37795 15524
rect 37737 15515 37795 15521
rect 38010 15512 38016 15564
rect 38068 15512 38074 15564
rect 39114 15512 39120 15564
rect 39172 15552 39178 15564
rect 39209 15555 39267 15561
rect 39209 15552 39221 15555
rect 39172 15524 39221 15552
rect 39172 15512 39178 15524
rect 39209 15521 39221 15524
rect 39255 15521 39267 15555
rect 39209 15515 39267 15521
rect 39942 15512 39948 15564
rect 40000 15512 40006 15564
rect 40218 15512 40224 15564
rect 40276 15512 40282 15564
rect 42518 15512 42524 15564
rect 42576 15512 42582 15564
rect 34333 15487 34391 15493
rect 34333 15453 34345 15487
rect 34379 15453 34391 15487
rect 34333 15447 34391 15453
rect 35342 15444 35348 15496
rect 35400 15444 35406 15496
rect 35529 15487 35587 15493
rect 35529 15453 35541 15487
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 38841 15487 38899 15493
rect 38841 15453 38853 15487
rect 38887 15484 38899 15487
rect 38887 15456 38976 15484
rect 38887 15453 38899 15456
rect 38841 15447 38899 15453
rect 33060 15416 33088 15444
rect 33413 15419 33471 15425
rect 33413 15416 33425 15419
rect 33060 15388 33425 15416
rect 33413 15385 33425 15388
rect 33459 15385 33471 15419
rect 33413 15379 33471 15385
rect 27580 15320 29040 15348
rect 33229 15351 33287 15357
rect 27580 15308 27586 15320
rect 33229 15317 33241 15351
rect 33275 15348 33287 15351
rect 33704 15348 33732 15444
rect 33275 15320 33732 15348
rect 33275 15317 33287 15320
rect 33229 15311 33287 15317
rect 35434 15308 35440 15360
rect 35492 15308 35498 15360
rect 35544 15348 35572 15447
rect 37182 15376 37188 15428
rect 37240 15376 37246 15428
rect 38102 15348 38108 15360
rect 35544 15320 38108 15348
rect 38102 15308 38108 15320
rect 38160 15308 38166 15360
rect 38194 15308 38200 15360
rect 38252 15308 38258 15360
rect 38948 15357 38976 15456
rect 39298 15444 39304 15496
rect 39356 15484 39362 15496
rect 39574 15484 39580 15496
rect 39356 15456 39580 15484
rect 39356 15444 39362 15456
rect 39574 15444 39580 15456
rect 39632 15444 39638 15496
rect 41598 15444 41604 15496
rect 41656 15484 41662 15496
rect 41785 15487 41843 15493
rect 41785 15484 41797 15487
rect 41656 15456 41797 15484
rect 41656 15444 41662 15456
rect 41785 15453 41797 15456
rect 41831 15453 41843 15487
rect 41785 15447 41843 15453
rect 41969 15487 42027 15493
rect 41969 15453 41981 15487
rect 42015 15484 42027 15487
rect 42058 15484 42064 15496
rect 42015 15456 42064 15484
rect 42015 15453 42027 15456
rect 41969 15447 42027 15453
rect 42058 15444 42064 15456
rect 42116 15444 42122 15496
rect 40862 15376 40868 15428
rect 40920 15376 40926 15428
rect 42794 15376 42800 15428
rect 42852 15376 42858 15428
rect 43346 15376 43352 15428
rect 43404 15376 43410 15428
rect 38933 15351 38991 15357
rect 38933 15317 38945 15351
rect 38979 15317 38991 15351
rect 38933 15311 38991 15317
rect 44266 15308 44272 15360
rect 44324 15308 44330 15360
rect 1104 15258 44620 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 44620 15258
rect 1104 15184 44620 15206
rect 5905 15147 5963 15153
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 6730 15144 6736 15156
rect 5951 15116 6736 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 10502 15104 10508 15156
rect 10560 15144 10566 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 10560 15116 10885 15144
rect 10560 15104 10566 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 10873 15107 10931 15113
rect 12066 15104 12072 15156
rect 12124 15104 12130 15156
rect 18322 15104 18328 15156
rect 18380 15104 18386 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20070 15144 20076 15156
rect 19659 15116 20076 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20533 15147 20591 15153
rect 20533 15144 20545 15147
rect 20404 15116 20545 15144
rect 20404 15104 20410 15116
rect 20533 15113 20545 15116
rect 20579 15113 20591 15147
rect 20533 15107 20591 15113
rect 20901 15147 20959 15153
rect 20901 15113 20913 15147
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 3697 15079 3755 15085
rect 3697 15045 3709 15079
rect 3743 15076 3755 15079
rect 3786 15076 3792 15088
rect 3743 15048 3792 15076
rect 3743 15045 3755 15048
rect 3697 15039 3755 15045
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 9030 15036 9036 15088
rect 9088 15036 9094 15088
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 3326 14968 3332 15020
rect 3384 15008 3390 15020
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3384 14980 3433 15008
rect 3384 14968 3390 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 4764 14980 4830 15008
rect 4764 14968 4770 14980
rect 5534 14968 5540 15020
rect 5592 14968 5598 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8757 15011 8815 15017
rect 8757 15008 8769 15011
rect 8352 14980 8769 15008
rect 8352 14968 8358 14980
rect 8757 14977 8769 14980
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 12084 15008 12112 15104
rect 18340 15076 18368 15104
rect 20438 15076 20444 15088
rect 17880 15048 18368 15076
rect 19366 15048 20444 15076
rect 17880 15017 17908 15048
rect 20438 15036 20444 15048
rect 20496 15036 20502 15088
rect 11103 14980 12112 15008
rect 17865 15011 17923 15017
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 17865 14977 17877 15011
rect 17911 14977 17923 15011
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 17865 14971 17923 14977
rect 20088 14980 20361 15008
rect 20088 14952 20116 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 20916 15008 20944 15107
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21232 15116 21925 15144
rect 21232 15104 21238 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 22646 15144 22652 15156
rect 21913 15107 21971 15113
rect 22388 15116 22652 15144
rect 22097 15079 22155 15085
rect 22097 15076 22109 15079
rect 20763 14980 20944 15008
rect 21100 15048 22109 15076
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 5626 14900 5632 14952
rect 5684 14900 5690 14952
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 18141 14943 18199 14949
rect 10551 14912 17264 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 6362 14832 6368 14884
rect 6420 14872 6426 14884
rect 8754 14872 8760 14884
rect 6420 14844 8760 14872
rect 6420 14832 6426 14844
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 14182 14832 14188 14884
rect 14240 14872 14246 14884
rect 16482 14872 16488 14884
rect 14240 14844 16488 14872
rect 14240 14832 14246 14844
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 17126 14804 17132 14816
rect 12308 14776 17132 14804
rect 12308 14764 12314 14776
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 17236 14804 17264 14912
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18506 14940 18512 14952
rect 18187 14912 18512 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 18690 14900 18696 14952
rect 18748 14940 18754 14952
rect 18748 14912 19196 14940
rect 18748 14900 18754 14912
rect 19168 14872 19196 14912
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 21100 14940 21128 15048
rect 22097 15045 22109 15048
rect 22143 15076 22155 15079
rect 22388 15076 22416 15116
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 22741 15147 22799 15153
rect 22741 15113 22753 15147
rect 22787 15144 22799 15147
rect 24210 15144 24216 15156
rect 22787 15116 24216 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 35986 15144 35992 15156
rect 24964 15116 27844 15144
rect 22143 15048 22416 15076
rect 22143 15045 22155 15048
rect 22097 15039 22155 15045
rect 21266 14968 21272 15020
rect 21324 14968 21330 15020
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21468 14980 21833 15008
rect 20211 14912 21128 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21468 14872 21496 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22370 15008 22376 15020
rect 21968 14980 22376 15008
rect 21968 14968 21974 14980
rect 22370 14968 22376 14980
rect 22428 15008 22434 15020
rect 24964 15017 24992 15116
rect 27816 15088 27844 15116
rect 32784 15116 35992 15144
rect 26694 15076 26700 15088
rect 26450 15048 26700 15076
rect 26694 15036 26700 15048
rect 26752 15076 26758 15088
rect 26970 15076 26976 15088
rect 26752 15048 26976 15076
rect 26752 15036 26758 15048
rect 26970 15036 26976 15048
rect 27028 15076 27034 15088
rect 27522 15076 27528 15088
rect 27028 15048 27528 15076
rect 27028 15036 27034 15048
rect 27522 15036 27528 15048
rect 27580 15036 27586 15088
rect 27798 15036 27804 15088
rect 27856 15036 27862 15088
rect 32784 15020 32812 15116
rect 24949 15011 25007 15017
rect 22428 14980 22968 15008
rect 22428 14968 22434 14980
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14909 21603 14943
rect 21545 14903 21603 14909
rect 19168 14844 21496 14872
rect 21560 14872 21588 14903
rect 22646 14900 22652 14952
rect 22704 14940 22710 14952
rect 22940 14949 22968 14980
rect 24949 14977 24961 15011
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 26436 14980 31754 15008
rect 22833 14943 22891 14949
rect 22833 14940 22845 14943
rect 22704 14912 22845 14940
rect 22704 14900 22710 14912
rect 22833 14909 22845 14912
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 22925 14943 22983 14949
rect 22925 14909 22937 14943
rect 22971 14909 22983 14943
rect 22925 14903 22983 14909
rect 25222 14900 25228 14952
rect 25280 14900 25286 14952
rect 25314 14900 25320 14952
rect 25372 14940 25378 14952
rect 26436 14940 26464 14980
rect 25372 14912 26464 14940
rect 26697 14943 26755 14949
rect 25372 14900 25378 14912
rect 26697 14909 26709 14943
rect 26743 14940 26755 14943
rect 27525 14943 27583 14949
rect 27525 14940 27537 14943
rect 26743 14912 27537 14940
rect 26743 14909 26755 14912
rect 26697 14903 26755 14909
rect 27525 14909 27537 14912
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 21910 14872 21916 14884
rect 21560 14844 21916 14872
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 22097 14875 22155 14881
rect 22097 14872 22109 14875
rect 22060 14844 22109 14872
rect 22060 14832 22066 14844
rect 22097 14841 22109 14844
rect 22143 14841 22155 14875
rect 22097 14835 22155 14841
rect 22186 14832 22192 14884
rect 22244 14872 22250 14884
rect 22373 14875 22431 14881
rect 22373 14872 22385 14875
rect 22244 14844 22385 14872
rect 22244 14832 22250 14844
rect 22373 14841 22385 14844
rect 22419 14841 22431 14875
rect 22373 14835 22431 14841
rect 26234 14832 26240 14884
rect 26292 14872 26298 14884
rect 26973 14875 27031 14881
rect 26973 14872 26985 14875
rect 26292 14844 26985 14872
rect 26292 14832 26298 14844
rect 26973 14841 26985 14844
rect 27019 14841 27031 14875
rect 26973 14835 27031 14841
rect 31478 14804 31484 14816
rect 17236 14776 31484 14804
rect 31478 14764 31484 14776
rect 31536 14764 31542 14816
rect 31726 14804 31754 14980
rect 32766 14968 32772 15020
rect 32824 14968 32830 15020
rect 35084 15017 35112 15116
rect 35986 15104 35992 15116
rect 36044 15104 36050 15156
rect 38010 15104 38016 15156
rect 38068 15104 38074 15156
rect 39574 15104 39580 15156
rect 39632 15104 39638 15156
rect 43533 15147 43591 15153
rect 43533 15113 43545 15147
rect 43579 15144 43591 15147
rect 43990 15144 43996 15156
rect 43579 15116 43996 15144
rect 43579 15113 43591 15116
rect 43533 15107 43591 15113
rect 43990 15104 43996 15116
rect 44048 15104 44054 15156
rect 35345 15079 35403 15085
rect 35345 15045 35357 15079
rect 35391 15076 35403 15079
rect 35434 15076 35440 15088
rect 35391 15048 35440 15076
rect 35391 15045 35403 15048
rect 35345 15039 35403 15045
rect 35434 15036 35440 15048
rect 35492 15036 35498 15088
rect 38028 15076 38056 15104
rect 35069 15011 35127 15017
rect 33045 14943 33103 14949
rect 33045 14909 33057 14943
rect 33091 14940 33103 14943
rect 33594 14940 33600 14952
rect 33091 14912 33600 14940
rect 33091 14909 33103 14912
rect 33045 14903 33103 14909
rect 33594 14900 33600 14912
rect 33652 14900 33658 14952
rect 34164 14940 34192 14994
rect 35069 14977 35081 15011
rect 35115 14977 35127 15011
rect 35069 14971 35127 14977
rect 36556 14940 36584 15062
rect 37844 15048 38056 15076
rect 38105 15079 38163 15085
rect 37844 15017 37872 15048
rect 38105 15045 38117 15079
rect 38151 15076 38163 15079
rect 38194 15076 38200 15088
rect 38151 15048 38200 15076
rect 38151 15045 38163 15048
rect 38105 15039 38163 15045
rect 38194 15036 38200 15048
rect 38252 15036 38258 15088
rect 43625 15079 43683 15085
rect 43625 15076 43637 15079
rect 42996 15048 43637 15076
rect 42996 15017 43024 15048
rect 43625 15045 43637 15048
rect 43671 15045 43683 15079
rect 43625 15039 43683 15045
rect 37829 15011 37887 15017
rect 37829 14977 37841 15011
rect 37875 14977 37887 15011
rect 42981 15011 43039 15017
rect 39238 14994 41414 15008
rect 37829 14971 37887 14977
rect 39224 14980 41414 14994
rect 37182 14940 37188 14952
rect 34164 14912 37188 14940
rect 37182 14900 37188 14912
rect 37240 14940 37246 14952
rect 39224 14940 39252 14980
rect 37240 14912 39252 14940
rect 37240 14900 37246 14912
rect 34517 14875 34575 14881
rect 34517 14841 34529 14875
rect 34563 14872 34575 14875
rect 34606 14872 34612 14884
rect 34563 14844 34612 14872
rect 34563 14841 34575 14844
rect 34517 14835 34575 14841
rect 34606 14832 34612 14844
rect 34664 14832 34670 14884
rect 41386 14872 41414 14980
rect 42981 14977 42993 15011
rect 43027 14977 43039 15011
rect 42981 14971 43039 14977
rect 43254 14968 43260 15020
rect 43312 15008 43318 15020
rect 43349 15011 43407 15017
rect 43349 15008 43361 15011
rect 43312 14980 43361 15008
rect 43312 14968 43318 14980
rect 43349 14977 43361 14980
rect 43395 14977 43407 15011
rect 43349 14971 43407 14977
rect 44266 14968 44272 15020
rect 44324 14968 44330 15020
rect 42613 14943 42671 14949
rect 42613 14909 42625 14943
rect 42659 14940 42671 14943
rect 42794 14940 42800 14952
rect 42659 14912 42800 14940
rect 42659 14909 42671 14912
rect 42613 14903 42671 14909
rect 42794 14900 42800 14912
rect 42852 14900 42858 14952
rect 43070 14900 43076 14952
rect 43128 14900 43134 14952
rect 43346 14872 43352 14884
rect 41386 14844 43352 14872
rect 43346 14832 43352 14844
rect 43404 14832 43410 14884
rect 36078 14804 36084 14816
rect 31726 14776 36084 14804
rect 36078 14764 36084 14776
rect 36136 14764 36142 14816
rect 36814 14764 36820 14816
rect 36872 14764 36878 14816
rect 1104 14714 44620 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 44620 14714
rect 1104 14640 44620 14662
rect 5166 14560 5172 14612
rect 5224 14560 5230 14612
rect 12710 14560 12716 14612
rect 12768 14560 12774 14612
rect 14185 14603 14243 14609
rect 14185 14569 14197 14603
rect 14231 14600 14243 14603
rect 14550 14600 14556 14612
rect 14231 14572 14556 14600
rect 14231 14569 14243 14572
rect 14185 14563 14243 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 16080 14572 16497 14600
rect 16080 14560 16086 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 16592 14572 17080 14600
rect 5184 14464 5212 14560
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 11977 14535 12035 14541
rect 11977 14532 11989 14535
rect 7984 14504 11989 14532
rect 7984 14492 7990 14504
rect 11977 14501 11989 14504
rect 12023 14501 12035 14535
rect 16592 14532 16620 14572
rect 11977 14495 12035 14501
rect 13188 14504 16620 14532
rect 17052 14532 17080 14572
rect 17126 14560 17132 14612
rect 17184 14600 17190 14612
rect 19150 14600 19156 14612
rect 17184 14572 19156 14600
rect 17184 14560 17190 14572
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20128 14572 25176 14600
rect 20128 14560 20134 14572
rect 22830 14532 22836 14544
rect 17052 14504 22836 14532
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 5184 14436 5365 14464
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11664 14368 11897 14396
rect 11664 14356 11670 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12618 14356 12624 14408
rect 12676 14356 12682 14408
rect 13188 14405 13216 14504
rect 22830 14492 22836 14504
rect 22888 14492 22894 14544
rect 25148 14532 25176 14572
rect 25222 14560 25228 14612
rect 25280 14560 25286 14612
rect 25314 14560 25320 14612
rect 25372 14560 25378 14612
rect 27154 14560 27160 14612
rect 27212 14600 27218 14612
rect 34885 14603 34943 14609
rect 27212 14572 31754 14600
rect 27212 14560 27218 14572
rect 25332 14532 25360 14560
rect 25148 14504 25360 14532
rect 25685 14535 25743 14541
rect 25685 14501 25697 14535
rect 25731 14532 25743 14535
rect 25958 14532 25964 14544
rect 25731 14504 25964 14532
rect 25731 14501 25743 14504
rect 25685 14495 25743 14501
rect 25958 14492 25964 14504
rect 26016 14492 26022 14544
rect 26053 14535 26111 14541
rect 26053 14501 26065 14535
rect 26099 14532 26111 14535
rect 26510 14532 26516 14544
rect 26099 14504 26516 14532
rect 26099 14501 26111 14504
rect 26053 14495 26111 14501
rect 26510 14492 26516 14504
rect 26568 14492 26574 14544
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 14829 14467 14887 14473
rect 14829 14464 14841 14467
rect 13596 14436 14841 14464
rect 13596 14424 13602 14436
rect 14829 14433 14841 14436
rect 14875 14464 14887 14467
rect 16301 14467 16359 14473
rect 14875 14436 16252 14464
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 12728 14368 12909 14396
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 12728 14328 12756 14368
rect 12897 14365 12909 14368
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 15764 14405 15792 14436
rect 16224 14408 16252 14436
rect 16301 14433 16313 14467
rect 16347 14464 16359 14467
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16347 14436 16405 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16393 14433 16405 14436
rect 16439 14433 16451 14467
rect 16393 14427 16451 14433
rect 16482 14424 16488 14476
rect 16540 14424 16546 14476
rect 16577 14472 16635 14473
rect 16577 14467 16804 14472
rect 16577 14433 16589 14467
rect 16623 14464 16804 14467
rect 19334 14464 19340 14476
rect 16623 14444 19340 14464
rect 16623 14433 16635 14444
rect 16776 14436 19340 14444
rect 16577 14427 16635 14433
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 22002 14464 22008 14476
rect 21140 14436 22008 14464
rect 21140 14424 21146 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 27430 14424 27436 14476
rect 27488 14464 27494 14476
rect 27798 14464 27804 14476
rect 27488 14436 27804 14464
rect 27488 14424 27494 14436
rect 27798 14424 27804 14436
rect 27856 14464 27862 14476
rect 30466 14464 30472 14476
rect 27856 14436 30472 14464
rect 27856 14424 27862 14436
rect 30466 14424 30472 14436
rect 30524 14424 30530 14476
rect 31726 14464 31754 14572
rect 34885 14569 34897 14603
rect 34931 14600 34943 14603
rect 35342 14600 35348 14612
rect 34931 14572 35348 14600
rect 34931 14569 34943 14572
rect 34885 14563 34943 14569
rect 35342 14560 35348 14572
rect 35400 14560 35406 14612
rect 39942 14560 39948 14612
rect 40000 14560 40006 14612
rect 43254 14560 43260 14612
rect 43312 14560 43318 14612
rect 35161 14467 35219 14473
rect 35161 14464 35173 14467
rect 31726 14436 35173 14464
rect 35161 14433 35173 14436
rect 35207 14433 35219 14467
rect 36814 14464 36820 14476
rect 35161 14427 35219 14433
rect 35360 14436 35756 14464
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14332 14368 14565 14396
rect 14332 14356 14338 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15838 14356 15844 14408
rect 15896 14356 15902 14408
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15988 14368 16037 14396
rect 15988 14356 15994 14368
rect 16025 14365 16037 14368
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 16114 14356 16120 14408
rect 16172 14356 16178 14408
rect 16206 14356 16212 14408
rect 16264 14356 16270 14408
rect 16500 14396 16528 14424
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16500 14368 16681 14396
rect 16669 14365 16681 14368
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 16816 14368 21128 14396
rect 16816 14356 16822 14368
rect 21100 14340 21128 14368
rect 25406 14356 25412 14408
rect 25464 14356 25470 14408
rect 25501 14399 25559 14405
rect 25501 14365 25513 14399
rect 25547 14365 25559 14399
rect 25501 14359 25559 14365
rect 25777 14399 25835 14405
rect 25777 14365 25789 14399
rect 25823 14396 25835 14399
rect 26234 14396 26240 14408
rect 25823 14368 26240 14396
rect 25823 14365 25835 14368
rect 25777 14359 25835 14365
rect 12584 14300 12756 14328
rect 14645 14331 14703 14337
rect 12584 14288 12590 14300
rect 14645 14297 14657 14331
rect 14691 14328 14703 14331
rect 18874 14328 18880 14340
rect 14691 14300 18880 14328
rect 14691 14297 14703 14300
rect 14645 14291 14703 14297
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 21082 14288 21088 14340
rect 21140 14288 21146 14340
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5776 14232 6009 14260
rect 5776 14220 5782 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 18230 14260 18236 14272
rect 13136 14232 18236 14260
rect 13136 14220 13142 14232
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 25516 14260 25544 14359
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14396 31263 14399
rect 31294 14396 31300 14408
rect 31251 14368 31300 14396
rect 31251 14365 31263 14368
rect 31205 14359 31263 14365
rect 31294 14356 31300 14368
rect 31352 14356 31358 14408
rect 31389 14399 31447 14405
rect 31389 14365 31401 14399
rect 31435 14396 31447 14399
rect 31662 14396 31668 14408
rect 31435 14368 31668 14396
rect 31435 14365 31447 14368
rect 31389 14359 31447 14365
rect 31662 14356 31668 14368
rect 31720 14356 31726 14408
rect 34701 14399 34759 14405
rect 34701 14365 34713 14399
rect 34747 14365 34759 14399
rect 34701 14359 34759 14365
rect 34885 14399 34943 14405
rect 34885 14365 34897 14399
rect 34931 14396 34943 14399
rect 35360 14396 35388 14436
rect 35728 14408 35756 14436
rect 36372 14436 36820 14464
rect 34931 14368 35388 14396
rect 34931 14365 34943 14368
rect 34885 14359 34943 14365
rect 26970 14288 26976 14340
rect 27028 14288 27034 14340
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 27525 14331 27583 14337
rect 27525 14328 27537 14331
rect 27304 14300 27537 14328
rect 27304 14288 27310 14300
rect 27525 14297 27537 14300
rect 27571 14297 27583 14331
rect 34716 14328 34744 14359
rect 35434 14356 35440 14408
rect 35492 14356 35498 14408
rect 35710 14356 35716 14408
rect 35768 14356 35774 14408
rect 35989 14399 36047 14405
rect 35989 14365 36001 14399
rect 36035 14396 36047 14399
rect 36078 14396 36084 14408
rect 36035 14368 36084 14396
rect 36035 14365 36047 14368
rect 35989 14359 36047 14365
rect 36078 14356 36084 14368
rect 36136 14356 36142 14408
rect 36372 14405 36400 14436
rect 36814 14424 36820 14436
rect 36872 14464 36878 14476
rect 37001 14467 37059 14473
rect 37001 14464 37013 14467
rect 36872 14436 37013 14464
rect 36872 14424 36878 14436
rect 37001 14433 37013 14436
rect 37047 14433 37059 14467
rect 39960 14464 39988 14560
rect 43073 14535 43131 14541
rect 43073 14501 43085 14535
rect 43119 14532 43131 14535
rect 43349 14535 43407 14541
rect 43349 14532 43361 14535
rect 43119 14504 43361 14532
rect 43119 14501 43131 14504
rect 43073 14495 43131 14501
rect 43349 14501 43361 14504
rect 43395 14501 43407 14535
rect 43349 14495 43407 14501
rect 41325 14467 41383 14473
rect 41325 14464 41337 14467
rect 39960 14436 41337 14464
rect 37001 14427 37059 14433
rect 41325 14433 41337 14436
rect 41371 14433 41383 14467
rect 41325 14427 41383 14433
rect 43714 14424 43720 14476
rect 43772 14424 43778 14476
rect 36357 14399 36415 14405
rect 36357 14365 36369 14399
rect 36403 14365 36415 14399
rect 36357 14359 36415 14365
rect 36449 14331 36507 14337
rect 36449 14328 36461 14331
rect 34716 14300 36461 14328
rect 27525 14291 27583 14297
rect 36449 14297 36461 14300
rect 36495 14297 36507 14331
rect 36449 14291 36507 14297
rect 41598 14288 41604 14340
rect 41656 14288 41662 14340
rect 42242 14288 42248 14340
rect 42300 14288 42306 14340
rect 18840 14232 25544 14260
rect 18840 14220 18846 14232
rect 31294 14220 31300 14272
rect 31352 14220 31358 14272
rect 1104 14170 44620 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 44620 14170
rect 1104 14096 44620 14118
rect 5534 14056 5540 14068
rect 5368 14028 5540 14056
rect 4614 13812 4620 13864
rect 4672 13812 4678 13864
rect 5368 13861 5396 14028
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 7282 14056 7288 14068
rect 5736 14028 7288 14056
rect 5736 13929 5764 14028
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7340 14028 7849 14056
rect 7340 14016 7346 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12434 14056 12440 14068
rect 12299 14028 12440 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 14516 14028 14565 14056
rect 14516 14016 14522 14028
rect 14553 14025 14565 14028
rect 14599 14025 14611 14059
rect 14553 14019 14611 14025
rect 15558 14059 15616 14065
rect 15558 14025 15570 14059
rect 15604 14056 15616 14059
rect 15838 14056 15844 14068
rect 15604 14028 15844 14056
rect 15604 14025 15616 14028
rect 15558 14019 15616 14025
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16172 14028 16681 14056
rect 16172 14016 16178 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 17218 14056 17224 14068
rect 16669 14019 16727 14025
rect 17052 14028 17224 14056
rect 13078 13988 13084 14000
rect 11992 13960 13084 13988
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13821 5411 13855
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5353 13815 5411 13821
rect 5460 13824 5641 13852
rect 4632 13784 4660 13812
rect 5460 13784 5488 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 7116 13852 7144 13883
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7248 13892 7297 13920
rect 7248 13880 7254 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 11992 13929 12020 13960
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13630 13948 13636 14000
rect 13688 13988 13694 14000
rect 15657 13991 15715 13997
rect 15657 13988 15669 13991
rect 13688 13960 14228 13988
rect 13688 13948 13694 13960
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 12526 13880 12532 13932
rect 12584 13880 12590 13932
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 13538 13920 13544 13932
rect 12676 13892 13544 13920
rect 12676 13880 12682 13892
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14200 13920 14228 13960
rect 15304 13960 15669 13988
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14200 13892 14289 13920
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 7116 13824 9628 13852
rect 5629 13815 5687 13821
rect 7484 13793 7512 13824
rect 4632 13756 5488 13784
rect 7469 13787 7527 13793
rect 7469 13753 7481 13787
rect 7515 13753 7527 13787
rect 7469 13747 7527 13753
rect 9600 13728 9628 13824
rect 12250 13812 12256 13864
rect 12308 13812 12314 13864
rect 14182 13852 14188 13864
rect 12820 13824 14188 13852
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 12820 13784 12848 13824
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14366 13812 14372 13864
rect 14424 13812 14430 13864
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 15304 13852 15332 13960
rect 15657 13957 15669 13960
rect 15703 13988 15715 13991
rect 15930 13988 15936 14000
rect 15703 13960 15936 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 15930 13948 15936 13960
rect 15988 13988 15994 14000
rect 17052 13988 17080 14028
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 18509 14059 18567 14065
rect 18509 14025 18521 14059
rect 18555 14056 18567 14059
rect 18690 14056 18696 14068
rect 18555 14028 18696 14056
rect 18555 14025 18567 14028
rect 18509 14019 18567 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 18782 14016 18788 14068
rect 18840 14016 18846 14068
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 21919 14059 21977 14065
rect 21919 14056 21931 14059
rect 18932 14028 21931 14056
rect 18932 14016 18938 14028
rect 21919 14025 21931 14028
rect 21965 14025 21977 14059
rect 21919 14019 21977 14025
rect 22005 14059 22063 14065
rect 22005 14025 22017 14059
rect 22051 14056 22063 14059
rect 22554 14056 22560 14068
rect 22051 14028 22560 14056
rect 22051 14025 22063 14028
rect 22005 14019 22063 14025
rect 22554 14016 22560 14028
rect 22612 14016 22618 14068
rect 22738 14016 22744 14068
rect 22796 14016 22802 14068
rect 22830 14016 22836 14068
rect 22888 14016 22894 14068
rect 30926 14016 30932 14068
rect 30984 14056 30990 14068
rect 30984 14028 31248 14056
rect 30984 14016 30990 14028
rect 15988 13960 17080 13988
rect 15988 13948 15994 13960
rect 17126 13948 17132 14000
rect 17184 13988 17190 14000
rect 20714 13988 20720 14000
rect 17184 13960 18828 13988
rect 17184 13948 17190 13960
rect 18800 13942 18828 13960
rect 19168 13960 20720 13988
rect 15378 13880 15384 13932
rect 15436 13880 15442 13932
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13889 15531 13923
rect 18046 13920 18052 13932
rect 15473 13883 15531 13889
rect 16868 13892 18052 13920
rect 14608 13824 15332 13852
rect 14608 13812 14614 13824
rect 11664 13756 12848 13784
rect 11664 13744 11670 13756
rect 12894 13744 12900 13796
rect 12952 13784 12958 13796
rect 15488 13784 15516 13883
rect 16868 13861 16896 13892
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 18322 13920 18328 13932
rect 18156 13892 18328 13920
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 12952 13756 15516 13784
rect 12952 13744 12958 13756
rect 4062 13676 4068 13728
rect 4120 13676 4126 13728
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6788 13688 6837 13716
rect 6788 13676 6794 13688
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11204 13688 12081 13716
rect 11204 13676 11210 13688
rect 12069 13685 12081 13688
rect 12115 13685 12127 13719
rect 12069 13679 12127 13685
rect 14458 13676 14464 13728
rect 14516 13716 14522 13728
rect 16868 13716 16896 13815
rect 16942 13812 16948 13864
rect 17000 13812 17006 13864
rect 17034 13812 17040 13864
rect 17092 13812 17098 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17310 13852 17316 13864
rect 17175 13824 17316 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 18156 13784 18184 13892
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18800 13929 19104 13942
rect 19168 13929 19196 13960
rect 20714 13948 20720 13960
rect 20772 13948 20778 14000
rect 21821 13991 21879 13997
rect 21821 13957 21833 13991
rect 21867 13988 21879 13991
rect 22370 13988 22376 14000
rect 21867 13960 22376 13988
rect 21867 13957 21879 13960
rect 21821 13951 21879 13957
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 23201 13991 23259 13997
rect 23201 13957 23213 13991
rect 23247 13988 23259 13991
rect 24670 13988 24676 14000
rect 23247 13960 24676 13988
rect 23247 13957 23259 13960
rect 23201 13951 23259 13957
rect 24670 13948 24676 13960
rect 24728 13948 24734 14000
rect 28077 13991 28135 13997
rect 28077 13957 28089 13991
rect 28123 13988 28135 13991
rect 31110 13988 31116 14000
rect 28123 13960 31116 13988
rect 28123 13957 28135 13960
rect 28077 13951 28135 13957
rect 31110 13948 31116 13960
rect 31168 13948 31174 14000
rect 31220 13988 31248 14028
rect 35434 14016 35440 14068
rect 35492 14056 35498 14068
rect 36265 14059 36323 14065
rect 36265 14056 36277 14059
rect 35492 14028 36277 14056
rect 35492 14016 35498 14028
rect 36265 14025 36277 14028
rect 36311 14025 36323 14059
rect 36265 14019 36323 14025
rect 39942 14016 39948 14068
rect 40000 14016 40006 14068
rect 41598 14016 41604 14068
rect 41656 14056 41662 14068
rect 42429 14059 42487 14065
rect 42429 14056 42441 14059
rect 41656 14028 42441 14056
rect 41656 14016 41662 14028
rect 42429 14025 42441 14028
rect 42475 14025 42487 14059
rect 42429 14019 42487 14025
rect 43346 14016 43352 14068
rect 43404 14016 43410 14068
rect 43530 14016 43536 14068
rect 43588 14016 43594 14068
rect 31481 13991 31539 13997
rect 31481 13988 31493 13991
rect 31220 13960 31493 13988
rect 31481 13957 31493 13960
rect 31527 13988 31539 13991
rect 31570 13988 31576 14000
rect 31527 13960 31576 13988
rect 31527 13957 31539 13960
rect 31481 13951 31539 13957
rect 31570 13948 31576 13960
rect 31628 13948 31634 14000
rect 36417 13991 36475 13997
rect 36417 13988 36429 13991
rect 34808 13960 36429 13988
rect 34808 13932 34836 13960
rect 36417 13957 36429 13960
rect 36463 13957 36475 13991
rect 36417 13951 36475 13957
rect 36633 13991 36691 13997
rect 36633 13957 36645 13991
rect 36679 13957 36691 13991
rect 39960 13988 39988 14016
rect 43364 13988 43392 14016
rect 39960 13960 40448 13988
rect 41998 13960 43392 13988
rect 36633 13951 36691 13957
rect 18800 13923 19119 13929
rect 18800 13914 19073 13923
rect 19061 13889 19073 13914
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 19246 13923 19304 13929
rect 19246 13889 19258 13923
rect 19292 13920 19304 13923
rect 20070 13920 20076 13932
rect 19292 13892 20076 13920
rect 19292 13889 19304 13892
rect 19246 13883 19304 13889
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 18966 13861 18972 13875
rect 18288 13824 18368 13852
rect 18288 13812 18294 13824
rect 17276 13756 18184 13784
rect 17276 13744 17282 13756
rect 14516 13688 16896 13716
rect 14516 13676 14522 13688
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 17862 13716 17868 13728
rect 17092 13688 17868 13716
rect 17092 13676 17098 13688
rect 17862 13676 17868 13688
rect 17920 13716 17926 13728
rect 18049 13719 18107 13725
rect 18049 13716 18061 13719
rect 17920 13688 18061 13716
rect 17920 13676 17926 13688
rect 18049 13685 18061 13688
rect 18095 13685 18107 13719
rect 18340 13716 18368 13824
rect 18965 13823 18972 13861
rect 19024 13823 19030 13875
rect 19168 13852 19196 13883
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 22094 13929 22100 13932
rect 22081 13923 22100 13929
rect 22081 13889 22093 13923
rect 22081 13883 22100 13889
rect 22094 13880 22100 13883
rect 22152 13880 22158 13932
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 22204 13892 22477 13920
rect 22204 13852 22232 13892
rect 22465 13889 22477 13892
rect 22511 13920 22523 13923
rect 23106 13920 23112 13932
rect 22511 13892 23112 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 23293 13923 23351 13929
rect 23293 13889 23305 13923
rect 23339 13920 23351 13923
rect 23937 13923 23995 13929
rect 23339 13892 23520 13920
rect 23339 13889 23351 13892
rect 23293 13883 23351 13889
rect 19076 13824 19196 13852
rect 19306 13824 22232 13852
rect 18965 13821 18977 13823
rect 19011 13821 19023 13823
rect 18965 13815 19023 13821
rect 18874 13744 18880 13796
rect 18932 13784 18938 13796
rect 19076 13784 19104 13824
rect 18932 13756 19104 13784
rect 18932 13744 18938 13756
rect 19306 13716 19334 13824
rect 22278 13812 22284 13864
rect 22336 13812 22342 13864
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13821 22431 13855
rect 22373 13815 22431 13821
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 23308 13852 23336 13883
rect 23492 13864 23520 13892
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 22603 13824 23336 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 22388 13784 22416 13815
rect 23382 13812 23388 13864
rect 23440 13812 23446 13864
rect 23474 13812 23480 13864
rect 23532 13812 23538 13864
rect 22738 13784 22744 13796
rect 22388 13756 22744 13784
rect 22738 13744 22744 13756
rect 22796 13744 22802 13796
rect 22830 13744 22836 13796
rect 22888 13784 22894 13796
rect 23952 13784 23980 13883
rect 29086 13880 29092 13932
rect 29144 13880 29150 13932
rect 29917 13923 29975 13929
rect 29917 13920 29929 13923
rect 29196 13892 29929 13920
rect 22888 13756 23980 13784
rect 29104 13784 29132 13880
rect 29196 13864 29224 13892
rect 29917 13889 29929 13892
rect 29963 13920 29975 13923
rect 30006 13920 30012 13932
rect 29963 13892 30012 13920
rect 29963 13889 29975 13892
rect 29917 13883 29975 13889
rect 30006 13880 30012 13892
rect 30064 13880 30070 13932
rect 30098 13880 30104 13932
rect 30156 13929 30162 13932
rect 30156 13923 30205 13929
rect 30156 13889 30159 13923
rect 30193 13889 30205 13923
rect 30156 13883 30205 13889
rect 30156 13880 30162 13883
rect 30926 13880 30932 13932
rect 30984 13880 30990 13932
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13889 31263 13923
rect 31205 13883 31263 13889
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13889 31447 13923
rect 31389 13883 31447 13889
rect 29178 13812 29184 13864
rect 29236 13812 29242 13864
rect 29825 13855 29883 13861
rect 29825 13821 29837 13855
rect 29871 13852 29883 13855
rect 29871 13824 30236 13852
rect 29871 13821 29883 13824
rect 29825 13815 29883 13821
rect 29730 13784 29736 13796
rect 29104 13756 29736 13784
rect 22888 13744 22894 13756
rect 29730 13744 29736 13756
rect 29788 13784 29794 13796
rect 30055 13787 30113 13793
rect 30055 13784 30067 13787
rect 29788 13756 30067 13784
rect 29788 13744 29794 13756
rect 30055 13753 30067 13756
rect 30101 13753 30113 13787
rect 30208 13784 30236 13824
rect 30282 13812 30288 13864
rect 30340 13812 30346 13864
rect 30650 13812 30656 13864
rect 30708 13812 30714 13864
rect 30742 13812 30748 13864
rect 30800 13812 30806 13864
rect 31018 13812 31024 13864
rect 31076 13852 31082 13864
rect 31220 13852 31248 13883
rect 31076 13824 31248 13852
rect 31404 13852 31432 13883
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 31757 13923 31815 13929
rect 31757 13920 31769 13923
rect 31720 13892 31769 13920
rect 31720 13880 31726 13892
rect 31757 13889 31769 13892
rect 31803 13889 31815 13923
rect 31757 13883 31815 13889
rect 34701 13923 34759 13929
rect 34701 13889 34713 13923
rect 34747 13920 34759 13923
rect 34790 13920 34796 13932
rect 34747 13892 34796 13920
rect 34747 13889 34759 13892
rect 34701 13883 34759 13889
rect 34790 13880 34796 13892
rect 34848 13880 34854 13932
rect 34885 13923 34943 13929
rect 34885 13889 34897 13923
rect 34931 13920 34943 13923
rect 34977 13923 35035 13929
rect 34977 13920 34989 13923
rect 34931 13892 34989 13920
rect 34931 13889 34943 13892
rect 34885 13883 34943 13889
rect 34977 13889 34989 13892
rect 35023 13889 35035 13923
rect 34977 13883 35035 13889
rect 35802 13880 35808 13932
rect 35860 13880 35866 13932
rect 31478 13852 31484 13864
rect 31404 13824 31484 13852
rect 31076 13812 31082 13824
rect 31478 13812 31484 13824
rect 31536 13852 31542 13864
rect 31573 13855 31631 13861
rect 31573 13852 31585 13855
rect 31536 13824 31585 13852
rect 31536 13812 31542 13824
rect 31573 13821 31585 13824
rect 31619 13821 31631 13855
rect 31573 13815 31631 13821
rect 35621 13855 35679 13861
rect 35621 13821 35633 13855
rect 35667 13852 35679 13855
rect 36078 13852 36084 13864
rect 35667 13824 36084 13852
rect 35667 13821 35679 13824
rect 35621 13815 35679 13821
rect 36078 13812 36084 13824
rect 36136 13852 36142 13864
rect 36648 13852 36676 13951
rect 39022 13880 39028 13932
rect 39080 13880 39086 13932
rect 40420 13929 40448 13960
rect 40405 13923 40463 13929
rect 40405 13889 40417 13923
rect 40451 13920 40463 13923
rect 40497 13923 40555 13929
rect 40497 13920 40509 13923
rect 40451 13892 40509 13920
rect 40451 13889 40463 13892
rect 40405 13883 40463 13889
rect 40497 13889 40509 13892
rect 40543 13889 40555 13923
rect 40497 13883 40555 13889
rect 43070 13880 43076 13932
rect 43128 13920 43134 13932
rect 43349 13923 43407 13929
rect 43349 13920 43361 13923
rect 43128 13892 43361 13920
rect 43128 13880 43134 13892
rect 43349 13889 43361 13892
rect 43395 13889 43407 13923
rect 43548 13920 43576 14016
rect 44082 13920 44088 13932
rect 43548 13892 44088 13920
rect 43349 13883 43407 13889
rect 36136 13824 36676 13852
rect 36136 13812 36142 13824
rect 40126 13812 40132 13864
rect 40184 13812 40190 13864
rect 40770 13812 40776 13864
rect 40828 13812 40834 13864
rect 42245 13855 42303 13861
rect 42245 13821 42257 13855
rect 42291 13852 42303 13855
rect 42981 13855 43039 13861
rect 42981 13852 42993 13855
rect 42291 13824 42993 13852
rect 42291 13821 42303 13824
rect 42245 13815 42303 13821
rect 42981 13821 42993 13824
rect 43027 13821 43039 13855
rect 43364 13852 43392 13883
rect 44082 13880 44088 13892
rect 44140 13920 44146 13932
rect 44177 13923 44235 13929
rect 44177 13920 44189 13923
rect 44140 13892 44189 13920
rect 44140 13880 44146 13892
rect 44177 13889 44189 13892
rect 44223 13889 44235 13923
rect 44177 13883 44235 13889
rect 43364 13824 44036 13852
rect 42981 13815 43039 13821
rect 30466 13784 30472 13796
rect 30208 13756 30472 13784
rect 30055 13747 30113 13753
rect 30466 13744 30472 13756
rect 30524 13784 30530 13796
rect 30926 13784 30932 13796
rect 30524 13756 30932 13784
rect 30524 13744 30530 13756
rect 30926 13744 30932 13756
rect 30984 13744 30990 13796
rect 32950 13784 32956 13796
rect 31220 13756 32956 13784
rect 18340 13688 19334 13716
rect 18049 13679 18107 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22462 13716 22468 13728
rect 22152 13688 22468 13716
rect 22152 13676 22158 13688
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 22554 13676 22560 13728
rect 22612 13716 22618 13728
rect 23382 13716 23388 13728
rect 22612 13688 23388 13716
rect 22612 13676 22618 13688
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 23753 13719 23811 13725
rect 23753 13685 23765 13719
rect 23799 13716 23811 13719
rect 23842 13716 23848 13728
rect 23799 13688 23848 13716
rect 23799 13685 23811 13688
rect 23753 13679 23811 13685
rect 23842 13676 23848 13688
rect 23900 13716 23906 13728
rect 24762 13716 24768 13728
rect 23900 13688 24768 13716
rect 23900 13676 23906 13688
rect 24762 13676 24768 13688
rect 24820 13676 24826 13728
rect 26878 13676 26884 13728
rect 26936 13716 26942 13728
rect 31220 13716 31248 13756
rect 32950 13744 32956 13756
rect 33008 13744 33014 13796
rect 44008 13793 44036 13824
rect 43993 13787 44051 13793
rect 43993 13753 44005 13787
rect 44039 13753 44051 13787
rect 43993 13747 44051 13753
rect 26936 13688 31248 13716
rect 26936 13676 26942 13688
rect 31386 13676 31392 13728
rect 31444 13716 31450 13728
rect 31481 13719 31539 13725
rect 31481 13716 31493 13719
rect 31444 13688 31493 13716
rect 31444 13676 31450 13688
rect 31481 13685 31493 13688
rect 31527 13685 31539 13719
rect 31481 13679 31539 13685
rect 31941 13719 31999 13725
rect 31941 13685 31953 13719
rect 31987 13716 31999 13719
rect 32674 13716 32680 13728
rect 31987 13688 32680 13716
rect 31987 13685 31999 13688
rect 31941 13679 31999 13685
rect 32674 13676 32680 13688
rect 32732 13676 32738 13728
rect 34698 13676 34704 13728
rect 34756 13676 34762 13728
rect 35894 13676 35900 13728
rect 35952 13676 35958 13728
rect 36449 13719 36507 13725
rect 36449 13685 36461 13719
rect 36495 13716 36507 13719
rect 36814 13716 36820 13728
rect 36495 13688 36820 13716
rect 36495 13685 36507 13688
rect 36449 13679 36507 13685
rect 36814 13676 36820 13688
rect 36872 13676 36878 13728
rect 38657 13719 38715 13725
rect 38657 13685 38669 13719
rect 38703 13716 38715 13719
rect 39574 13716 39580 13728
rect 38703 13688 39580 13716
rect 38703 13685 38715 13688
rect 38657 13679 38715 13685
rect 39574 13676 39580 13688
rect 39632 13676 39638 13728
rect 43254 13676 43260 13728
rect 43312 13676 43318 13728
rect 1104 13626 44620 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 44620 13626
rect 1104 13552 44620 13574
rect 7423 13515 7481 13521
rect 7423 13481 7435 13515
rect 7469 13512 7481 13515
rect 7650 13512 7656 13524
rect 7469 13484 7656 13512
rect 7469 13481 7481 13484
rect 7423 13475 7481 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11974 13512 11980 13524
rect 11655 13484 11980 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12308 13484 13584 13512
rect 12308 13472 12314 13484
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 13556 13444 13584 13484
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13688 13484 13737 13512
rect 13688 13472 13694 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 14277 13515 14335 13521
rect 14277 13481 14289 13515
rect 14323 13512 14335 13515
rect 14366 13512 14372 13524
rect 14323 13484 14372 13512
rect 14323 13481 14335 13484
rect 14277 13475 14335 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 17034 13512 17040 13524
rect 14660 13484 17040 13512
rect 14550 13444 14556 13456
rect 10376 13416 13400 13444
rect 13556 13416 14556 13444
rect 10376 13404 10382 13416
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13376 3847 13379
rect 5629 13379 5687 13385
rect 5629 13376 5641 13379
rect 3835 13348 5641 13376
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 5629 13345 5641 13348
rect 5675 13376 5687 13379
rect 5810 13376 5816 13388
rect 5675 13348 5816 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 5920 13348 6776 13376
rect 5920 13320 5948 13348
rect 5902 13308 5908 13320
rect 5198 13280 5908 13308
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6748 13252 6776 13348
rect 7926 13336 7932 13388
rect 7984 13336 7990 13388
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 8036 13348 10885 13376
rect 4062 13200 4068 13252
rect 4120 13200 4126 13252
rect 6730 13200 6736 13252
rect 6788 13200 6794 13252
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6914 13172 6920 13184
rect 5583 13144 6920 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 8036 13181 8064 13348
rect 10873 13345 10885 13348
rect 10919 13376 10931 13379
rect 11238 13376 11244 13388
rect 10919 13348 11244 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 11238 13336 11244 13348
rect 11296 13336 11302 13388
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8496 13280 8769 13308
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 7248 13144 8033 13172
rect 7248 13132 7254 13144
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8110 13132 8116 13184
rect 8168 13132 8174 13184
rect 8496 13181 8524 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10152 13184 10180 13271
rect 11422 13268 11428 13320
rect 11480 13268 11486 13320
rect 11532 13308 11560 13339
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 13372 13376 13400 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 14660 13376 14688 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17126 13472 17132 13524
rect 17184 13472 17190 13524
rect 17218 13472 17224 13524
rect 17276 13512 17282 13524
rect 17957 13515 18015 13521
rect 17276 13484 17816 13512
rect 17276 13472 17282 13484
rect 17310 13444 17316 13456
rect 13372 13348 14688 13376
rect 12066 13308 12072 13320
rect 11532 13280 12072 13308
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 13372 13317 13400 13348
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14090 13308 14096 13320
rect 13587 13280 14096 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 14660 13317 14688 13348
rect 15028 13416 17316 13444
rect 15028 13320 15056 13416
rect 17310 13404 17316 13416
rect 17368 13444 17374 13456
rect 17368 13416 17540 13444
rect 17368 13404 17374 13416
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 15160 13348 16773 13376
rect 15160 13336 15166 13348
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 16942 13336 16948 13388
rect 17000 13336 17006 13388
rect 17512 13385 17540 13416
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 10336 13212 10609 13240
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 10336 13181 10364 13212
rect 10597 13209 10609 13212
rect 10643 13240 10655 13243
rect 11330 13240 11336 13252
rect 10643 13212 11336 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 14550 13200 14556 13252
rect 14608 13200 14614 13252
rect 10321 13175 10379 13181
rect 10321 13141 10333 13175
rect 10367 13141 10379 13175
rect 10321 13135 10379 13141
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 12250 13172 12256 13184
rect 11296 13144 12256 13172
rect 11296 13132 11302 13144
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 14936 13172 14964 13271
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 16868 13240 16896 13271
rect 16632 13212 16896 13240
rect 17236 13240 17264 13271
rect 17402 13268 17408 13320
rect 17460 13268 17466 13320
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 17788 13317 17816 13484
rect 17957 13481 17969 13515
rect 18003 13512 18015 13515
rect 22278 13512 22284 13524
rect 18003 13484 22284 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23566 13512 23572 13524
rect 23523 13484 23572 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 25041 13515 25099 13521
rect 25041 13481 25053 13515
rect 25087 13512 25099 13515
rect 25406 13512 25412 13524
rect 25087 13484 25412 13512
rect 25087 13481 25099 13484
rect 25041 13475 25099 13481
rect 25406 13472 25412 13484
rect 25464 13472 25470 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 30742 13512 30748 13524
rect 27028 13484 27568 13512
rect 27028 13472 27034 13484
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 18141 13447 18199 13453
rect 18141 13444 18153 13447
rect 18104 13416 18153 13444
rect 18104 13404 18110 13416
rect 18141 13413 18153 13416
rect 18187 13413 18199 13447
rect 18141 13407 18199 13413
rect 20714 13404 20720 13456
rect 20772 13404 20778 13456
rect 20901 13447 20959 13453
rect 20901 13413 20913 13447
rect 20947 13444 20959 13447
rect 20947 13416 23704 13444
rect 20947 13413 20959 13416
rect 20901 13407 20959 13413
rect 18506 13376 18512 13388
rect 17972 13348 18512 13376
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17972 13240 18000 13348
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 21821 13379 21879 13385
rect 21821 13345 21833 13379
rect 21867 13376 21879 13379
rect 21910 13376 21916 13388
rect 21867 13348 21916 13376
rect 21867 13345 21879 13348
rect 21821 13339 21879 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22554 13336 22560 13388
rect 22612 13336 22618 13388
rect 23566 13376 23572 13388
rect 22664 13348 23572 13376
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13308 18107 13311
rect 18138 13308 18144 13320
rect 18095 13280 18144 13308
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18524 13308 18552 13336
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 18524 13280 20453 13308
rect 18233 13271 18291 13277
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 18248 13240 18276 13271
rect 20898 13268 20904 13320
rect 20956 13268 20962 13320
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13308 21695 13311
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 21683 13280 22477 13308
rect 21683 13277 21695 13280
rect 21637 13271 21695 13277
rect 22465 13277 22477 13280
rect 22511 13308 22523 13311
rect 22664 13308 22692 13348
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 22511 13280 22692 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 22738 13268 22744 13320
rect 22796 13268 22802 13320
rect 23014 13268 23020 13320
rect 23072 13268 23078 13320
rect 23109 13311 23167 13317
rect 23109 13277 23121 13311
rect 23155 13277 23167 13311
rect 23109 13271 23167 13277
rect 17236 13212 18000 13240
rect 18064 13212 18276 13240
rect 16632 13200 16638 13212
rect 18064 13184 18092 13212
rect 19334 13200 19340 13252
rect 19392 13200 19398 13252
rect 21450 13200 21456 13252
rect 21508 13240 21514 13252
rect 21545 13243 21603 13249
rect 21545 13240 21557 13243
rect 21508 13212 21557 13240
rect 21508 13200 21514 13212
rect 21545 13209 21557 13212
rect 21591 13240 21603 13243
rect 22756 13240 22784 13268
rect 23124 13240 23152 13271
rect 23198 13268 23204 13320
rect 23256 13268 23262 13320
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 23382 13308 23388 13320
rect 23339 13280 23388 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23676 13308 23704 13416
rect 24121 13379 24179 13385
rect 24121 13345 24133 13379
rect 24167 13376 24179 13379
rect 25590 13376 25596 13388
rect 24167 13348 25596 13376
rect 24167 13345 24179 13348
rect 24121 13339 24179 13345
rect 25590 13336 25596 13348
rect 25648 13336 25654 13388
rect 27430 13336 27436 13388
rect 27488 13336 27494 13388
rect 27540 13376 27568 13484
rect 30116 13484 30748 13512
rect 30116 13376 30144 13484
rect 30742 13472 30748 13484
rect 30800 13472 30806 13524
rect 31018 13472 31024 13524
rect 31076 13472 31082 13524
rect 31202 13472 31208 13524
rect 31260 13512 31266 13524
rect 31478 13512 31484 13524
rect 31260 13484 31484 13512
rect 31260 13472 31266 13484
rect 31478 13472 31484 13484
rect 31536 13472 31542 13524
rect 32950 13472 32956 13524
rect 33008 13512 33014 13524
rect 34425 13515 34483 13521
rect 33008 13484 34192 13512
rect 33008 13472 33014 13484
rect 30190 13404 30196 13456
rect 30248 13404 30254 13456
rect 27540 13348 28856 13376
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 23676 13280 23765 13308
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 23900 13280 23980 13308
rect 23900 13268 23906 13280
rect 21591 13212 22692 13240
rect 22756 13212 23152 13240
rect 21591 13209 21603 13212
rect 21545 13203 21603 13209
rect 17494 13172 17500 13184
rect 14936 13144 17500 13172
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 18046 13132 18052 13184
rect 18104 13132 18110 13184
rect 19352 13172 19380 13200
rect 21177 13175 21235 13181
rect 21177 13172 21189 13175
rect 19352 13144 21189 13172
rect 21177 13141 21189 13144
rect 21223 13141 21235 13175
rect 21177 13135 21235 13141
rect 22002 13132 22008 13184
rect 22060 13132 22066 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22373 13175 22431 13181
rect 22373 13172 22385 13175
rect 22152 13144 22385 13172
rect 22152 13132 22158 13144
rect 22373 13141 22385 13144
rect 22419 13141 22431 13175
rect 22664 13172 22692 13212
rect 22922 13172 22928 13184
rect 22664 13144 22928 13172
rect 22373 13135 22431 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 23124 13172 23152 13212
rect 23569 13243 23627 13249
rect 23569 13209 23581 13243
rect 23615 13240 23627 13243
rect 23658 13240 23664 13252
rect 23615 13212 23664 13240
rect 23615 13209 23627 13212
rect 23569 13203 23627 13209
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 23952 13240 23980 13280
rect 24210 13268 24216 13320
rect 24268 13268 24274 13320
rect 24397 13311 24455 13317
rect 24397 13277 24409 13311
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 23860 13212 23980 13240
rect 23860 13172 23888 13212
rect 23124 13144 23888 13172
rect 23934 13132 23940 13184
rect 23992 13172 23998 13184
rect 24412 13172 24440 13271
rect 24578 13268 24584 13320
rect 24636 13268 24642 13320
rect 24670 13268 24676 13320
rect 24728 13268 24734 13320
rect 24762 13268 24768 13320
rect 24820 13268 24826 13320
rect 28828 13294 28856 13348
rect 30024 13348 30144 13376
rect 30208 13376 30236 13404
rect 30208 13348 30328 13376
rect 29730 13268 29736 13320
rect 29788 13268 29794 13320
rect 30024 13317 30052 13348
rect 30009 13311 30067 13317
rect 30009 13277 30021 13311
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 30098 13268 30104 13320
rect 30156 13308 30162 13320
rect 30300 13317 30328 13348
rect 32490 13336 32496 13388
rect 32548 13336 32554 13388
rect 30193 13311 30251 13317
rect 30193 13308 30205 13311
rect 30156 13280 30205 13308
rect 30156 13268 30162 13280
rect 30193 13277 30205 13280
rect 30239 13277 30251 13311
rect 30193 13271 30251 13277
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13277 30343 13311
rect 30285 13271 30343 13277
rect 30374 13268 30380 13320
rect 30432 13268 30438 13320
rect 30558 13268 30564 13320
rect 30616 13268 30622 13320
rect 30650 13268 30656 13320
rect 30708 13268 30714 13320
rect 31205 13311 31263 13317
rect 31205 13277 31217 13311
rect 31251 13308 31263 13311
rect 31386 13308 31392 13320
rect 31251 13280 31392 13308
rect 31251 13277 31263 13280
rect 31205 13271 31263 13277
rect 31386 13268 31392 13280
rect 31444 13268 31450 13320
rect 31478 13268 31484 13320
rect 31536 13268 31542 13320
rect 31662 13268 31668 13320
rect 31720 13268 31726 13320
rect 34164 13317 34192 13484
rect 34425 13481 34437 13515
rect 34471 13512 34483 13515
rect 35802 13512 35808 13524
rect 34471 13484 35808 13512
rect 34471 13481 34483 13484
rect 34425 13475 34483 13481
rect 32217 13311 32275 13317
rect 32217 13277 32229 13311
rect 32263 13277 32275 13311
rect 32217 13271 32275 13277
rect 34149 13311 34207 13317
rect 34149 13277 34161 13311
rect 34195 13277 34207 13311
rect 34149 13271 34207 13277
rect 27709 13243 27767 13249
rect 27709 13209 27721 13243
rect 27755 13240 27767 13243
rect 27982 13240 27988 13252
rect 27755 13212 27988 13240
rect 27755 13209 27767 13212
rect 27709 13203 27767 13209
rect 27982 13200 27988 13212
rect 28040 13200 28046 13252
rect 31754 13240 31760 13252
rect 29012 13212 31760 13240
rect 23992 13144 24440 13172
rect 23992 13132 23998 13144
rect 26142 13132 26148 13184
rect 26200 13172 26206 13184
rect 29012 13172 29040 13212
rect 31754 13200 31760 13212
rect 31812 13200 31818 13252
rect 26200 13144 29040 13172
rect 26200 13132 26206 13144
rect 29178 13132 29184 13184
rect 29236 13132 29242 13184
rect 29546 13132 29552 13184
rect 29604 13132 29610 13184
rect 30466 13132 30472 13184
rect 30524 13172 30530 13184
rect 30837 13175 30895 13181
rect 30837 13172 30849 13175
rect 30524 13144 30849 13172
rect 30524 13132 30530 13144
rect 30837 13141 30849 13144
rect 30883 13141 30895 13175
rect 30837 13135 30895 13141
rect 30926 13132 30932 13184
rect 30984 13172 30990 13184
rect 32232 13172 32260 13271
rect 34440 13240 34468 13475
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 37550 13472 37556 13524
rect 37608 13512 37614 13524
rect 39022 13512 39028 13524
rect 37608 13484 39028 13512
rect 37608 13472 37614 13484
rect 39022 13472 39028 13484
rect 39080 13472 39086 13524
rect 39114 13472 39120 13524
rect 39172 13512 39178 13524
rect 40681 13515 40739 13521
rect 40681 13512 40693 13515
rect 39172 13484 40693 13512
rect 39172 13472 39178 13484
rect 40681 13481 40693 13484
rect 40727 13481 40739 13515
rect 40681 13475 40739 13481
rect 40770 13472 40776 13524
rect 40828 13512 40834 13524
rect 40865 13515 40923 13521
rect 40865 13512 40877 13515
rect 40828 13484 40877 13512
rect 40828 13472 40834 13484
rect 40865 13481 40877 13484
rect 40911 13481 40923 13515
rect 40865 13475 40923 13481
rect 44082 13472 44088 13524
rect 44140 13472 44146 13524
rect 38381 13447 38439 13453
rect 38381 13413 38393 13447
rect 38427 13444 38439 13447
rect 38427 13416 41092 13444
rect 38427 13413 38439 13416
rect 38381 13407 38439 13413
rect 34701 13379 34759 13385
rect 34701 13345 34713 13379
rect 34747 13376 34759 13379
rect 36078 13376 36084 13388
rect 34747 13348 36084 13376
rect 34747 13345 34759 13348
rect 34701 13339 34759 13345
rect 36078 13336 36084 13348
rect 36136 13336 36142 13388
rect 36170 13336 36176 13388
rect 36228 13336 36234 13388
rect 36449 13379 36507 13385
rect 36449 13345 36461 13379
rect 36495 13376 36507 13379
rect 38289 13379 38347 13385
rect 38289 13376 38301 13379
rect 36495 13348 38301 13376
rect 36495 13345 36507 13348
rect 36449 13339 36507 13345
rect 38289 13345 38301 13348
rect 38335 13345 38347 13379
rect 38289 13339 38347 13345
rect 38304 13308 38332 13339
rect 38930 13336 38936 13388
rect 38988 13376 38994 13388
rect 39025 13379 39083 13385
rect 39025 13376 39037 13379
rect 38988 13348 39037 13376
rect 38988 13336 38994 13348
rect 39025 13345 39037 13348
rect 39071 13345 39083 13379
rect 39025 13339 39083 13345
rect 39114 13336 39120 13388
rect 39172 13336 39178 13388
rect 39206 13336 39212 13388
rect 39264 13376 39270 13388
rect 39853 13379 39911 13385
rect 39853 13376 39865 13379
rect 39264 13348 39865 13376
rect 39264 13336 39270 13348
rect 39853 13345 39865 13348
rect 39899 13345 39911 13379
rect 39853 13339 39911 13345
rect 40497 13379 40555 13385
rect 40497 13345 40509 13379
rect 40543 13376 40555 13379
rect 40543 13348 40816 13376
rect 40543 13345 40555 13348
rect 40497 13339 40555 13345
rect 38304 13280 38700 13308
rect 36262 13240 36268 13252
rect 33718 13212 34468 13240
rect 35742 13212 36268 13240
rect 30984 13144 32260 13172
rect 30984 13132 30990 13144
rect 33318 13132 33324 13184
rect 33376 13172 33382 13184
rect 33796 13172 33824 13212
rect 36262 13200 36268 13212
rect 36320 13240 36326 13252
rect 36320 13212 36676 13240
rect 36320 13200 36326 13212
rect 33376 13144 33824 13172
rect 33376 13132 33382 13144
rect 33962 13132 33968 13184
rect 34020 13132 34026 13184
rect 34330 13132 34336 13184
rect 34388 13172 34394 13184
rect 36541 13175 36599 13181
rect 36541 13172 36553 13175
rect 34388 13144 36553 13172
rect 34388 13132 34394 13144
rect 36541 13141 36553 13144
rect 36587 13141 36599 13175
rect 36648 13172 36676 13212
rect 37550 13200 37556 13252
rect 37608 13240 37614 13252
rect 38013 13243 38071 13249
rect 37608 13212 37688 13240
rect 37608 13200 37614 13212
rect 37660 13172 37688 13212
rect 38013 13209 38025 13243
rect 38059 13240 38071 13243
rect 38378 13240 38384 13252
rect 38059 13212 38384 13240
rect 38059 13209 38071 13212
rect 38013 13203 38071 13209
rect 38378 13200 38384 13212
rect 38436 13200 38442 13252
rect 38562 13249 38568 13252
rect 38540 13243 38568 13249
rect 38540 13209 38552 13243
rect 38540 13203 38568 13209
rect 38562 13200 38568 13203
rect 38620 13200 38626 13252
rect 38672 13240 38700 13280
rect 39298 13268 39304 13320
rect 39356 13268 39362 13320
rect 39574 13268 39580 13320
rect 39632 13308 39638 13320
rect 40788 13317 40816 13348
rect 41064 13317 41092 13416
rect 42613 13379 42671 13385
rect 42613 13345 42625 13379
rect 42659 13376 42671 13379
rect 43254 13376 43260 13388
rect 42659 13348 43260 13376
rect 42659 13345 42671 13348
rect 42613 13339 42671 13345
rect 43254 13336 43260 13348
rect 43312 13336 43318 13388
rect 40589 13311 40647 13317
rect 40589 13308 40601 13311
rect 39632 13280 40601 13308
rect 39632 13268 39638 13280
rect 40589 13277 40601 13280
rect 40635 13277 40647 13311
rect 40589 13271 40647 13277
rect 40773 13311 40831 13317
rect 40773 13277 40785 13311
rect 40819 13277 40831 13311
rect 40773 13271 40831 13277
rect 41049 13311 41107 13317
rect 41049 13277 41061 13311
rect 41095 13277 41107 13311
rect 42337 13311 42395 13317
rect 42337 13308 42349 13311
rect 41049 13271 41107 13277
rect 41386 13280 42349 13308
rect 38838 13240 38844 13252
rect 38672 13212 38844 13240
rect 38838 13200 38844 13212
rect 38896 13240 38902 13252
rect 39666 13240 39672 13252
rect 38896 13212 39672 13240
rect 38896 13200 38902 13212
rect 39666 13200 39672 13212
rect 39724 13240 39730 13252
rect 41386 13240 41414 13280
rect 42337 13277 42349 13280
rect 42383 13277 42395 13311
rect 42337 13271 42395 13277
rect 39724 13212 41414 13240
rect 39724 13200 39730 13212
rect 43346 13200 43352 13252
rect 43404 13200 43410 13252
rect 36648 13144 37688 13172
rect 36541 13135 36599 13141
rect 38654 13132 38660 13184
rect 38712 13132 38718 13184
rect 38749 13175 38807 13181
rect 38749 13141 38761 13175
rect 38795 13172 38807 13175
rect 39390 13172 39396 13184
rect 38795 13144 39396 13172
rect 38795 13141 38807 13144
rect 38749 13135 38807 13141
rect 39390 13132 39396 13144
rect 39448 13132 39454 13184
rect 39482 13132 39488 13184
rect 39540 13132 39546 13184
rect 1104 13082 44620 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 44620 13082
rect 1104 13008 44620 13030
rect 4019 12971 4077 12977
rect 4019 12937 4031 12971
rect 4065 12968 4077 12971
rect 4614 12968 4620 12980
rect 4065 12940 4620 12968
rect 4065 12937 4077 12940
rect 4019 12931 4077 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6052 12940 6377 12968
rect 6052 12928 6058 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 11422 12968 11428 12980
rect 10551 12940 11428 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11609 12971 11667 12977
rect 11609 12937 11621 12971
rect 11655 12968 11667 12971
rect 12894 12968 12900 12980
rect 11655 12940 12900 12968
rect 11655 12937 11667 12940
rect 11609 12931 11667 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15657 12971 15715 12977
rect 15657 12968 15669 12971
rect 15436 12940 15669 12968
rect 15436 12928 15442 12940
rect 15657 12937 15669 12940
rect 15703 12937 15715 12971
rect 15657 12931 15715 12937
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16942 12968 16948 12980
rect 16255 12940 16948 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20898 12968 20904 12980
rect 20027 12940 20904 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 23014 12968 23020 12980
rect 21008 12940 23020 12968
rect 4706 12860 4712 12912
rect 4764 12860 4770 12912
rect 9582 12900 9588 12912
rect 5828 12872 7972 12900
rect 9338 12872 9588 12900
rect 5828 12844 5856 12872
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5718 12832 5724 12844
rect 5491 12804 5724 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5810 12792 5816 12844
rect 5868 12792 5874 12844
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 7650 12832 7656 12844
rect 7423 12804 7656 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7944 12841 7972 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12900 10195 12903
rect 10226 12900 10232 12912
rect 10183 12872 10232 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10353 12903 10411 12909
rect 10353 12869 10365 12903
rect 10399 12900 10411 12903
rect 10686 12900 10692 12912
rect 10399 12872 10692 12900
rect 10399 12869 10411 12872
rect 10353 12863 10411 12869
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 10796 12872 11284 12900
rect 10796 12841 10824 12872
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 7282 12764 7288 12776
rect 6788 12736 7288 12764
rect 6788 12724 6794 12736
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 8110 12764 8116 12776
rect 7791 12736 8116 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 8570 12764 8576 12776
rect 8343 12736 8576 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9723 12767 9781 12773
rect 9723 12733 9735 12767
rect 9769 12764 9781 12767
rect 10134 12764 10140 12776
rect 9769 12736 10140 12764
rect 9769 12733 9781 12736
rect 9723 12727 9781 12733
rect 10134 12724 10140 12736
rect 10192 12764 10198 12776
rect 11164 12764 11192 12795
rect 11256 12773 11284 12872
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 11940 12872 12020 12900
rect 11940 12860 11946 12872
rect 11992 12841 12020 12872
rect 13538 12860 13544 12912
rect 13596 12900 13602 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 13596 12872 16068 12900
rect 13596 12860 13602 12872
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12832 11667 12835
rect 11977 12835 12035 12841
rect 11655 12804 11928 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 10192 12736 11192 12764
rect 11241 12767 11299 12773
rect 10192 12724 10198 12736
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11514 12764 11520 12776
rect 11287 12736 11520 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11900 12764 11928 12804
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 14734 12792 14740 12844
rect 14792 12792 14798 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15013 12835 15071 12841
rect 14875 12804 14964 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 12710 12764 12716 12776
rect 11900 12736 12716 12764
rect 11701 12727 11759 12733
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10336 12668 10609 12696
rect 10336 12637 10364 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 11716 12696 11744 12727
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 11020 12668 11744 12696
rect 11020 12656 11026 12668
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 13004 12696 13032 12727
rect 14936 12708 14964 12804
rect 15013 12801 15025 12835
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 15028 12764 15056 12795
rect 15378 12792 15384 12844
rect 15436 12792 15442 12844
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 15838 12792 15844 12844
rect 15896 12792 15902 12844
rect 16040 12841 16068 12872
rect 16408 12872 17785 12900
rect 16408 12844 16436 12872
rect 17773 12869 17785 12872
rect 17819 12900 17831 12903
rect 18782 12900 18788 12912
rect 17819 12872 18460 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16500 12804 16957 12832
rect 15488 12764 15516 12792
rect 15028 12736 15516 12764
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 16500 12764 16528 12804
rect 16945 12801 16957 12804
rect 16991 12832 17003 12835
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 16991 12804 17233 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17494 12792 17500 12844
rect 17552 12792 17558 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 15703 12736 16528 12764
rect 16669 12767 16727 12773
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15948 12708 15976 12736
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 17972 12764 18000 12795
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 18104 12804 18153 12832
rect 18104 12792 18110 12804
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18230 12792 18236 12844
rect 18288 12792 18294 12844
rect 18432 12841 18460 12872
rect 18524 12872 18788 12900
rect 18524 12844 18552 12872
rect 18782 12860 18788 12872
rect 18840 12900 18846 12912
rect 19153 12903 19211 12909
rect 18840 12872 19012 12900
rect 18840 12860 18846 12872
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 18506 12792 18512 12844
rect 18564 12792 18570 12844
rect 18984 12841 19012 12872
rect 19153 12869 19165 12903
rect 19199 12900 19211 12903
rect 21008 12900 21036 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 23750 12968 23756 12980
rect 23256 12940 23756 12968
rect 23256 12928 23262 12940
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 23845 12971 23903 12977
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24210 12968 24216 12980
rect 23891 12940 24216 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24210 12928 24216 12940
rect 24268 12968 24274 12980
rect 24397 12971 24455 12977
rect 24397 12968 24409 12971
rect 24268 12940 24409 12968
rect 24268 12928 24274 12940
rect 24397 12937 24409 12940
rect 24443 12937 24455 12971
rect 24397 12931 24455 12937
rect 25498 12928 25504 12980
rect 25556 12928 25562 12980
rect 25608 12940 26464 12968
rect 25608 12900 25636 12940
rect 19199 12872 21036 12900
rect 21100 12872 22416 12900
rect 19199 12869 19211 12872
rect 19153 12863 19211 12869
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 18969 12835 19027 12841
rect 18647 12804 18920 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 16715 12736 18000 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 11848 12668 13032 12696
rect 11848 12656 11854 12668
rect 14918 12656 14924 12708
rect 14976 12696 14982 12708
rect 14976 12668 15601 12696
rect 14976 12656 14982 12668
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11296 12600 11897 12628
rect 11296 12588 11302 12600
rect 11885 12597 11897 12600
rect 11931 12597 11943 12631
rect 11885 12591 11943 12597
rect 15010 12588 15016 12640
rect 15068 12588 15074 12640
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 15573 12628 15601 12668
rect 15930 12656 15936 12708
rect 15988 12656 15994 12708
rect 16022 12656 16028 12708
rect 16080 12696 16086 12708
rect 16684 12696 16712 12727
rect 18690 12724 18696 12776
rect 18748 12724 18754 12776
rect 18892 12764 18920 12804
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12832 19671 12835
rect 19978 12832 19984 12844
rect 19659 12804 19984 12832
rect 19659 12801 19671 12804
rect 19613 12795 19671 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21100 12832 21128 12872
rect 20772 12804 21128 12832
rect 20772 12792 20778 12804
rect 21910 12792 21916 12844
rect 21968 12792 21974 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12801 22155 12835
rect 22097 12795 22155 12801
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 18892 12736 19349 12764
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 19518 12724 19524 12776
rect 19576 12724 19582 12776
rect 21928 12764 21956 12792
rect 22112 12764 22140 12795
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22388 12841 22416 12872
rect 23492 12872 25636 12900
rect 25961 12903 26019 12909
rect 22281 12835 22339 12841
rect 22281 12832 22293 12835
rect 22244 12804 22293 12832
rect 22244 12792 22250 12804
rect 22281 12801 22293 12804
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 22465 12835 22523 12841
rect 22465 12801 22477 12835
rect 22511 12832 22523 12835
rect 22649 12835 22707 12841
rect 22511 12804 22600 12832
rect 22511 12801 22523 12804
rect 22465 12795 22523 12801
rect 22572 12764 22600 12804
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 23382 12832 23388 12844
rect 22695 12804 23388 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 23382 12792 23388 12804
rect 23440 12792 23446 12844
rect 22830 12764 22836 12776
rect 21928 12756 22232 12764
rect 21928 12736 22416 12756
rect 22204 12728 22416 12736
rect 16080 12668 16712 12696
rect 17681 12699 17739 12705
rect 16080 12656 16086 12668
rect 17681 12665 17693 12699
rect 17727 12696 17739 12699
rect 18785 12699 18843 12705
rect 18785 12696 18797 12699
rect 17727 12668 18797 12696
rect 17727 12665 17739 12668
rect 17681 12659 17739 12665
rect 18785 12665 18797 12668
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 19150 12656 19156 12708
rect 19208 12696 19214 12708
rect 21821 12699 21879 12705
rect 21821 12696 21833 12699
rect 19208 12668 21833 12696
rect 19208 12656 19214 12668
rect 21821 12665 21833 12668
rect 21867 12665 21879 12699
rect 22388 12696 22416 12728
rect 22572 12736 22836 12764
rect 22572 12696 22600 12736
rect 22830 12724 22836 12736
rect 22888 12724 22894 12776
rect 22922 12724 22928 12776
rect 22980 12764 22986 12776
rect 23492 12773 23520 12872
rect 25961 12869 25973 12903
rect 26007 12900 26019 12903
rect 26234 12900 26240 12912
rect 26007 12872 26240 12900
rect 26007 12869 26019 12872
rect 25961 12863 26019 12869
rect 26234 12860 26240 12872
rect 26292 12860 26298 12912
rect 26436 12900 26464 12940
rect 26970 12928 26976 12980
rect 27028 12928 27034 12980
rect 29546 12928 29552 12980
rect 29604 12928 29610 12980
rect 30650 12928 30656 12980
rect 30708 12968 30714 12980
rect 30837 12971 30895 12977
rect 30837 12968 30849 12971
rect 30708 12940 30849 12968
rect 30708 12928 30714 12940
rect 30837 12937 30849 12940
rect 30883 12937 30895 12971
rect 30837 12931 30895 12937
rect 31294 12928 31300 12980
rect 31352 12928 31358 12980
rect 31570 12928 31576 12980
rect 31628 12928 31634 12980
rect 32585 12971 32643 12977
rect 32585 12937 32597 12971
rect 32631 12968 32643 12971
rect 32766 12968 32772 12980
rect 32631 12940 32772 12968
rect 32631 12937 32643 12940
rect 32585 12931 32643 12937
rect 32766 12928 32772 12940
rect 32824 12928 32830 12980
rect 35069 12971 35127 12977
rect 35069 12937 35081 12971
rect 35115 12968 35127 12971
rect 36170 12968 36176 12980
rect 35115 12940 36176 12968
rect 35115 12937 35127 12940
rect 35069 12931 35127 12937
rect 36170 12928 36176 12940
rect 36228 12928 36234 12980
rect 38838 12968 38844 12980
rect 37292 12940 38844 12968
rect 26436 12872 27384 12900
rect 23555 12835 23613 12841
rect 23555 12801 23567 12835
rect 23601 12832 23613 12835
rect 23601 12804 24256 12832
rect 23601 12801 23613 12804
rect 23555 12795 23613 12801
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 22980 12736 23489 12764
rect 22980 12724 22986 12736
rect 23477 12733 23489 12736
rect 23523 12733 23535 12767
rect 23477 12727 23535 12733
rect 22388 12668 22600 12696
rect 24228 12696 24256 12804
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 25866 12792 25872 12844
rect 25924 12792 25930 12844
rect 26436 12841 26464 12872
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 26602 12792 26608 12844
rect 26660 12792 26666 12844
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 26712 12804 27261 12832
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 26050 12764 26056 12776
rect 24627 12736 26056 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 26050 12724 26056 12736
rect 26108 12764 26114 12776
rect 26712 12764 26740 12804
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27356 12773 27384 12872
rect 27614 12792 27620 12844
rect 27672 12792 27678 12844
rect 28810 12792 28816 12844
rect 28868 12792 28874 12844
rect 29178 12792 29184 12844
rect 29236 12792 29242 12844
rect 29564 12832 29592 12928
rect 31312 12900 31340 12928
rect 31036 12872 31340 12900
rect 29641 12835 29699 12841
rect 29641 12832 29653 12835
rect 29564 12804 29653 12832
rect 29641 12801 29653 12804
rect 29687 12801 29699 12835
rect 29641 12795 29699 12801
rect 29914 12792 29920 12844
rect 29972 12832 29978 12844
rect 30282 12832 30288 12844
rect 29972 12804 30288 12832
rect 29972 12792 29978 12804
rect 30282 12792 30288 12804
rect 30340 12832 30346 12844
rect 31036 12841 31064 12872
rect 30469 12835 30527 12841
rect 30469 12832 30481 12835
rect 30340 12804 30481 12832
rect 30340 12792 30346 12804
rect 30469 12801 30481 12804
rect 30515 12801 30527 12835
rect 30469 12795 30527 12801
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12801 31079 12835
rect 31021 12795 31079 12801
rect 31113 12835 31171 12841
rect 31113 12801 31125 12835
rect 31159 12801 31171 12835
rect 31113 12795 31171 12801
rect 26973 12767 27031 12773
rect 26973 12764 26985 12767
rect 26108 12736 26740 12764
rect 26804 12736 26985 12764
rect 26108 12724 26114 12736
rect 26326 12696 26332 12708
rect 24228 12668 26332 12696
rect 21821 12659 21879 12665
rect 26326 12656 26332 12668
rect 26384 12656 26390 12708
rect 26804 12705 26832 12736
rect 26973 12733 26985 12736
rect 27019 12733 27031 12767
rect 26973 12727 27031 12733
rect 27341 12767 27399 12773
rect 27341 12733 27353 12767
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 28629 12767 28687 12773
rect 28629 12733 28641 12767
rect 28675 12733 28687 12767
rect 31128 12764 31156 12795
rect 31202 12792 31208 12844
rect 31260 12832 31266 12844
rect 31297 12835 31355 12841
rect 31297 12832 31309 12835
rect 31260 12804 31309 12832
rect 31260 12792 31266 12804
rect 31297 12801 31309 12804
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 31389 12835 31447 12841
rect 31389 12801 31401 12835
rect 31435 12832 31447 12835
rect 31588 12832 31616 12928
rect 32674 12860 32680 12912
rect 32732 12860 32738 12912
rect 35345 12903 35403 12909
rect 32876 12872 34376 12900
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31435 12804 31616 12832
rect 31726 12804 32137 12832
rect 31435 12801 31447 12804
rect 31389 12795 31447 12801
rect 31726 12764 31754 12804
rect 32125 12801 32137 12804
rect 32171 12832 32183 12835
rect 32306 12832 32312 12844
rect 32171 12804 32312 12832
rect 32171 12801 32183 12804
rect 32125 12795 32183 12801
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 32398 12792 32404 12844
rect 32456 12792 32462 12844
rect 32876 12832 32904 12872
rect 34348 12844 34376 12872
rect 35345 12869 35357 12903
rect 35391 12900 35403 12903
rect 35894 12900 35900 12912
rect 35391 12872 35900 12900
rect 35391 12869 35403 12872
rect 35345 12863 35403 12869
rect 35894 12860 35900 12872
rect 35952 12860 35958 12912
rect 32784 12804 32904 12832
rect 31128 12736 31754 12764
rect 32217 12767 32275 12773
rect 28629 12727 28687 12733
rect 32217 12733 32229 12767
rect 32263 12764 32275 12767
rect 32784 12764 32812 12804
rect 32950 12792 32956 12844
rect 33008 12792 33014 12844
rect 33226 12832 33232 12844
rect 33060 12804 33232 12832
rect 32263 12736 32812 12764
rect 32263 12733 32275 12736
rect 32217 12727 32275 12733
rect 26789 12699 26847 12705
rect 26789 12665 26801 12699
rect 26835 12665 26847 12699
rect 28644 12696 28672 12727
rect 32858 12724 32864 12776
rect 32916 12724 32922 12776
rect 32398 12696 32404 12708
rect 26789 12659 26847 12665
rect 27080 12668 32404 12696
rect 16114 12628 16120 12640
rect 15573 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16758 12588 16764 12640
rect 16816 12588 16822 12640
rect 17126 12588 17132 12640
rect 17184 12588 17190 12640
rect 17310 12588 17316 12640
rect 17368 12588 17374 12640
rect 17770 12588 17776 12640
rect 17828 12588 17834 12640
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 18322 12628 18328 12640
rect 18196 12600 18328 12628
rect 18196 12588 18202 12600
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22244 12600 22661 12628
rect 22244 12588 22250 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 23937 12631 23995 12637
rect 23937 12628 23949 12631
rect 23532 12600 23949 12628
rect 23532 12588 23538 12600
rect 23937 12597 23949 12600
rect 23983 12597 23995 12631
rect 23937 12591 23995 12597
rect 25590 12588 25596 12640
rect 25648 12628 25654 12640
rect 26421 12631 26479 12637
rect 26421 12628 26433 12631
rect 25648 12600 26433 12628
rect 25648 12588 25654 12600
rect 26421 12597 26433 12600
rect 26467 12597 26479 12631
rect 26421 12591 26479 12597
rect 26510 12588 26516 12640
rect 26568 12628 26574 12640
rect 27080 12628 27108 12668
rect 32398 12656 32404 12668
rect 32456 12696 32462 12708
rect 33060 12696 33088 12804
rect 33226 12792 33232 12804
rect 33284 12792 33290 12844
rect 34330 12792 34336 12844
rect 34388 12792 34394 12844
rect 34698 12792 34704 12844
rect 34756 12832 34762 12844
rect 34977 12835 35035 12841
rect 34977 12832 34989 12835
rect 34756 12804 34989 12832
rect 34756 12792 34762 12804
rect 34977 12801 34989 12804
rect 35023 12801 35035 12835
rect 34977 12795 35035 12801
rect 35161 12835 35219 12841
rect 35161 12801 35173 12835
rect 35207 12832 35219 12835
rect 35710 12832 35716 12844
rect 35207 12804 35716 12832
rect 35207 12801 35219 12804
rect 35161 12795 35219 12801
rect 35710 12792 35716 12804
rect 35768 12832 35774 12844
rect 35805 12835 35863 12841
rect 35805 12832 35817 12835
rect 35768 12804 35817 12832
rect 35768 12792 35774 12804
rect 35805 12801 35817 12804
rect 35851 12801 35863 12835
rect 35986 12835 36044 12841
rect 35986 12832 35998 12835
rect 35805 12795 35863 12801
rect 35912 12804 35998 12832
rect 34790 12724 34796 12776
rect 34848 12764 34854 12776
rect 35912 12764 35940 12804
rect 35986 12801 35998 12804
rect 36032 12801 36044 12835
rect 35986 12795 36044 12801
rect 36078 12792 36084 12844
rect 36136 12792 36142 12844
rect 37292 12841 37320 12940
rect 38838 12928 38844 12940
rect 38896 12928 38902 12980
rect 39025 12971 39083 12977
rect 39025 12937 39037 12971
rect 39071 12968 39083 12971
rect 39206 12968 39212 12980
rect 39071 12940 39212 12968
rect 39071 12937 39083 12940
rect 39025 12931 39083 12937
rect 39132 12909 39160 12940
rect 39206 12928 39212 12940
rect 39264 12928 39270 12980
rect 39298 12928 39304 12980
rect 39356 12928 39362 12980
rect 39482 12928 39488 12980
rect 39540 12928 39546 12980
rect 39761 12971 39819 12977
rect 39761 12937 39773 12971
rect 39807 12968 39819 12971
rect 40126 12968 40132 12980
rect 39807 12940 40132 12968
rect 39807 12937 39819 12940
rect 39761 12931 39819 12937
rect 40126 12928 40132 12940
rect 40184 12928 40190 12980
rect 39117 12903 39175 12909
rect 39117 12869 39129 12903
rect 39163 12869 39175 12903
rect 39316 12900 39344 12928
rect 39316 12872 39436 12900
rect 39117 12863 39175 12869
rect 37277 12835 37335 12841
rect 37277 12801 37289 12835
rect 37323 12801 37335 12835
rect 37277 12795 37335 12801
rect 38562 12792 38568 12844
rect 38620 12792 38626 12844
rect 39022 12832 39028 12844
rect 38686 12804 39028 12832
rect 39022 12792 39028 12804
rect 39080 12792 39086 12844
rect 39301 12835 39359 12841
rect 39301 12801 39313 12835
rect 39347 12801 39359 12835
rect 39301 12795 39359 12801
rect 34848 12736 35940 12764
rect 34848 12724 34854 12736
rect 36262 12724 36268 12776
rect 36320 12724 36326 12776
rect 37550 12724 37556 12776
rect 37608 12724 37614 12776
rect 32456 12668 33088 12696
rect 35621 12699 35679 12705
rect 32456 12656 32462 12668
rect 35621 12665 35633 12699
rect 35667 12696 35679 12699
rect 36280 12696 36308 12724
rect 35667 12668 36308 12696
rect 35667 12665 35679 12668
rect 35621 12659 35679 12665
rect 26568 12600 27108 12628
rect 26568 12588 26574 12600
rect 27154 12588 27160 12640
rect 27212 12628 27218 12640
rect 27433 12631 27491 12637
rect 27433 12628 27445 12631
rect 27212 12600 27445 12628
rect 27212 12588 27218 12600
rect 27433 12597 27445 12600
rect 27479 12597 27491 12631
rect 27433 12591 27491 12597
rect 27522 12588 27528 12640
rect 27580 12588 27586 12640
rect 28994 12588 29000 12640
rect 29052 12588 29058 12640
rect 30285 12631 30343 12637
rect 30285 12597 30297 12631
rect 30331 12628 30343 12631
rect 31478 12628 31484 12640
rect 30331 12600 31484 12628
rect 30331 12597 30343 12600
rect 30285 12591 30343 12597
rect 31478 12588 31484 12600
rect 31536 12588 31542 12640
rect 32122 12588 32128 12640
rect 32180 12588 32186 12640
rect 32490 12588 32496 12640
rect 32548 12628 32554 12640
rect 32677 12631 32735 12637
rect 32677 12628 32689 12631
rect 32548 12600 32689 12628
rect 32548 12588 32554 12600
rect 32677 12597 32689 12600
rect 32723 12597 32735 12631
rect 32677 12591 32735 12597
rect 33137 12631 33195 12637
rect 33137 12597 33149 12631
rect 33183 12628 33195 12631
rect 38580 12628 38608 12792
rect 39316 12696 39344 12795
rect 39408 12764 39436 12872
rect 39500 12832 39528 12928
rect 39577 12835 39635 12841
rect 39577 12832 39589 12835
rect 39500 12804 39589 12832
rect 39577 12801 39589 12804
rect 39623 12801 39635 12835
rect 39577 12795 39635 12801
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 39408 12736 39497 12764
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 39574 12696 39580 12708
rect 39316 12668 39580 12696
rect 39574 12656 39580 12668
rect 39632 12656 39638 12708
rect 33183 12600 38608 12628
rect 33183 12597 33195 12600
rect 33137 12591 33195 12597
rect 1104 12538 44620 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 44620 12538
rect 1104 12464 44620 12486
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10318 12424 10324 12436
rect 10275 12396 10324 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10870 12384 10876 12436
rect 10928 12384 10934 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 11664 12396 11836 12424
rect 11664 12384 11670 12396
rect 10778 12356 10784 12368
rect 9646 12328 10784 12356
rect 9646 12288 9674 12328
rect 10778 12316 10784 12328
rect 10836 12356 10842 12368
rect 11698 12356 11704 12368
rect 10836 12328 11704 12356
rect 10836 12316 10842 12328
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 11808 12297 11836 12396
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 14090 12384 14096 12436
rect 14148 12384 14154 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14884 12396 14933 12424
rect 14884 12384 14890 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 14921 12387 14979 12393
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15436 12396 15761 12424
rect 15436 12384 15442 12396
rect 15749 12393 15761 12396
rect 15795 12424 15807 12427
rect 15838 12424 15844 12436
rect 15795 12396 15844 12424
rect 15795 12393 15807 12396
rect 15749 12387 15807 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 17129 12427 17187 12433
rect 17129 12393 17141 12427
rect 17175 12424 17187 12427
rect 17586 12424 17592 12436
rect 17175 12396 17592 12424
rect 17175 12393 17187 12396
rect 17129 12387 17187 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18690 12384 18696 12436
rect 18748 12424 18754 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18748 12396 19257 12424
rect 18748 12384 18754 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 19981 12427 20039 12433
rect 19981 12424 19993 12427
rect 19576 12396 19993 12424
rect 19576 12384 19582 12396
rect 19981 12393 19993 12396
rect 20027 12393 20039 12427
rect 19981 12387 20039 12393
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 23106 12424 23112 12436
rect 22152 12396 23112 12424
rect 22152 12384 22158 12396
rect 23106 12384 23112 12396
rect 23164 12384 23170 12436
rect 23566 12384 23572 12436
rect 23624 12424 23630 12436
rect 25869 12427 25927 12433
rect 25869 12424 25881 12427
rect 23624 12396 25881 12424
rect 23624 12384 23630 12396
rect 25869 12393 25881 12396
rect 25915 12393 25927 12427
rect 26510 12424 26516 12436
rect 25869 12387 25927 12393
rect 26252 12396 26516 12424
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13814 12356 13820 12368
rect 12768 12328 13820 12356
rect 12768 12316 12774 12328
rect 13814 12316 13820 12328
rect 13872 12356 13878 12368
rect 15102 12356 15108 12368
rect 13872 12328 15108 12356
rect 13872 12316 13878 12328
rect 7208 12260 9674 12288
rect 11793 12291 11851 12297
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7208 12161 7236 12260
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 13998 12288 14004 12300
rect 11793 12251 11851 12257
rect 13004 12260 14004 12288
rect 9784 12192 10548 12220
rect 9784 12164 9812 12192
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6880 12124 7205 12152
rect 6880 12112 6886 12124
rect 7193 12121 7205 12124
rect 7239 12121 7251 12155
rect 7193 12115 7251 12121
rect 9766 12112 9772 12164
rect 9824 12112 9830 12164
rect 9950 12112 9956 12164
rect 10008 12112 10014 12164
rect 10520 12152 10548 12192
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10652 12192 10977 12220
rect 10652 12180 10658 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11296 12192 11345 12220
rect 11296 12180 11302 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12214 11759 12223
rect 13004 12220 13032 12260
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 11900 12214 13032 12220
rect 11747 12192 13032 12214
rect 11747 12189 11928 12192
rect 11701 12186 11928 12189
rect 11701 12183 11759 12186
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 14476 12229 14504 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 15197 12359 15255 12365
rect 15197 12325 15209 12359
rect 15243 12356 15255 12359
rect 15243 12328 18092 12356
rect 15243 12325 15255 12328
rect 15197 12319 15255 12325
rect 15010 12288 15016 12300
rect 14660 12260 15016 12288
rect 14660 12229 14688 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 17770 12288 17776 12300
rect 16868 12260 17776 12288
rect 14277 12223 14335 12229
rect 13136 12214 14228 12220
rect 14277 12214 14289 12223
rect 13136 12192 14289 12214
rect 13136 12180 13142 12192
rect 14200 12189 14289 12192
rect 14323 12189 14335 12223
rect 14200 12186 14335 12189
rect 14277 12183 14335 12186
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 11425 12155 11483 12161
rect 11425 12152 11437 12155
rect 10520 12124 11437 12152
rect 11425 12121 11437 12124
rect 11471 12152 11483 12155
rect 14090 12152 14096 12164
rect 11471 12124 14096 12152
rect 11471 12121 11483 12124
rect 11425 12115 11483 12121
rect 14090 12112 14096 12124
rect 14148 12112 14154 12164
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5684 12056 5733 12084
rect 5684 12044 5690 12056
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 5721 12047 5779 12053
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 10318 12084 10324 12096
rect 7708 12056 10324 12084
rect 7708 12044 7714 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 10468 12056 11621 12084
rect 10468 12044 10474 12056
rect 11609 12053 11621 12056
rect 11655 12084 11667 12087
rect 11698 12084 11704 12096
rect 11655 12056 11704 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 11698 12044 11704 12056
rect 11756 12084 11762 12096
rect 12526 12084 12532 12096
rect 11756 12056 12532 12084
rect 11756 12044 11762 12056
rect 12526 12044 12532 12056
rect 12584 12084 12590 12096
rect 14384 12084 14412 12183
rect 14752 12152 14780 12183
rect 14660 12124 14780 12152
rect 14660 12096 14688 12124
rect 12584 12056 14412 12084
rect 12584 12044 12590 12056
rect 14642 12044 14648 12096
rect 14700 12044 14706 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15120 12084 15148 12183
rect 15286 12180 15292 12232
rect 15344 12180 15350 12232
rect 15378 12180 15384 12232
rect 15436 12180 15442 12232
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15672 12152 15700 12183
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15804 12192 15853 12220
rect 15804 12180 15810 12192
rect 15841 12189 15853 12192
rect 15887 12220 15899 12223
rect 16758 12220 16764 12232
rect 15887 12192 16764 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 16868 12229 16896 12260
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 18064 12164 18092 12328
rect 19426 12316 19432 12368
rect 19484 12356 19490 12368
rect 19794 12356 19800 12368
rect 19484 12328 19800 12356
rect 19484 12316 19490 12328
rect 19794 12316 19800 12328
rect 19852 12316 19858 12368
rect 22189 12359 22247 12365
rect 22189 12325 22201 12359
rect 22235 12356 22247 12359
rect 22462 12356 22468 12368
rect 22235 12328 22468 12356
rect 22235 12325 22247 12328
rect 22189 12319 22247 12325
rect 22462 12316 22468 12328
rect 22520 12356 22526 12368
rect 24397 12359 24455 12365
rect 24397 12356 24409 12359
rect 22520 12328 24409 12356
rect 22520 12316 22526 12328
rect 24397 12325 24409 12328
rect 24443 12325 24455 12359
rect 26252 12356 26280 12396
rect 26510 12384 26516 12396
rect 26568 12384 26574 12436
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 27614 12424 27620 12436
rect 26660 12396 27620 12424
rect 26660 12384 26666 12396
rect 27614 12384 27620 12396
rect 27672 12384 27678 12436
rect 29181 12427 29239 12433
rect 29181 12393 29193 12427
rect 29227 12424 29239 12427
rect 30558 12424 30564 12436
rect 29227 12396 30564 12424
rect 29227 12393 29239 12396
rect 29181 12387 29239 12393
rect 30558 12384 30564 12396
rect 30616 12384 30622 12436
rect 24397 12319 24455 12325
rect 24964 12328 26280 12356
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 18748 12192 19533 12220
rect 18748 12180 18754 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19812 12220 19840 12316
rect 21910 12288 21916 12300
rect 21560 12260 21916 12288
rect 21560 12232 21588 12260
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 23290 12248 23296 12300
rect 23348 12288 23354 12300
rect 24964 12288 24992 12328
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 26384 12328 28212 12356
rect 26384 12316 26390 12328
rect 23348 12260 24992 12288
rect 25041 12291 25099 12297
rect 23348 12248 23354 12260
rect 25041 12257 25053 12291
rect 25087 12288 25099 12291
rect 25130 12288 25136 12300
rect 25087 12260 25136 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 25130 12248 25136 12260
rect 25188 12288 25194 12300
rect 26050 12288 26056 12300
rect 25188 12260 26056 12288
rect 25188 12248 25194 12260
rect 26050 12248 26056 12260
rect 26108 12288 26114 12300
rect 26421 12291 26479 12297
rect 26421 12288 26433 12291
rect 26108 12260 26433 12288
rect 26108 12248 26114 12260
rect 26421 12257 26433 12260
rect 26467 12257 26479 12291
rect 26421 12251 26479 12257
rect 26970 12248 26976 12300
rect 27028 12248 27034 12300
rect 27062 12248 27068 12300
rect 27120 12288 27126 12300
rect 27157 12291 27215 12297
rect 27157 12288 27169 12291
rect 27120 12260 27169 12288
rect 27120 12248 27126 12260
rect 27157 12257 27169 12260
rect 27203 12257 27215 12291
rect 27157 12251 27215 12257
rect 27341 12291 27399 12297
rect 27341 12257 27353 12291
rect 27387 12288 27399 12291
rect 27614 12288 27620 12300
rect 27387 12260 27620 12288
rect 27387 12257 27399 12260
rect 27341 12251 27399 12257
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 27893 12291 27951 12297
rect 27893 12257 27905 12291
rect 27939 12288 27951 12291
rect 27985 12291 28043 12297
rect 27985 12288 27997 12291
rect 27939 12260 27997 12288
rect 27939 12257 27951 12260
rect 27893 12251 27951 12257
rect 27985 12257 27997 12260
rect 28031 12257 28043 12291
rect 28184 12288 28212 12328
rect 29730 12288 29736 12300
rect 28184 12260 28304 12288
rect 27985 12251 28043 12257
rect 19889 12223 19947 12229
rect 19889 12220 19901 12223
rect 19812 12192 19901 12220
rect 19521 12183 19579 12189
rect 19889 12189 19901 12192
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 20070 12180 20076 12232
rect 20128 12180 20134 12232
rect 21542 12180 21548 12232
rect 21600 12180 21606 12232
rect 22002 12180 22008 12232
rect 22060 12180 22066 12232
rect 26329 12223 26387 12229
rect 26329 12189 26341 12223
rect 26375 12220 26387 12223
rect 26988 12220 27016 12248
rect 28276 12229 28304 12260
rect 29196 12260 29736 12288
rect 29196 12229 29224 12260
rect 29730 12248 29736 12260
rect 29788 12248 29794 12300
rect 35437 12291 35495 12297
rect 35437 12288 35449 12291
rect 33980 12260 35449 12288
rect 33980 12232 34008 12260
rect 35437 12257 35449 12260
rect 35483 12288 35495 12291
rect 38194 12288 38200 12300
rect 35483 12260 38200 12288
rect 35483 12257 35495 12260
rect 35437 12251 35495 12257
rect 38194 12248 38200 12260
rect 38252 12248 38258 12300
rect 28169 12223 28227 12229
rect 26375 12192 27016 12220
rect 27264 12192 28028 12220
rect 26375 12189 26387 12192
rect 26329 12183 26387 12189
rect 15672 12124 16252 12152
rect 16224 12096 16252 12124
rect 18046 12112 18052 12164
rect 18104 12152 18110 12164
rect 19150 12152 19156 12164
rect 18104 12124 19156 12152
rect 18104 12112 18110 12124
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19978 12152 19984 12164
rect 19444 12124 19984 12152
rect 16022 12084 16028 12096
rect 14792 12056 16028 12084
rect 14792 12044 14798 12056
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16942 12084 16948 12096
rect 16632 12056 16948 12084
rect 16632 12044 16638 12056
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 19444 12093 19472 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 24302 12112 24308 12164
rect 24360 12152 24366 12164
rect 24360 12124 24900 12152
rect 24360 12112 24366 12124
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12053 19487 12087
rect 19429 12047 19487 12053
rect 19613 12087 19671 12093
rect 19613 12053 19625 12087
rect 19659 12084 19671 12087
rect 20346 12084 20352 12096
rect 19659 12056 20352 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 21821 12087 21879 12093
rect 21821 12084 21833 12087
rect 21784 12056 21833 12084
rect 21784 12044 21790 12056
rect 21821 12053 21833 12056
rect 21867 12053 21879 12087
rect 21821 12047 21879 12053
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 22646 12084 22652 12096
rect 21968 12056 22652 12084
rect 21968 12044 21974 12056
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 24762 12044 24768 12096
rect 24820 12044 24826 12096
rect 24872 12093 24900 12124
rect 26234 12112 26240 12164
rect 26292 12152 26298 12164
rect 27264 12152 27292 12192
rect 26292 12124 27292 12152
rect 26292 12112 26298 12124
rect 27430 12112 27436 12164
rect 27488 12152 27494 12164
rect 27525 12155 27583 12161
rect 27525 12152 27537 12155
rect 27488 12124 27537 12152
rect 27488 12112 27494 12124
rect 27525 12121 27537 12124
rect 27571 12121 27583 12155
rect 27525 12115 27583 12121
rect 27614 12112 27620 12164
rect 27672 12152 27678 12164
rect 28000 12161 28028 12192
rect 28169 12189 28181 12223
rect 28215 12189 28227 12223
rect 28169 12183 28227 12189
rect 28261 12223 28319 12229
rect 28261 12189 28273 12223
rect 28307 12189 28319 12223
rect 28261 12183 28319 12189
rect 29181 12223 29239 12229
rect 29181 12189 29193 12223
rect 29227 12189 29239 12223
rect 29181 12183 29239 12189
rect 27709 12155 27767 12161
rect 27709 12152 27721 12155
rect 27672 12124 27721 12152
rect 27672 12112 27678 12124
rect 27709 12121 27721 12124
rect 27755 12121 27767 12155
rect 27709 12115 27767 12121
rect 27985 12155 28043 12161
rect 27985 12121 27997 12155
rect 28031 12121 28043 12155
rect 27985 12115 28043 12121
rect 28184 12152 28212 12183
rect 29362 12180 29368 12232
rect 29420 12220 29426 12232
rect 30098 12220 30104 12232
rect 29420 12192 30104 12220
rect 29420 12180 29426 12192
rect 30098 12180 30104 12192
rect 30156 12180 30162 12232
rect 30282 12180 30288 12232
rect 30340 12180 30346 12232
rect 31110 12180 31116 12232
rect 31168 12180 31174 12232
rect 33962 12180 33968 12232
rect 34020 12180 34026 12232
rect 34514 12180 34520 12232
rect 34572 12220 34578 12232
rect 34790 12220 34796 12232
rect 34572 12192 34796 12220
rect 34572 12180 34578 12192
rect 34790 12180 34796 12192
rect 34848 12220 34854 12232
rect 34885 12223 34943 12229
rect 34885 12220 34897 12223
rect 34848 12192 34897 12220
rect 34848 12180 34854 12192
rect 34885 12189 34897 12192
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 35066 12180 35072 12232
rect 35124 12180 35130 12232
rect 30300 12152 30328 12180
rect 28184 12124 30328 12152
rect 31128 12152 31156 12180
rect 37921 12155 37979 12161
rect 37921 12152 37933 12155
rect 31128 12124 37933 12152
rect 24857 12087 24915 12093
rect 24857 12053 24869 12087
rect 24903 12084 24915 12087
rect 26697 12087 26755 12093
rect 26697 12084 26709 12087
rect 24903 12056 26709 12084
rect 24903 12053 24915 12056
rect 24857 12047 24915 12053
rect 26697 12053 26709 12056
rect 26743 12053 26755 12087
rect 26697 12047 26755 12053
rect 27065 12087 27123 12093
rect 27065 12053 27077 12087
rect 27111 12084 27123 12087
rect 28184 12084 28212 12124
rect 37921 12121 37933 12124
rect 37967 12152 37979 12155
rect 40494 12152 40500 12164
rect 37967 12124 40500 12152
rect 37967 12121 37979 12124
rect 37921 12115 37979 12121
rect 40494 12112 40500 12124
rect 40552 12152 40558 12164
rect 42518 12152 42524 12164
rect 40552 12124 42524 12152
rect 40552 12112 40558 12124
rect 42518 12112 42524 12124
rect 42576 12112 42582 12164
rect 27111 12056 28212 12084
rect 27111 12053 27123 12056
rect 27065 12047 27123 12053
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 34977 12087 35035 12093
rect 34977 12084 34989 12087
rect 34848 12056 34989 12084
rect 34848 12044 34854 12056
rect 34977 12053 34989 12056
rect 35023 12053 35035 12087
rect 34977 12047 35035 12053
rect 36078 12044 36084 12096
rect 36136 12044 36142 12096
rect 39022 12044 39028 12096
rect 39080 12084 39086 12096
rect 39209 12087 39267 12093
rect 39209 12084 39221 12087
rect 39080 12056 39221 12084
rect 39080 12044 39086 12056
rect 39209 12053 39221 12056
rect 39255 12084 39267 12087
rect 39666 12084 39672 12096
rect 39255 12056 39672 12084
rect 39255 12053 39267 12056
rect 39209 12047 39267 12053
rect 39666 12044 39672 12056
rect 39724 12044 39730 12096
rect 1104 11994 44620 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 44620 11994
rect 1104 11920 44620 11942
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10042 11880 10048 11892
rect 9999 11852 10048 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10686 11840 10692 11892
rect 10744 11840 10750 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 10928 11852 11283 11880
rect 10928 11840 10934 11852
rect 9582 11744 9588 11756
rect 8970 11716 9588 11744
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9674 11704 9680 11756
rect 9732 11704 9738 11756
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10468 11716 10640 11744
rect 10468 11704 10474 11716
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 5684 11648 7573 11676
rect 5684 11636 5690 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7834 11636 7840 11688
rect 7892 11636 7898 11688
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9692 11676 9720 11704
rect 10612 11685 10640 11716
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 11255 11753 11283 11852
rect 11698 11840 11704 11892
rect 11756 11840 11762 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 11974 11880 11980 11892
rect 11931 11852 11980 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12342 11840 12348 11892
rect 12400 11840 12406 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12860 11852 13001 11880
rect 12860 11840 12866 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 12989 11843 13047 11849
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13188 11852 16988 11880
rect 12360 11812 12388 11840
rect 13096 11812 13124 11840
rect 11900 11784 12848 11812
rect 10868 11747 10926 11753
rect 10868 11744 10880 11747
rect 10744 11716 10880 11744
rect 10744 11704 10750 11716
rect 10868 11713 10880 11716
rect 10914 11713 10926 11747
rect 10868 11707 10926 11713
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11240 11747 11298 11753
rect 11240 11713 11252 11747
rect 11286 11713 11298 11747
rect 11240 11707 11298 11713
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11422 11744 11428 11756
rect 11379 11716 11428 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 9355 11648 9720 11676
rect 10597 11679 10655 11685
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10778 11636 10784 11688
rect 10836 11676 10842 11688
rect 10980 11676 11008 11707
rect 10836 11648 11008 11676
rect 10836 11636 10842 11648
rect 10505 11611 10563 11617
rect 10505 11577 10517 11611
rect 10551 11608 10563 11611
rect 11072 11608 11100 11707
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11538 11620 11566 11707
rect 11900 11676 11928 11784
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12618 11744 12624 11756
rect 12391 11716 12624 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 11624 11648 11928 11676
rect 10551 11580 10916 11608
rect 11072 11580 11192 11608
rect 10551 11577 10563 11580
rect 10505 11571 10563 11577
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10778 11540 10784 11552
rect 10459 11512 10784 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10888 11540 10916 11580
rect 11054 11540 11060 11552
rect 10888 11512 11060 11540
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11164 11540 11192 11580
rect 11514 11568 11520 11620
rect 11572 11568 11578 11620
rect 11624 11540 11652 11648
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12728 11676 12756 11704
rect 12299 11648 12756 11676
rect 12820 11676 12848 11784
rect 12912 11784 13124 11812
rect 12912 11756 12940 11784
rect 12894 11704 12900 11756
rect 12952 11704 12958 11756
rect 13188 11753 13216 11852
rect 15856 11784 16896 11812
rect 15856 11753 15884 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 15841 11747 15899 11753
rect 13403 11716 13860 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13188 11676 13216 11707
rect 12820 11648 13216 11676
rect 13449 11679 13507 11685
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 11164 11512 11652 11540
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12710 11540 12716 11552
rect 12584 11512 12716 11540
rect 12584 11500 12590 11512
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13464 11540 13492 11639
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 13832 11676 13860 11716
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16163 11716 16681 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16669 11713 16681 11716
rect 16715 11744 16727 11747
rect 16758 11744 16764 11756
rect 16715 11716 16764 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 14550 11685 14556 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 13832 11648 14381 11676
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 14507 11679 14556 11685
rect 14507 11645 14519 11679
rect 14553 11645 14556 11679
rect 14507 11639 14556 11645
rect 14550 11636 14556 11639
rect 14608 11636 14614 11688
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 14700 11648 15056 11676
rect 14700 11636 14706 11648
rect 14090 11568 14096 11620
rect 14148 11568 14154 11620
rect 15028 11608 15056 11648
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 15562 11676 15568 11688
rect 15252 11648 15568 11676
rect 15252 11636 15258 11648
rect 15562 11636 15568 11648
rect 15620 11676 15626 11688
rect 15856 11676 15884 11707
rect 15620 11648 15884 11676
rect 15620 11636 15626 11648
rect 15930 11636 15936 11688
rect 15988 11636 15994 11688
rect 16040 11676 16068 11707
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16868 11753 16896 11784
rect 16960 11753 16988 11852
rect 17310 11840 17316 11892
rect 17368 11840 17374 11892
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11880 18015 11883
rect 18966 11880 18972 11892
rect 18003 11852 18972 11880
rect 18003 11849 18015 11852
rect 17957 11843 18015 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 22094 11840 22100 11892
rect 22152 11840 22158 11892
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 24489 11883 24547 11889
rect 24489 11849 24501 11883
rect 24535 11880 24547 11883
rect 24670 11880 24676 11892
rect 24535 11852 24676 11880
rect 24535 11849 24547 11852
rect 24489 11843 24547 11849
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 34422 11840 34428 11892
rect 34480 11840 34486 11892
rect 34606 11889 34612 11892
rect 34593 11883 34612 11889
rect 34593 11849 34605 11883
rect 34593 11843 34612 11849
rect 34606 11840 34612 11843
rect 34664 11840 34670 11892
rect 35066 11840 35072 11892
rect 35124 11880 35130 11892
rect 35621 11883 35679 11889
rect 35621 11880 35633 11883
rect 35124 11852 35633 11880
rect 35124 11840 35130 11852
rect 35621 11849 35633 11852
rect 35667 11849 35679 11883
rect 35621 11843 35679 11849
rect 37550 11840 37556 11892
rect 37608 11880 37614 11892
rect 37829 11883 37887 11889
rect 37829 11880 37841 11883
rect 37608 11852 37841 11880
rect 37608 11840 37614 11852
rect 37829 11849 37841 11852
rect 37875 11849 37887 11883
rect 37829 11843 37887 11849
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 16206 11676 16212 11688
rect 16040 11648 16212 11676
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 15654 11608 15660 11620
rect 15028 11580 15660 11608
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 15841 11611 15899 11617
rect 15841 11577 15853 11611
rect 15887 11608 15899 11611
rect 15948 11608 15976 11636
rect 15887 11580 15976 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 17052 11608 17080 11707
rect 18138 11704 18144 11756
rect 18196 11704 18202 11756
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 22480 11753 22508 11840
rect 28810 11812 28816 11824
rect 23584 11784 28816 11812
rect 22373 11747 22431 11753
rect 22373 11713 22385 11747
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 22465 11747 22523 11753
rect 22465 11713 22477 11747
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 22557 11747 22615 11753
rect 22557 11713 22569 11747
rect 22603 11713 22615 11747
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 22557 11707 22615 11713
rect 22664 11716 22753 11744
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 21082 11676 21088 11688
rect 20864 11648 21088 11676
rect 20864 11636 20870 11648
rect 21082 11636 21088 11648
rect 21140 11676 21146 11688
rect 22002 11676 22008 11688
rect 21140 11648 22008 11676
rect 21140 11636 21146 11648
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 22388 11676 22416 11707
rect 22388 11648 22508 11676
rect 16080 11580 17080 11608
rect 16080 11568 16086 11580
rect 22480 11552 22508 11648
rect 22572 11620 22600 11707
rect 22554 11568 22560 11620
rect 22612 11568 22618 11620
rect 22664 11552 22692 11716
rect 22741 11713 22753 11716
rect 22787 11744 22799 11747
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 22787 11716 23213 11744
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23201 11713 23213 11716
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 23216 11676 23244 11707
rect 23290 11704 23296 11756
rect 23348 11744 23354 11756
rect 23584 11753 23612 11784
rect 28810 11772 28816 11784
rect 28868 11772 28874 11824
rect 34793 11815 34851 11821
rect 34793 11781 34805 11815
rect 34839 11781 34851 11815
rect 38654 11812 38660 11824
rect 34793 11775 34851 11781
rect 35544 11784 38660 11812
rect 23385 11747 23443 11753
rect 23385 11744 23397 11747
rect 23348 11716 23397 11744
rect 23348 11704 23354 11716
rect 23385 11713 23397 11716
rect 23431 11713 23443 11747
rect 23385 11707 23443 11713
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 24670 11704 24676 11756
rect 24728 11704 24734 11756
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25590 11744 25596 11756
rect 25004 11716 25596 11744
rect 25004 11704 25010 11716
rect 25590 11704 25596 11716
rect 25648 11704 25654 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 27706 11744 27712 11756
rect 27387 11716 27712 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 27706 11704 27712 11716
rect 27764 11704 27770 11756
rect 23477 11679 23535 11685
rect 23477 11676 23489 11679
rect 23216 11648 23489 11676
rect 23477 11645 23489 11648
rect 23523 11645 23535 11679
rect 23477 11639 23535 11645
rect 27430 11636 27436 11688
rect 27488 11636 27494 11688
rect 27522 11636 27528 11688
rect 27580 11636 27586 11688
rect 28828 11676 28856 11772
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 31662 11744 31668 11756
rect 30800 11716 31668 11744
rect 30800 11704 30806 11716
rect 31662 11704 31668 11716
rect 31720 11744 31726 11756
rect 31757 11747 31815 11753
rect 31757 11744 31769 11747
rect 31720 11716 31769 11744
rect 31720 11704 31726 11716
rect 31757 11713 31769 11716
rect 31803 11713 31815 11747
rect 34808 11744 34836 11775
rect 35342 11744 35348 11756
rect 34808 11716 35348 11744
rect 31757 11707 31815 11713
rect 35342 11704 35348 11716
rect 35400 11744 35406 11756
rect 35437 11747 35495 11753
rect 35437 11744 35449 11747
rect 35400 11716 35449 11744
rect 35400 11704 35406 11716
rect 35437 11713 35449 11716
rect 35483 11713 35495 11747
rect 35437 11707 35495 11713
rect 32858 11676 32864 11688
rect 28828 11648 32864 11676
rect 32858 11636 32864 11648
rect 32916 11676 32922 11688
rect 35544 11676 35572 11784
rect 38654 11772 38660 11784
rect 38712 11772 38718 11824
rect 37921 11747 37979 11753
rect 37921 11713 37933 11747
rect 37967 11744 37979 11747
rect 37967 11716 38424 11744
rect 37967 11713 37979 11716
rect 37921 11707 37979 11713
rect 32916 11648 35572 11676
rect 32916 11636 32922 11648
rect 36170 11636 36176 11688
rect 36228 11636 36234 11688
rect 38396 11685 38424 11716
rect 38470 11704 38476 11756
rect 38528 11744 38534 11756
rect 38841 11747 38899 11753
rect 38841 11744 38853 11747
rect 38528 11716 38853 11744
rect 38528 11704 38534 11716
rect 38841 11713 38853 11716
rect 38887 11713 38899 11747
rect 38841 11707 38899 11713
rect 38381 11679 38439 11685
rect 38381 11645 38393 11679
rect 38427 11645 38439 11679
rect 38381 11639 38439 11645
rect 24762 11568 24768 11620
rect 24820 11608 24826 11620
rect 24857 11611 24915 11617
rect 24857 11608 24869 11611
rect 24820 11580 24869 11608
rect 24820 11568 24826 11580
rect 24857 11577 24869 11580
rect 24903 11608 24915 11611
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 24903 11580 26985 11608
rect 24903 11577 24915 11580
rect 24857 11571 24915 11577
rect 26973 11577 26985 11580
rect 27019 11577 27031 11611
rect 26973 11571 27031 11577
rect 14642 11540 14648 11552
rect 13464 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15289 11543 15347 11549
rect 15289 11509 15301 11543
rect 15335 11540 15347 11543
rect 22002 11540 22008 11552
rect 15335 11512 22008 11540
rect 15335 11509 15347 11512
rect 15289 11503 15347 11509
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 22462 11500 22468 11552
rect 22520 11500 22526 11552
rect 22646 11500 22652 11552
rect 22704 11500 22710 11552
rect 22830 11500 22836 11552
rect 22888 11540 22894 11552
rect 22925 11543 22983 11549
rect 22925 11540 22937 11543
rect 22888 11512 22937 11540
rect 22888 11500 22894 11512
rect 22925 11509 22937 11512
rect 22971 11540 22983 11543
rect 23198 11540 23204 11552
rect 22971 11512 23204 11540
rect 22971 11509 22983 11512
rect 22925 11503 22983 11509
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 27448 11540 27476 11636
rect 31570 11568 31576 11620
rect 31628 11608 31634 11620
rect 32214 11608 32220 11620
rect 31628 11580 32220 11608
rect 31628 11568 31634 11580
rect 32214 11568 32220 11580
rect 32272 11608 32278 11620
rect 32950 11608 32956 11620
rect 32272 11580 32956 11608
rect 32272 11568 32278 11580
rect 32950 11568 32956 11580
rect 33008 11568 33014 11620
rect 36446 11608 36452 11620
rect 34624 11580 36452 11608
rect 29546 11540 29552 11552
rect 27448 11512 29552 11540
rect 29546 11500 29552 11512
rect 29604 11500 29610 11552
rect 31294 11500 31300 11552
rect 31352 11540 31358 11552
rect 34624 11549 34652 11580
rect 36446 11568 36452 11580
rect 36504 11568 36510 11620
rect 31665 11543 31723 11549
rect 31665 11540 31677 11543
rect 31352 11512 31677 11540
rect 31352 11500 31358 11512
rect 31665 11509 31677 11512
rect 31711 11509 31723 11543
rect 31665 11503 31723 11509
rect 34609 11543 34667 11549
rect 34609 11509 34621 11543
rect 34655 11509 34667 11543
rect 34609 11503 34667 11509
rect 34698 11500 34704 11552
rect 34756 11540 34762 11552
rect 34885 11543 34943 11549
rect 34885 11540 34897 11543
rect 34756 11512 34897 11540
rect 34756 11500 34762 11512
rect 34885 11509 34897 11512
rect 34931 11509 34943 11543
rect 34885 11503 34943 11509
rect 38749 11543 38807 11549
rect 38749 11509 38761 11543
rect 38795 11540 38807 11543
rect 38930 11540 38936 11552
rect 38795 11512 38936 11540
rect 38795 11509 38807 11512
rect 38749 11503 38807 11509
rect 38930 11500 38936 11512
rect 38988 11500 38994 11552
rect 1104 11450 44620 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 44620 11450
rect 1104 11376 44620 11398
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7834 11336 7840 11348
rect 7607 11308 7840 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 10781 11339 10839 11345
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 10962 11336 10968 11348
rect 10827 11308 10968 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 10612 11268 10640 11299
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 11839 11308 12020 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 11808 11268 11836 11299
rect 7438 11240 7965 11268
rect 10612 11240 11836 11268
rect 11992 11268 12020 11308
rect 12066 11296 12072 11348
rect 12124 11296 12130 11348
rect 13078 11336 13084 11348
rect 12176 11308 13084 11336
rect 12176 11268 12204 11308
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13170 11296 13176 11348
rect 13228 11296 13234 11348
rect 14108 11308 14504 11336
rect 11992 11240 12204 11268
rect 12437 11271 12495 11277
rect 7438 11200 7466 11240
rect 7392 11172 7466 11200
rect 7653 11203 7711 11209
rect 7392 11144 7420 11172
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7699 11172 7849 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 7937 11144 7965 11240
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7650 11064 7656 11076
rect 7340 11036 7656 11064
rect 7340 11024 7346 11036
rect 7650 11024 7656 11036
rect 7708 11064 7714 11076
rect 7760 11064 7788 11095
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9732 11104 9781 11132
rect 9732 11092 9738 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9769 11095 9827 11101
rect 9876 11104 10425 11132
rect 7708 11036 7788 11064
rect 7708 11024 7714 11036
rect 9876 11008 9904 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10778 11132 10784 11144
rect 10643 11104 10784 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10888 11064 10916 11095
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11164 11141 11192 11240
rect 12437 11237 12449 11271
rect 12483 11268 12495 11271
rect 14108 11268 14136 11308
rect 12483 11240 14136 11268
rect 12483 11237 12495 11240
rect 12437 11231 12495 11237
rect 11330 11200 11336 11212
rect 11256 11172 11336 11200
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 11020 11104 11161 11132
rect 11020 11092 11026 11104
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 11256 11064 11284 11172
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11200 11759 11203
rect 11882 11200 11888 11212
rect 11747 11172 11888 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11992 11172 12265 11200
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11348 11104 11621 11132
rect 11348 11076 11376 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 10428 11036 10916 11064
rect 10980 11036 11284 11064
rect 10428 11008 10456 11036
rect 9858 10956 9864 11008
rect 9916 10956 9922 11008
rect 10410 10956 10416 11008
rect 10468 10956 10474 11008
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 10980 11005 11008 11036
rect 11330 11024 11336 11076
rect 11388 11024 11394 11076
rect 11992 11005 12020 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12207 11104 12296 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12268 11076 12296 11104
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 13188 11132 13216 11163
rect 13262 11160 13268 11212
rect 13320 11160 13326 11212
rect 14476 11200 14504 11308
rect 14550 11296 14556 11348
rect 14608 11296 14614 11348
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14700 11308 14933 11336
rect 14700 11296 14706 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 14921 11299 14979 11305
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 16022 11336 16028 11348
rect 15344 11308 16028 11336
rect 15344 11296 15350 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 18472 11308 18521 11336
rect 18472 11296 18478 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 19978 11336 19984 11348
rect 18739 11308 19984 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 14734 11228 14740 11280
rect 14792 11268 14798 11280
rect 18708 11268 18736 11299
rect 19978 11296 19984 11308
rect 20036 11336 20042 11348
rect 20438 11336 20444 11348
rect 20036 11308 20444 11336
rect 20036 11296 20042 11308
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 21726 11296 21732 11348
rect 21784 11296 21790 11348
rect 22189 11339 22247 11345
rect 22189 11305 22201 11339
rect 22235 11336 22247 11339
rect 22278 11336 22284 11348
rect 22235 11308 22284 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 24670 11296 24676 11348
rect 24728 11336 24734 11348
rect 24949 11339 25007 11345
rect 24949 11336 24961 11339
rect 24728 11308 24961 11336
rect 24728 11296 24734 11308
rect 24949 11305 24961 11308
rect 24995 11305 25007 11339
rect 24949 11299 25007 11305
rect 27246 11296 27252 11348
rect 27304 11336 27310 11348
rect 27985 11339 28043 11345
rect 27985 11336 27997 11339
rect 27304 11308 27997 11336
rect 27304 11296 27310 11308
rect 27985 11305 27997 11308
rect 28031 11305 28043 11339
rect 27985 11299 28043 11305
rect 29546 11296 29552 11348
rect 29604 11296 29610 11348
rect 29914 11296 29920 11348
rect 29972 11296 29978 11348
rect 32030 11296 32036 11348
rect 32088 11336 32094 11348
rect 32582 11336 32588 11348
rect 32088 11308 32588 11336
rect 32088 11296 32094 11308
rect 32582 11296 32588 11308
rect 32640 11296 32646 11348
rect 32858 11296 32864 11348
rect 32916 11296 32922 11348
rect 34698 11296 34704 11348
rect 34756 11296 34762 11348
rect 34790 11296 34796 11348
rect 34848 11336 34854 11348
rect 34958 11339 35016 11345
rect 34958 11336 34970 11339
rect 34848 11308 34970 11336
rect 34848 11296 34854 11308
rect 34958 11305 34970 11308
rect 35004 11305 35016 11339
rect 34958 11299 35016 11305
rect 36446 11296 36452 11348
rect 36504 11296 36510 11348
rect 38930 11296 38936 11348
rect 38988 11296 38994 11348
rect 14792 11240 15240 11268
rect 14792 11228 14798 11240
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 13372 11172 13584 11200
rect 14476 11172 15117 11200
rect 13372 11141 13400 11172
rect 13556 11144 13584 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15212 11200 15240 11240
rect 17972 11240 18736 11268
rect 15271 11203 15329 11209
rect 15271 11200 15283 11203
rect 15212 11172 15283 11200
rect 15105 11163 15163 11169
rect 15271 11169 15283 11172
rect 15317 11169 15329 11203
rect 15271 11163 15329 11169
rect 12584 11104 13216 11132
rect 12584 11092 12590 11104
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 12986 11024 12992 11076
rect 13044 11024 13050 11076
rect 13188 11064 13216 11104
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13446 11092 13452 11144
rect 13504 11092 13510 11144
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 14083 11135 14141 11141
rect 14083 11132 14095 11135
rect 13924 11104 14095 11132
rect 13464 11064 13492 11092
rect 13924 11076 13952 11104
rect 14083 11101 14095 11104
rect 14129 11101 14141 11135
rect 14083 11095 14141 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 13188 11036 13492 11064
rect 13906 11024 13912 11076
rect 13964 11024 13970 11076
rect 14182 11024 14188 11076
rect 14240 11024 14246 11076
rect 14384 11064 14412 11095
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14516 11104 14657 11132
rect 14516 11092 14522 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14384 11036 14749 11064
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 15120 11064 15148 11163
rect 15378 11160 15384 11212
rect 15436 11160 15442 11212
rect 15186 11135 15244 11141
rect 15186 11101 15198 11135
rect 15232 11132 15244 11135
rect 17218 11132 17224 11144
rect 15232 11104 17224 11132
rect 15232 11101 15244 11104
rect 15186 11095 15244 11101
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 17972 11141 18000 11240
rect 18046 11160 18052 11212
rect 18104 11200 18110 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 18104 11172 18613 11200
rect 18104 11160 18110 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 20254 11200 20260 11212
rect 18601 11163 18659 11169
rect 19536 11172 20260 11200
rect 19536 11144 19564 11172
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11101 18015 11135
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17957 11095 18015 11101
rect 18064 11104 18245 11132
rect 16114 11064 16120 11076
rect 15120 11036 16120 11064
rect 14737 11027 14795 11033
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 17678 11064 17684 11076
rect 16816 11036 17684 11064
rect 16816 11024 16822 11036
rect 17678 11024 17684 11036
rect 17736 11064 17742 11076
rect 18064 11064 18092 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 18414 11132 18420 11144
rect 18371 11104 18420 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18748 11104 18889 11132
rect 18748 11092 18754 11104
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19426 11132 19432 11144
rect 19300 11104 19432 11132
rect 19300 11092 19306 11104
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19518 11092 19524 11144
rect 19576 11092 19582 11144
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 20346 11132 20352 11144
rect 19751 11104 20352 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 21266 11132 21272 11144
rect 20548 11104 21272 11132
rect 17736 11036 18092 11064
rect 17736 11024 17742 11036
rect 18138 11024 18144 11076
rect 18196 11024 18202 11076
rect 20548 11064 20576 11104
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11132 21695 11135
rect 21744 11132 21772 11296
rect 22738 11228 22744 11280
rect 22796 11268 22802 11280
rect 23474 11268 23480 11280
rect 22796 11240 23480 11268
rect 22796 11228 22802 11240
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 27614 11228 27620 11280
rect 27672 11268 27678 11280
rect 29932 11268 29960 11296
rect 31757 11271 31815 11277
rect 31757 11268 31769 11271
rect 27672 11240 29960 11268
rect 31128 11240 31769 11268
rect 27672 11228 27678 11240
rect 22925 11203 22983 11209
rect 22925 11200 22937 11203
rect 21836 11172 22937 11200
rect 21836 11141 21864 11172
rect 22925 11169 22937 11172
rect 22971 11169 22983 11203
rect 24946 11200 24952 11212
rect 22925 11163 22983 11169
rect 24872 11172 24952 11200
rect 21683 11104 21772 11132
rect 21821 11135 21879 11141
rect 21683 11101 21695 11104
rect 21637 11095 21695 11101
rect 21821 11101 21833 11135
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 22002 11092 22008 11144
rect 22060 11092 22066 11144
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22281 11135 22339 11141
rect 22281 11132 22293 11135
rect 22152 11104 22293 11132
rect 22152 11092 22158 11104
rect 22281 11101 22293 11104
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22796 11104 22845 11132
rect 22796 11092 22802 11104
rect 22833 11101 22845 11104
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23072 11104 24348 11132
rect 23072 11092 23078 11104
rect 18248 11036 20576 11064
rect 10965 10999 11023 11005
rect 10965 10996 10977 10999
rect 10560 10968 10977 10996
rect 10560 10956 10566 10968
rect 10965 10965 10977 10968
rect 11011 10965 11023 10999
rect 10965 10959 11023 10965
rect 11977 10999 12035 11005
rect 11977 10965 11989 10999
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 18248 10996 18276 11036
rect 20622 11024 20628 11076
rect 20680 11024 20686 11076
rect 20714 11024 20720 11076
rect 20772 11064 20778 11076
rect 21913 11067 21971 11073
rect 21913 11064 21925 11067
rect 20772 11036 21925 11064
rect 20772 11024 20778 11036
rect 21913 11033 21925 11036
rect 21959 11064 21971 11067
rect 22186 11064 22192 11076
rect 21959 11036 22192 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 12124 10968 18276 10996
rect 12124 10956 12130 10968
rect 19058 10956 19064 11008
rect 19116 10956 19122 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19613 10999 19671 11005
rect 19613 10996 19625 10999
rect 19484 10968 19625 10996
rect 19484 10956 19490 10968
rect 19613 10965 19625 10968
rect 19659 10965 19671 10999
rect 20640 10996 20668 11024
rect 24320 11008 24348 11104
rect 24486 11092 24492 11144
rect 24544 11132 24550 11144
rect 24872 11141 24900 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 24857 11135 24915 11141
rect 24857 11132 24869 11135
rect 24544 11104 24869 11132
rect 24544 11092 24550 11104
rect 24857 11101 24869 11104
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11101 25099 11135
rect 25041 11095 25099 11101
rect 25056 11008 25084 11095
rect 27890 11092 27896 11144
rect 27948 11092 27954 11144
rect 28077 11135 28135 11141
rect 28077 11101 28089 11135
rect 28123 11132 28135 11135
rect 28626 11132 28632 11144
rect 28123 11104 28632 11132
rect 28123 11101 28135 11104
rect 28077 11095 28135 11101
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 29730 11092 29736 11144
rect 29788 11092 29794 11144
rect 29822 11092 29828 11144
rect 29880 11092 29886 11144
rect 31128 11141 31156 11240
rect 31757 11237 31769 11240
rect 31803 11268 31815 11271
rect 32674 11268 32680 11280
rect 31803 11240 32680 11268
rect 31803 11237 31815 11240
rect 31757 11231 31815 11237
rect 32674 11228 32680 11240
rect 32732 11228 32738 11280
rect 32769 11271 32827 11277
rect 32769 11237 32781 11271
rect 32815 11268 32827 11271
rect 32876 11268 32904 11296
rect 34716 11268 34744 11296
rect 32815 11240 32904 11268
rect 34348 11240 34744 11268
rect 32815 11237 32827 11240
rect 32769 11231 32827 11237
rect 31294 11160 31300 11212
rect 31352 11160 31358 11212
rect 32582 11160 32588 11212
rect 32640 11160 32646 11212
rect 33137 11203 33195 11209
rect 33137 11169 33149 11203
rect 33183 11200 33195 11203
rect 33226 11200 33232 11212
rect 33183 11172 33232 11200
rect 33183 11169 33195 11172
rect 33137 11163 33195 11169
rect 33226 11160 33232 11172
rect 33284 11160 33290 11212
rect 33778 11160 33784 11212
rect 33836 11200 33842 11212
rect 33965 11203 34023 11209
rect 33965 11200 33977 11203
rect 33836 11172 33977 11200
rect 33836 11160 33842 11172
rect 33965 11169 33977 11172
rect 34011 11169 34023 11203
rect 33965 11163 34023 11169
rect 31113 11135 31171 11141
rect 31113 11101 31125 11135
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 31570 11092 31576 11144
rect 31628 11092 31634 11144
rect 31662 11092 31668 11144
rect 31720 11092 31726 11144
rect 31849 11135 31907 11141
rect 31849 11101 31861 11135
rect 31895 11132 31907 11135
rect 32030 11132 32036 11144
rect 31895 11104 32036 11132
rect 31895 11101 31907 11104
rect 31849 11095 31907 11101
rect 32030 11092 32036 11104
rect 32088 11092 32094 11144
rect 32125 11135 32183 11141
rect 32125 11101 32137 11135
rect 32171 11132 32183 11135
rect 32214 11132 32220 11144
rect 32171 11104 32220 11132
rect 32171 11101 32183 11104
rect 32125 11095 32183 11101
rect 32214 11092 32220 11104
rect 32272 11092 32278 11144
rect 29454 11024 29460 11076
rect 29512 11064 29518 11076
rect 30098 11064 30104 11076
rect 29512 11036 30104 11064
rect 29512 11024 29518 11036
rect 30098 11024 30104 11036
rect 30156 11064 30162 11076
rect 31389 11067 31447 11073
rect 31389 11064 31401 11067
rect 30156 11036 31401 11064
rect 30156 11024 30162 11036
rect 31389 11033 31401 11036
rect 31435 11033 31447 11067
rect 31680 11064 31708 11092
rect 32490 11064 32496 11076
rect 31680 11036 32496 11064
rect 31389 11027 31447 11033
rect 32490 11024 32496 11036
rect 32548 11024 32554 11076
rect 22830 10996 22836 11008
rect 20640 10968 22836 10996
rect 19613 10959 19671 10965
rect 22830 10956 22836 10968
rect 22888 10956 22894 11008
rect 24302 10956 24308 11008
rect 24360 10956 24366 11008
rect 25038 10956 25044 11008
rect 25096 10956 25102 11008
rect 30929 10999 30987 11005
rect 30929 10965 30941 10999
rect 30975 10996 30987 10999
rect 31110 10996 31116 11008
rect 30975 10968 31116 10996
rect 30975 10965 30987 10968
rect 30929 10959 30987 10965
rect 31110 10956 31116 10968
rect 31168 10956 31174 11008
rect 31938 10956 31944 11008
rect 31996 10996 32002 11008
rect 32125 10999 32183 11005
rect 32125 10996 32137 10999
rect 31996 10968 32137 10996
rect 31996 10956 32002 10968
rect 32125 10965 32137 10968
rect 32171 10965 32183 10999
rect 32600 10996 32628 11160
rect 34348 11141 34376 11240
rect 34425 11203 34483 11209
rect 34425 11169 34437 11203
rect 34471 11169 34483 11203
rect 34425 11163 34483 11169
rect 34701 11203 34759 11209
rect 34701 11169 34713 11203
rect 34747 11200 34759 11203
rect 35342 11200 35348 11212
rect 34747 11172 35348 11200
rect 34747 11169 34759 11172
rect 34701 11163 34759 11169
rect 34333 11135 34391 11141
rect 34333 11101 34345 11135
rect 34379 11101 34391 11135
rect 34333 11095 34391 11101
rect 34440 11064 34468 11163
rect 35342 11160 35348 11172
rect 35400 11160 35406 11212
rect 36464 11200 36492 11296
rect 41414 11228 41420 11280
rect 41472 11268 41478 11280
rect 42521 11271 42579 11277
rect 42521 11268 42533 11271
rect 41472 11240 42533 11268
rect 41472 11228 41478 11240
rect 42521 11237 42533 11240
rect 42567 11237 42579 11271
rect 42521 11231 42579 11237
rect 37093 11203 37151 11209
rect 37093 11200 37105 11203
rect 36464 11172 37105 11200
rect 37093 11169 37105 11172
rect 37139 11169 37151 11203
rect 37093 11163 37151 11169
rect 37274 11160 37280 11212
rect 37332 11200 37338 11212
rect 38013 11203 38071 11209
rect 38013 11200 38025 11203
rect 37332 11172 38025 11200
rect 37332 11160 37338 11172
rect 38013 11169 38025 11172
rect 38059 11200 38071 11203
rect 38470 11200 38476 11212
rect 38059 11172 38476 11200
rect 38059 11169 38071 11172
rect 38013 11163 38071 11169
rect 38470 11160 38476 11172
rect 38528 11160 38534 11212
rect 38654 11160 38660 11212
rect 38712 11200 38718 11212
rect 38749 11203 38807 11209
rect 38749 11200 38761 11203
rect 38712 11172 38761 11200
rect 38712 11160 38718 11172
rect 38749 11169 38761 11172
rect 38795 11169 38807 11203
rect 38749 11163 38807 11169
rect 42794 11160 42800 11212
rect 42852 11200 42858 11212
rect 42852 11172 42932 11200
rect 42852 11160 42858 11172
rect 36262 11132 36268 11144
rect 36110 11104 36268 11132
rect 36262 11092 36268 11104
rect 36320 11132 36326 11144
rect 37642 11132 37648 11144
rect 36320 11104 37648 11132
rect 36320 11092 36326 11104
rect 37642 11092 37648 11104
rect 37700 11092 37706 11144
rect 38102 11092 38108 11144
rect 38160 11092 38166 11144
rect 38194 11092 38200 11144
rect 38252 11132 38258 11144
rect 38381 11135 38439 11141
rect 38381 11132 38393 11135
rect 38252 11104 38393 11132
rect 38252 11092 38258 11104
rect 38381 11101 38393 11104
rect 38427 11101 38439 11135
rect 38381 11095 38439 11101
rect 38562 11092 38568 11144
rect 38620 11092 38626 11144
rect 39482 11092 39488 11144
rect 39540 11092 39546 11144
rect 42904 11118 42932 11172
rect 43990 11160 43996 11212
rect 44048 11160 44054 11212
rect 44266 11092 44272 11144
rect 44324 11092 44330 11144
rect 34606 11064 34612 11076
rect 34440 11036 34612 11064
rect 34606 11024 34612 11036
rect 34664 11064 34670 11076
rect 35066 11064 35072 11076
rect 34664 11036 35072 11064
rect 34664 11024 34670 11036
rect 35066 11024 35072 11036
rect 35124 11024 35130 11076
rect 32677 10999 32735 11005
rect 32677 10996 32689 10999
rect 32600 10968 32689 10996
rect 32125 10959 32183 10965
rect 32677 10965 32689 10968
rect 32723 10965 32735 10999
rect 32677 10959 32735 10965
rect 36538 10956 36544 11008
rect 36596 10956 36602 11008
rect 37366 10956 37372 11008
rect 37424 10956 37430 11008
rect 1104 10906 44620 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 44620 10906
rect 1104 10832 44620 10854
rect 6089 10795 6147 10801
rect 6089 10761 6101 10795
rect 6135 10761 6147 10795
rect 6089 10755 6147 10761
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10792 6975 10795
rect 7466 10792 7472 10804
rect 6963 10764 7472 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 6104 10724 6132 10755
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 12066 10792 12072 10804
rect 9646 10764 12072 10792
rect 9646 10724 9674 10764
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 12216 10764 12265 10792
rect 12216 10752 12222 10764
rect 12253 10761 12265 10764
rect 12299 10761 12311 10795
rect 12253 10755 12311 10761
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12986 10792 12992 10804
rect 12759 10764 12992 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15436 10764 15485 10792
rect 15436 10752 15442 10764
rect 15473 10761 15485 10764
rect 15519 10761 15531 10795
rect 15473 10755 15531 10761
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16908 10764 17141 10792
rect 16908 10752 16914 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17494 10792 17500 10804
rect 17276 10764 17500 10792
rect 17276 10752 17282 10764
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 18380 10764 18613 10792
rect 18380 10752 18386 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 18601 10755 18659 10761
rect 19426 10752 19432 10804
rect 19484 10752 19490 10804
rect 20162 10752 20168 10804
rect 20220 10752 20226 10804
rect 21450 10752 21456 10804
rect 21508 10792 21514 10804
rect 21508 10764 22048 10792
rect 21508 10752 21514 10764
rect 6104 10696 9674 10724
rect 11808 10696 12480 10724
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 7098 10656 7104 10668
rect 6595 10628 7104 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 4706 10588 4712 10600
rect 4663 10560 4712 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4356 10452 4384 10551
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 6730 10588 6736 10600
rect 6687 10560 6736 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7524 10560 7941 10588
rect 7524 10548 7530 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 7561 10523 7619 10529
rect 7561 10489 7573 10523
rect 7607 10520 7619 10523
rect 8036 10520 8064 10619
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 11480 10628 11621 10656
rect 11480 10616 11486 10628
rect 11609 10625 11621 10628
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 11808 10588 11836 10696
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12069 10619 12127 10625
rect 12176 10628 12357 10656
rect 9640 10560 11836 10588
rect 9640 10548 9646 10560
rect 7607 10492 8064 10520
rect 7607 10489 7619 10492
rect 7561 10483 7619 10489
rect 10686 10480 10692 10532
rect 10744 10480 10750 10532
rect 10778 10480 10784 10532
rect 10836 10520 10842 10532
rect 11514 10520 11520 10532
rect 10836 10492 11520 10520
rect 10836 10480 10842 10492
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 11790 10480 11796 10532
rect 11848 10520 11854 10532
rect 11900 10520 11928 10619
rect 11992 10532 12020 10619
rect 12084 10532 12112 10619
rect 11848 10492 11928 10520
rect 11848 10480 11854 10492
rect 11974 10480 11980 10532
rect 12032 10480 12038 10532
rect 12066 10480 12072 10532
rect 12124 10480 12130 10532
rect 4614 10452 4620 10464
rect 4356 10424 4620 10452
rect 4614 10412 4620 10424
rect 4672 10452 4678 10464
rect 5626 10452 5632 10464
rect 4672 10424 5632 10452
rect 4672 10412 4678 10424
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 7742 10412 7748 10464
rect 7800 10412 7806 10464
rect 10704 10452 10732 10480
rect 11882 10452 11888 10464
rect 10704 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10452 11946 10464
rect 12176 10452 12204 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12452 10588 12480 10696
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 14182 10724 14188 10736
rect 12860 10696 14188 10724
rect 12860 10684 12866 10696
rect 14182 10684 14188 10696
rect 14240 10724 14246 10736
rect 14734 10724 14740 10736
rect 14240 10696 14740 10724
rect 14240 10684 14246 10696
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 14884 10696 18092 10724
rect 14884 10684 14890 10696
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12618 10656 12624 10668
rect 12575 10628 12624 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13354 10656 13360 10668
rect 13136 10628 13360 10656
rect 13136 10616 13142 10628
rect 13354 10616 13360 10628
rect 13412 10656 13418 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 13412 10628 15393 10656
rect 13412 10616 13418 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 16206 10656 16212 10668
rect 15611 10628 16212 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 12452 10560 14504 10588
rect 14476 10520 14504 10560
rect 14734 10548 14740 10600
rect 14792 10588 14798 10600
rect 15580 10588 15608 10619
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10656 17463 10659
rect 17862 10656 17868 10668
rect 17451 10628 17868 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 18064 10665 18092 10696
rect 18230 10684 18236 10736
rect 18288 10724 18294 10736
rect 19242 10724 19248 10736
rect 18288 10696 19248 10724
rect 18288 10684 18294 10696
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 19444 10724 19472 10752
rect 22020 10736 22048 10764
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22152 10764 22385 10792
rect 22152 10752 22158 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 22563 10795 22621 10801
rect 22563 10761 22575 10795
rect 22609 10792 22621 10795
rect 22922 10792 22928 10804
rect 22609 10764 22928 10792
rect 22609 10761 22621 10764
rect 22563 10755 22621 10761
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 23106 10752 23112 10804
rect 23164 10752 23170 10804
rect 24121 10795 24179 10801
rect 24121 10761 24133 10795
rect 24167 10792 24179 10795
rect 24578 10792 24584 10804
rect 24167 10764 24584 10792
rect 24167 10761 24179 10764
rect 24121 10755 24179 10761
rect 24578 10752 24584 10764
rect 24636 10752 24642 10804
rect 25133 10795 25191 10801
rect 25133 10761 25145 10795
rect 25179 10761 25191 10795
rect 25133 10755 25191 10761
rect 25593 10795 25651 10801
rect 25593 10761 25605 10795
rect 25639 10792 25651 10795
rect 25866 10792 25872 10804
rect 25639 10764 25872 10792
rect 25639 10761 25651 10764
rect 25593 10755 25651 10761
rect 21545 10727 21603 10733
rect 21545 10724 21557 10727
rect 19444 10696 19656 10724
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 19058 10656 19064 10668
rect 18463 10628 19064 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 19628 10665 19656 10696
rect 20824 10696 21557 10724
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 19444 10628 19533 10656
rect 19444 10600 19472 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 20349 10659 20407 10665
rect 20349 10625 20361 10659
rect 20395 10656 20407 10659
rect 20714 10656 20720 10668
rect 20395 10628 20720 10656
rect 20395 10625 20407 10628
rect 20349 10619 20407 10625
rect 14792 10560 15608 10588
rect 14792 10548 14798 10560
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 17494 10588 17500 10600
rect 16172 10560 17500 10588
rect 16172 10548 16178 10560
rect 17494 10548 17500 10560
rect 17552 10588 17558 10600
rect 17681 10591 17739 10597
rect 17681 10588 17693 10591
rect 17552 10560 17693 10588
rect 17552 10548 17558 10560
rect 17681 10557 17693 10560
rect 17727 10557 17739 10591
rect 17681 10551 17739 10557
rect 17770 10548 17776 10600
rect 17828 10548 17834 10600
rect 18322 10548 18328 10600
rect 18380 10548 18386 10600
rect 19426 10548 19432 10600
rect 19484 10548 19490 10600
rect 18340 10520 18368 10548
rect 14476 10492 18368 10520
rect 19245 10523 19303 10529
rect 19245 10489 19257 10523
rect 19291 10520 19303 10523
rect 19904 10520 19932 10619
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20824 10665 20852 10696
rect 21545 10693 21557 10696
rect 21591 10693 21603 10727
rect 21545 10687 21603 10693
rect 22002 10684 22008 10736
rect 22060 10684 22066 10736
rect 23124 10724 23152 10752
rect 25148 10724 25176 10755
rect 25866 10752 25872 10764
rect 25924 10792 25930 10804
rect 26053 10795 26111 10801
rect 26053 10792 26065 10795
rect 25924 10764 26065 10792
rect 25924 10752 25930 10764
rect 26053 10761 26065 10764
rect 26099 10761 26111 10795
rect 26053 10755 26111 10761
rect 26421 10795 26479 10801
rect 26421 10761 26433 10795
rect 26467 10792 26479 10795
rect 27798 10792 27804 10804
rect 26467 10764 27804 10792
rect 26467 10761 26479 10764
rect 26421 10755 26479 10761
rect 27798 10752 27804 10764
rect 27856 10792 27862 10804
rect 27893 10795 27951 10801
rect 27893 10792 27905 10795
rect 27856 10764 27905 10792
rect 27856 10752 27862 10764
rect 27893 10761 27905 10764
rect 27939 10761 27951 10795
rect 29641 10795 29699 10801
rect 27893 10755 27951 10761
rect 28920 10764 29592 10792
rect 22756 10696 25176 10724
rect 26513 10727 26571 10733
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 22094 10656 22100 10668
rect 21683 10628 22100 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 20530 10548 20536 10600
rect 20588 10548 20594 10600
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10588 20683 10591
rect 21266 10588 21272 10600
rect 20671 10560 21272 10588
rect 20671 10557 20683 10560
rect 20625 10551 20683 10557
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 21468 10588 21496 10619
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 21542 10588 21548 10600
rect 21468 10560 21548 10588
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 19291 10492 19932 10520
rect 20073 10523 20131 10529
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 20073 10489 20085 10523
rect 20119 10520 20131 10523
rect 20441 10523 20499 10529
rect 20441 10520 20453 10523
rect 20119 10492 20453 10520
rect 20119 10489 20131 10492
rect 20073 10483 20131 10489
rect 20441 10489 20453 10492
rect 20487 10489 20499 10523
rect 22204 10520 22232 10619
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22336 10628 22477 10656
rect 22336 10616 22342 10628
rect 22465 10625 22477 10628
rect 22511 10656 22523 10659
rect 22511 10628 22600 10656
rect 22511 10625 22523 10628
rect 22465 10619 22523 10625
rect 22462 10520 22468 10532
rect 22204 10492 22468 10520
rect 20441 10483 20499 10489
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 11940 10424 12204 10452
rect 11940 10412 11946 10424
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 17402 10452 17408 10464
rect 14148 10424 17408 10452
rect 14148 10412 14154 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 18104 10424 18153 10452
rect 18104 10412 18110 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19705 10455 19763 10461
rect 19705 10452 19717 10455
rect 19484 10424 19717 10452
rect 19484 10412 19490 10424
rect 19705 10421 19717 10424
rect 19751 10421 19763 10455
rect 22572 10452 22600 10628
rect 22646 10616 22652 10668
rect 22704 10616 22710 10668
rect 22756 10665 22784 10696
rect 26513 10693 26525 10727
rect 26559 10724 26571 10727
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 26559 10696 27445 10724
rect 26559 10693 26571 10696
rect 26513 10687 26571 10693
rect 27433 10693 27445 10696
rect 27479 10724 27491 10727
rect 28077 10727 28135 10733
rect 28077 10724 28089 10727
rect 27479 10696 28089 10724
rect 27479 10693 27491 10696
rect 27433 10687 27491 10693
rect 28077 10693 28089 10696
rect 28123 10693 28135 10727
rect 28813 10727 28871 10733
rect 28813 10724 28825 10727
rect 28077 10687 28135 10693
rect 28368 10696 28825 10724
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 23492 10588 23520 10616
rect 24136 10588 24164 10619
rect 24670 10616 24676 10668
rect 24728 10616 24734 10668
rect 25498 10616 25504 10668
rect 25556 10616 25562 10668
rect 27338 10616 27344 10668
rect 27396 10616 27402 10668
rect 27706 10616 27712 10668
rect 27764 10656 27770 10668
rect 28368 10665 28396 10696
rect 28813 10693 28825 10696
rect 28859 10693 28871 10727
rect 28813 10687 28871 10693
rect 27801 10659 27859 10665
rect 27801 10656 27813 10659
rect 27764 10628 27813 10656
rect 27764 10616 27770 10628
rect 27801 10625 27813 10628
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 28353 10659 28411 10665
rect 28353 10625 28365 10659
rect 28399 10625 28411 10659
rect 28353 10619 28411 10625
rect 28626 10616 28632 10668
rect 28684 10656 28690 10668
rect 28920 10665 28948 10764
rect 29564 10736 29592 10764
rect 29641 10761 29653 10795
rect 29687 10792 29699 10795
rect 29730 10792 29736 10804
rect 29687 10764 29736 10792
rect 29687 10761 29699 10764
rect 29641 10755 29699 10761
rect 29730 10752 29736 10764
rect 29788 10752 29794 10804
rect 30282 10752 30288 10804
rect 30340 10752 30346 10804
rect 30466 10752 30472 10804
rect 30524 10752 30530 10804
rect 31938 10792 31944 10804
rect 30576 10764 31944 10792
rect 28994 10684 29000 10736
rect 29052 10724 29058 10736
rect 29273 10727 29331 10733
rect 29273 10724 29285 10727
rect 29052 10696 29285 10724
rect 29052 10684 29058 10696
rect 28721 10659 28779 10665
rect 28721 10656 28733 10659
rect 28684 10628 28733 10656
rect 28684 10616 28690 10628
rect 28721 10625 28733 10628
rect 28767 10625 28779 10659
rect 28721 10619 28779 10625
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 23492 10560 24164 10588
rect 24765 10591 24823 10597
rect 24765 10557 24777 10591
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 24949 10591 25007 10597
rect 24949 10557 24961 10591
rect 24995 10588 25007 10591
rect 25130 10588 25136 10600
rect 24995 10560 25136 10588
rect 24995 10557 25007 10560
rect 24949 10551 25007 10557
rect 24302 10480 24308 10532
rect 24360 10480 24366 10532
rect 24780 10520 24808 10551
rect 25130 10548 25136 10560
rect 25188 10588 25194 10600
rect 25685 10591 25743 10597
rect 25685 10588 25697 10591
rect 25188 10560 25697 10588
rect 25188 10548 25194 10560
rect 25685 10557 25697 10560
rect 25731 10557 25743 10591
rect 25685 10551 25743 10557
rect 26326 10548 26332 10600
rect 26384 10588 26390 10600
rect 26697 10591 26755 10597
rect 26697 10588 26709 10591
rect 26384 10560 26709 10588
rect 26384 10548 26390 10560
rect 26697 10557 26709 10560
rect 26743 10588 26755 10591
rect 27246 10588 27252 10600
rect 26743 10560 27252 10588
rect 26743 10557 26755 10560
rect 26697 10551 26755 10557
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 27430 10548 27436 10600
rect 27488 10588 27494 10600
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 27488 10560 27537 10588
rect 27488 10548 27494 10560
rect 27525 10557 27537 10560
rect 27571 10557 27583 10591
rect 27525 10551 27583 10557
rect 28077 10591 28135 10597
rect 28077 10557 28089 10591
rect 28123 10588 28135 10591
rect 28534 10588 28540 10600
rect 28123 10560 28540 10588
rect 28123 10557 28135 10560
rect 28077 10551 28135 10557
rect 28534 10548 28540 10560
rect 28592 10588 28598 10600
rect 29089 10591 29147 10597
rect 29089 10588 29101 10591
rect 28592 10560 29101 10588
rect 28592 10548 28598 10560
rect 29089 10557 29101 10560
rect 29135 10557 29147 10591
rect 29089 10551 29147 10557
rect 25038 10520 25044 10532
rect 24780 10492 25044 10520
rect 25038 10480 25044 10492
rect 25096 10520 25102 10532
rect 26973 10523 27031 10529
rect 26973 10520 26985 10523
rect 25096 10492 26985 10520
rect 25096 10480 25102 10492
rect 26973 10489 26985 10492
rect 27019 10489 27031 10523
rect 29196 10520 29224 10696
rect 29273 10693 29285 10696
rect 29319 10693 29331 10727
rect 29273 10687 29331 10693
rect 29454 10684 29460 10736
rect 29512 10684 29518 10736
rect 29546 10684 29552 10736
rect 29604 10724 29610 10736
rect 30484 10724 30512 10752
rect 30576 10733 30604 10764
rect 31938 10752 31944 10764
rect 31996 10792 32002 10804
rect 32214 10792 32220 10804
rect 31996 10764 32220 10792
rect 31996 10752 32002 10764
rect 32214 10752 32220 10764
rect 32272 10752 32278 10804
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 34848 10764 35112 10792
rect 34848 10752 34854 10764
rect 29604 10696 30512 10724
rect 30561 10727 30619 10733
rect 29604 10684 29610 10696
rect 30561 10693 30573 10727
rect 30607 10693 30619 10727
rect 30561 10687 30619 10693
rect 30653 10727 30711 10733
rect 30653 10693 30665 10727
rect 30699 10724 30711 10727
rect 30742 10724 30748 10736
rect 30699 10696 30748 10724
rect 30699 10693 30711 10696
rect 30653 10687 30711 10693
rect 30742 10684 30748 10696
rect 30800 10684 30806 10736
rect 31110 10684 31116 10736
rect 31168 10724 31174 10736
rect 31168 10696 32352 10724
rect 31168 10684 31174 10696
rect 31680 10668 31708 10696
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10656 29883 10659
rect 30374 10656 30380 10668
rect 29871 10628 30380 10656
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 30374 10616 30380 10628
rect 30432 10656 30438 10668
rect 30469 10659 30527 10665
rect 30469 10656 30481 10659
rect 30432 10628 30481 10656
rect 30432 10616 30438 10628
rect 30469 10625 30481 10628
rect 30515 10625 30527 10659
rect 30469 10619 30527 10625
rect 30834 10616 30840 10668
rect 30892 10616 30898 10668
rect 30929 10659 30987 10665
rect 30929 10625 30941 10659
rect 30975 10656 30987 10659
rect 31205 10659 31263 10665
rect 30975 10628 31156 10656
rect 30975 10625 30987 10628
rect 30929 10619 30987 10625
rect 29917 10591 29975 10597
rect 29917 10557 29929 10591
rect 29963 10557 29975 10591
rect 29917 10551 29975 10557
rect 26973 10483 27031 10489
rect 27080 10492 29224 10520
rect 29932 10520 29960 10551
rect 30006 10548 30012 10600
rect 30064 10548 30070 10600
rect 30101 10591 30159 10597
rect 30101 10557 30113 10591
rect 30147 10588 30159 10591
rect 31021 10591 31079 10597
rect 31021 10588 31033 10591
rect 30147 10560 31033 10588
rect 30147 10557 30159 10560
rect 30101 10551 30159 10557
rect 31021 10557 31033 10560
rect 31067 10557 31079 10591
rect 31021 10551 31079 10557
rect 31128 10520 31156 10628
rect 31205 10625 31217 10659
rect 31251 10656 31263 10659
rect 31573 10659 31631 10665
rect 31573 10656 31585 10659
rect 31251 10628 31585 10656
rect 31251 10625 31263 10628
rect 31205 10619 31263 10625
rect 31573 10625 31585 10628
rect 31619 10625 31631 10659
rect 31573 10619 31631 10625
rect 31220 10532 31248 10619
rect 31662 10616 31668 10668
rect 31720 10656 31726 10668
rect 31720 10628 31745 10656
rect 31720 10616 31726 10628
rect 31938 10616 31944 10668
rect 31996 10616 32002 10668
rect 32324 10665 32352 10696
rect 33778 10684 33784 10736
rect 33836 10684 33842 10736
rect 35084 10724 35112 10764
rect 35250 10752 35256 10804
rect 35308 10792 35314 10804
rect 35437 10795 35495 10801
rect 35437 10792 35449 10795
rect 35308 10764 35449 10792
rect 35308 10752 35314 10764
rect 35437 10761 35449 10764
rect 35483 10761 35495 10795
rect 36262 10792 36268 10804
rect 35437 10755 35495 10761
rect 35544 10764 36268 10792
rect 35544 10724 35572 10764
rect 36262 10752 36268 10764
rect 36320 10752 36326 10804
rect 37093 10795 37151 10801
rect 37093 10761 37105 10795
rect 37139 10792 37151 10795
rect 37274 10792 37280 10804
rect 37139 10764 37280 10792
rect 37139 10761 37151 10764
rect 37093 10755 37151 10761
rect 37274 10752 37280 10764
rect 37332 10752 37338 10804
rect 37366 10752 37372 10804
rect 37424 10752 37430 10804
rect 39025 10795 39083 10801
rect 39025 10761 39037 10795
rect 39071 10792 39083 10795
rect 39482 10792 39488 10804
rect 39071 10764 39488 10792
rect 39071 10761 39083 10764
rect 39025 10755 39083 10761
rect 39482 10752 39488 10764
rect 39540 10752 39546 10804
rect 35006 10696 35572 10724
rect 35621 10727 35679 10733
rect 35621 10693 35633 10727
rect 35667 10724 35679 10727
rect 36538 10724 36544 10736
rect 35667 10696 36544 10724
rect 35667 10693 35679 10696
rect 35621 10687 35679 10693
rect 36538 10684 36544 10696
rect 36596 10684 36602 10736
rect 37384 10724 37412 10752
rect 37553 10727 37611 10733
rect 37553 10724 37565 10727
rect 37384 10696 37565 10724
rect 37553 10693 37565 10696
rect 37599 10693 37611 10727
rect 37553 10687 37611 10693
rect 37642 10684 37648 10736
rect 37700 10724 37706 10736
rect 37700 10696 38042 10724
rect 37700 10684 37706 10696
rect 32125 10659 32183 10665
rect 32125 10656 32137 10659
rect 32048 10628 32137 10656
rect 32048 10600 32076 10628
rect 32125 10625 32137 10628
rect 32171 10625 32183 10659
rect 32125 10619 32183 10625
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32490 10616 32496 10668
rect 32548 10616 32554 10668
rect 32677 10659 32735 10665
rect 32677 10625 32689 10659
rect 32723 10656 32735 10659
rect 32950 10656 32956 10668
rect 32723 10628 32956 10656
rect 32723 10625 32735 10628
rect 32677 10619 32735 10625
rect 32950 10616 32956 10628
rect 33008 10616 33014 10668
rect 35066 10616 35072 10668
rect 35124 10656 35130 10668
rect 35345 10659 35403 10665
rect 35345 10656 35357 10659
rect 35124 10628 35357 10656
rect 35124 10616 35130 10628
rect 35345 10625 35357 10628
rect 35391 10656 35403 10659
rect 35526 10656 35532 10668
rect 35391 10628 35532 10656
rect 35391 10625 35403 10628
rect 35345 10619 35403 10625
rect 35526 10616 35532 10628
rect 35584 10616 35590 10668
rect 36078 10616 36084 10668
rect 36136 10656 36142 10668
rect 36817 10659 36875 10665
rect 36817 10656 36829 10659
rect 36136 10628 36829 10656
rect 36136 10616 36142 10628
rect 36817 10625 36829 10628
rect 36863 10625 36875 10659
rect 36817 10619 36875 10625
rect 37274 10616 37280 10668
rect 37332 10616 37338 10668
rect 31478 10548 31484 10600
rect 31536 10548 31542 10600
rect 32030 10548 32036 10600
rect 32088 10548 32094 10600
rect 32401 10591 32459 10597
rect 32401 10557 32413 10591
rect 32447 10557 32459 10591
rect 32401 10551 32459 10557
rect 29932 10492 30512 10520
rect 27080 10452 27108 10492
rect 30484 10464 30512 10492
rect 30760 10492 31156 10520
rect 30760 10464 30788 10492
rect 31202 10480 31208 10532
rect 31260 10480 31266 10532
rect 31938 10520 31944 10532
rect 31726 10492 31944 10520
rect 22572 10424 27108 10452
rect 19705 10415 19763 10421
rect 28258 10412 28264 10464
rect 28316 10412 28322 10464
rect 30466 10412 30472 10464
rect 30524 10412 30530 10464
rect 30742 10412 30748 10464
rect 30800 10412 30806 10464
rect 30834 10412 30840 10464
rect 30892 10452 30898 10464
rect 31389 10455 31447 10461
rect 31389 10452 31401 10455
rect 30892 10424 31401 10452
rect 30892 10412 30898 10424
rect 31389 10421 31401 10424
rect 31435 10452 31447 10455
rect 31726 10452 31754 10492
rect 31938 10480 31944 10492
rect 31996 10520 32002 10532
rect 32416 10520 32444 10551
rect 33502 10548 33508 10600
rect 33560 10548 33566 10600
rect 36725 10591 36783 10597
rect 36725 10557 36737 10591
rect 36771 10557 36783 10591
rect 36725 10551 36783 10557
rect 31996 10492 32444 10520
rect 36740 10520 36768 10551
rect 36906 10548 36912 10600
rect 36964 10588 36970 10600
rect 39117 10591 39175 10597
rect 39117 10588 39129 10591
rect 36964 10560 39129 10588
rect 36964 10548 36970 10560
rect 39117 10557 39129 10560
rect 39163 10557 39175 10591
rect 39117 10551 39175 10557
rect 39669 10591 39727 10597
rect 39669 10557 39681 10591
rect 39715 10588 39727 10591
rect 41414 10588 41420 10600
rect 39715 10560 41420 10588
rect 39715 10557 39727 10560
rect 39669 10551 39727 10557
rect 37182 10520 37188 10532
rect 36740 10492 37188 10520
rect 31996 10480 32002 10492
rect 37182 10480 37188 10492
rect 37240 10480 37246 10532
rect 38562 10480 38568 10532
rect 38620 10520 38626 10532
rect 39684 10520 39712 10551
rect 41414 10548 41420 10560
rect 41472 10548 41478 10600
rect 38620 10492 39712 10520
rect 38620 10480 38626 10492
rect 31435 10424 31754 10452
rect 31435 10421 31447 10424
rect 31389 10415 31447 10421
rect 32858 10412 32864 10464
rect 32916 10412 32922 10464
rect 35621 10455 35679 10461
rect 35621 10421 35633 10455
rect 35667 10452 35679 10455
rect 36170 10452 36176 10464
rect 35667 10424 36176 10452
rect 35667 10421 35679 10424
rect 35621 10415 35679 10421
rect 36170 10412 36176 10424
rect 36228 10412 36234 10464
rect 37366 10412 37372 10464
rect 37424 10452 37430 10464
rect 39022 10452 39028 10464
rect 37424 10424 39028 10452
rect 37424 10412 37430 10424
rect 39022 10412 39028 10424
rect 39080 10412 39086 10464
rect 1104 10362 44620 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 44620 10362
rect 1104 10288 44620 10310
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 4706 10248 4712 10260
rect 4663 10220 4712 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 10962 10248 10968 10260
rect 10244 10220 10968 10248
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10112 10011 10115
rect 10042 10112 10048 10124
rect 9999 10084 10048 10112
rect 9999 10081 10011 10084
rect 9953 10075 10011 10081
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 5166 10004 5172 10056
rect 5224 10004 5230 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10244 10053 10272 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 19245 10251 19303 10257
rect 19245 10248 19257 10251
rect 18012 10220 19257 10248
rect 18012 10208 18018 10220
rect 19245 10217 19257 10220
rect 19291 10217 19303 10251
rect 19245 10211 19303 10217
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 21968 10220 22017 10248
rect 21968 10208 21974 10220
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22278 10248 22284 10260
rect 22005 10211 22063 10217
rect 22112 10220 22284 10248
rect 10689 10183 10747 10189
rect 10689 10149 10701 10183
rect 10735 10149 10747 10183
rect 10689 10143 10747 10149
rect 10704 10112 10732 10143
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 12618 10180 12624 10192
rect 11848 10152 12624 10180
rect 11848 10140 11854 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 15703 10152 16252 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 12066 10112 12072 10124
rect 10520 10084 12072 10112
rect 10520 10053 10548 10084
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 13262 10072 13268 10124
rect 13320 10112 13326 10124
rect 13320 10084 15792 10112
rect 13320 10072 13326 10084
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9916 10016 10149 10044
rect 9916 10004 9922 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10336 9976 10364 10007
rect 10778 10004 10784 10056
rect 10836 10044 10842 10056
rect 10873 10047 10931 10053
rect 10873 10044 10885 10047
rect 10836 10016 10885 10044
rect 10836 10004 10842 10016
rect 10873 10013 10885 10016
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11330 10044 11336 10056
rect 11112 10016 11336 10044
rect 11112 10004 11118 10016
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 14734 10044 14740 10056
rect 11572 10016 14740 10044
rect 11572 10004 11578 10016
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15764 10053 15792 10084
rect 16114 10072 16120 10124
rect 16172 10072 16178 10124
rect 16224 10121 16252 10152
rect 18782 10140 18788 10192
rect 18840 10140 18846 10192
rect 18969 10183 19027 10189
rect 18969 10149 18981 10183
rect 19015 10180 19027 10183
rect 19797 10183 19855 10189
rect 19797 10180 19809 10183
rect 19015 10152 19809 10180
rect 19015 10149 19027 10152
rect 18969 10143 19027 10149
rect 19797 10149 19809 10152
rect 19843 10149 19855 10183
rect 19797 10143 19855 10149
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 18230 10072 18236 10124
rect 18288 10072 18294 10124
rect 18800 10112 18828 10140
rect 19061 10115 19119 10121
rect 19061 10112 19073 10115
rect 18800 10084 19073 10112
rect 19061 10081 19073 10084
rect 19107 10112 19119 10115
rect 22112 10112 22140 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 27798 10208 27804 10260
rect 27856 10208 27862 10260
rect 28169 10251 28227 10257
rect 28169 10217 28181 10251
rect 28215 10217 28227 10251
rect 28169 10211 28227 10217
rect 22186 10140 22192 10192
rect 22244 10140 22250 10192
rect 22462 10140 22468 10192
rect 22520 10180 22526 10192
rect 22738 10180 22744 10192
rect 22520 10152 22744 10180
rect 22520 10140 22526 10152
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 19107 10084 22140 10112
rect 22204 10112 22232 10140
rect 22204 10084 22324 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10044 15807 10047
rect 15838 10044 15844 10056
rect 15795 10016 15844 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 9999 9948 10364 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 15470 9976 15476 9988
rect 10744 9948 15476 9976
rect 10744 9936 10750 9948
rect 15470 9936 15476 9948
rect 15528 9976 15534 9988
rect 15580 9976 15608 10007
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 15528 9948 15608 9976
rect 15528 9936 15534 9948
rect 15654 9936 15660 9988
rect 15712 9976 15718 9988
rect 15948 9976 15976 10007
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 18248 9976 18276 10072
rect 18877 10047 18935 10053
rect 18786 10025 18844 10031
rect 18786 9991 18798 10025
rect 18832 9991 18844 10025
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19150 10044 19156 10056
rect 18923 10016 19156 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19426 10047 19484 10053
rect 19426 10013 19438 10047
rect 19472 10044 19484 10047
rect 19794 10044 19800 10056
rect 19472 10016 19800 10044
rect 19472 10013 19484 10016
rect 19426 10007 19484 10013
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 19978 10044 19984 10056
rect 19935 10016 19984 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 22296 10053 22324 10084
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 22152 10016 22201 10044
rect 22152 10004 22158 10016
rect 22189 10013 22201 10016
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10044 22339 10047
rect 22557 10047 22615 10053
rect 22327 10016 22508 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 18786 9988 18844 9991
rect 22480 9988 22508 10016
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 22922 10044 22928 10056
rect 22603 10016 22928 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 22922 10004 22928 10016
rect 22980 10004 22986 10056
rect 27816 10044 27844 10208
rect 28184 10180 28212 10211
rect 28258 10208 28264 10260
rect 28316 10248 28322 10260
rect 28445 10251 28503 10257
rect 28445 10248 28457 10251
rect 28316 10220 28457 10248
rect 28316 10208 28322 10220
rect 28445 10217 28457 10220
rect 28491 10217 28503 10251
rect 28445 10211 28503 10217
rect 28626 10208 28632 10260
rect 28684 10248 28690 10260
rect 28813 10251 28871 10257
rect 28813 10248 28825 10251
rect 28684 10220 28825 10248
rect 28684 10208 28690 10220
rect 28813 10217 28825 10220
rect 28859 10248 28871 10251
rect 29270 10248 29276 10260
rect 28859 10220 29276 10248
rect 28859 10217 28871 10220
rect 28813 10211 28871 10217
rect 29270 10208 29276 10220
rect 29328 10208 29334 10260
rect 29549 10251 29607 10257
rect 29549 10217 29561 10251
rect 29595 10248 29607 10251
rect 29822 10248 29828 10260
rect 29595 10220 29828 10248
rect 29595 10217 29607 10220
rect 29549 10211 29607 10217
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 31018 10208 31024 10260
rect 31076 10248 31082 10260
rect 31481 10251 31539 10257
rect 31481 10248 31493 10251
rect 31076 10220 31493 10248
rect 31076 10208 31082 10220
rect 31481 10217 31493 10220
rect 31527 10248 31539 10251
rect 31846 10248 31852 10260
rect 31527 10220 31852 10248
rect 31527 10217 31539 10220
rect 31481 10211 31539 10217
rect 31846 10208 31852 10220
rect 31904 10208 31910 10260
rect 37274 10208 37280 10260
rect 37332 10248 37338 10260
rect 37645 10251 37703 10257
rect 37645 10248 37657 10251
rect 37332 10220 37657 10248
rect 37332 10208 37338 10220
rect 37645 10217 37657 10220
rect 37691 10248 37703 10251
rect 38102 10248 38108 10260
rect 37691 10220 38108 10248
rect 37691 10217 37703 10220
rect 37645 10211 37703 10217
rect 38102 10208 38108 10220
rect 38160 10208 38166 10260
rect 29730 10180 29736 10192
rect 28184 10152 29736 10180
rect 29730 10140 29736 10152
rect 29788 10140 29794 10192
rect 28534 10072 28540 10124
rect 28592 10072 28598 10124
rect 29270 10072 29276 10124
rect 29328 10112 29334 10124
rect 31202 10112 31208 10124
rect 29328 10084 31208 10112
rect 29328 10072 29334 10084
rect 31202 10072 31208 10084
rect 31260 10072 31266 10124
rect 39022 10072 39028 10124
rect 39080 10112 39086 10124
rect 39393 10115 39451 10121
rect 39393 10112 39405 10115
rect 39080 10084 39405 10112
rect 39080 10072 39086 10084
rect 39393 10081 39405 10084
rect 39439 10081 39451 10115
rect 39393 10075 39451 10081
rect 27893 10047 27951 10053
rect 27893 10044 27905 10047
rect 27816 10016 27905 10044
rect 27893 10013 27905 10016
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 28077 10047 28135 10053
rect 28077 10013 28089 10047
rect 28123 10044 28135 10047
rect 28442 10044 28448 10056
rect 28123 10016 28448 10044
rect 28123 10013 28135 10016
rect 28077 10007 28135 10013
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 15712 9948 18276 9976
rect 15712 9936 15718 9948
rect 18782 9936 18788 9988
rect 18840 9936 18846 9988
rect 21910 9976 21916 9988
rect 19444 9948 21916 9976
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 10376 9880 10425 9908
rect 10376 9868 10382 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 15672 9908 15700 9936
rect 11480 9880 15700 9908
rect 16393 9911 16451 9917
rect 11480 9868 11486 9880
rect 16393 9877 16405 9911
rect 16439 9908 16451 9911
rect 16666 9908 16672 9920
rect 16439 9880 16672 9908
rect 16439 9877 16451 9880
rect 16393 9871 16451 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 19444 9917 19472 9948
rect 21910 9936 21916 9948
rect 21968 9936 21974 9988
rect 22370 9936 22376 9988
rect 22428 9936 22434 9988
rect 22462 9936 22468 9988
rect 22520 9936 22526 9988
rect 28353 9979 28411 9985
rect 28353 9945 28365 9979
rect 28399 9976 28411 9979
rect 28552 9976 28580 10072
rect 28626 10004 28632 10056
rect 28684 10004 28690 10056
rect 28902 10004 28908 10056
rect 28960 10004 28966 10056
rect 30009 10047 30067 10053
rect 30009 10044 30021 10047
rect 29748 10016 30021 10044
rect 29748 9985 29776 10016
rect 30009 10013 30021 10016
rect 30055 10013 30067 10047
rect 30009 10007 30067 10013
rect 30193 10047 30251 10053
rect 30193 10013 30205 10047
rect 30239 10044 30251 10047
rect 30466 10044 30472 10056
rect 30239 10016 30472 10044
rect 30239 10013 30251 10016
rect 30193 10007 30251 10013
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 28399 9948 29745 9976
rect 28399 9945 28411 9948
rect 28353 9939 28411 9945
rect 29733 9945 29745 9948
rect 29779 9945 29791 9979
rect 29733 9939 29791 9945
rect 29917 9979 29975 9985
rect 29917 9945 29929 9979
rect 29963 9976 29975 9979
rect 30208 9976 30236 10007
rect 30466 10004 30472 10016
rect 30524 10004 30530 10056
rect 31754 10004 31760 10056
rect 31812 10044 31818 10056
rect 32953 10047 33011 10053
rect 32953 10044 32965 10047
rect 31812 10016 32965 10044
rect 31812 10004 31818 10016
rect 32953 10013 32965 10016
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 37642 10004 37648 10056
rect 37700 10044 37706 10056
rect 37700 10016 38042 10044
rect 37700 10004 37706 10016
rect 29963 9948 30236 9976
rect 39117 9979 39175 9985
rect 29963 9945 29975 9948
rect 29917 9939 29975 9945
rect 39117 9945 39129 9979
rect 39163 9976 39175 9979
rect 40862 9976 40868 9988
rect 39163 9948 40868 9976
rect 39163 9945 39175 9948
rect 39117 9939 39175 9945
rect 40862 9936 40868 9948
rect 40920 9936 40926 9988
rect 19429 9911 19487 9917
rect 19429 9877 19441 9911
rect 19475 9877 19487 9911
rect 19429 9871 19487 9877
rect 19794 9868 19800 9920
rect 19852 9908 19858 9920
rect 20622 9908 20628 9920
rect 19852 9880 20628 9908
rect 19852 9868 19858 9880
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22922 9908 22928 9920
rect 22060 9880 22928 9908
rect 22060 9868 22066 9880
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 26970 9868 26976 9920
rect 27028 9908 27034 9920
rect 27709 9911 27767 9917
rect 27709 9908 27721 9911
rect 27028 9880 27721 9908
rect 27028 9868 27034 9880
rect 27709 9877 27721 9880
rect 27755 9877 27767 9911
rect 27709 9871 27767 9877
rect 30101 9911 30159 9917
rect 30101 9877 30113 9911
rect 30147 9908 30159 9911
rect 30742 9908 30748 9920
rect 30147 9880 30748 9908
rect 30147 9877 30159 9880
rect 30101 9871 30159 9877
rect 30742 9868 30748 9880
rect 30800 9868 30806 9920
rect 31570 9868 31576 9920
rect 31628 9908 31634 9920
rect 31754 9908 31760 9920
rect 31628 9880 31760 9908
rect 31628 9868 31634 9880
rect 31754 9868 31760 9880
rect 31812 9868 31818 9920
rect 1104 9818 44620 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 44620 9818
rect 1104 9744 44620 9766
rect 2685 9707 2743 9713
rect 2685 9673 2697 9707
rect 2731 9673 2743 9707
rect 2685 9667 2743 9673
rect 4525 9707 4583 9713
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 5166 9704 5172 9716
rect 4571 9676 5172 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 2700 9636 2728 9667
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 10778 9704 10784 9716
rect 10284 9676 10784 9704
rect 10284 9664 10290 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 12176 9676 17954 9704
rect 3053 9639 3111 9645
rect 3053 9636 3065 9639
rect 2700 9608 3065 9636
rect 3053 9605 3065 9608
rect 3099 9605 3111 9639
rect 4798 9636 4804 9648
rect 4278 9608 4804 9636
rect 3053 9599 3111 9605
rect 4798 9596 4804 9608
rect 4856 9636 4862 9648
rect 5718 9636 5724 9648
rect 4856 9608 5724 9636
rect 4856 9596 4862 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 11146 9596 11152 9648
rect 11204 9596 11210 9648
rect 2498 9528 2504 9580
rect 2556 9528 2562 9580
rect 10318 9577 10324 9580
rect 10296 9571 10324 9577
rect 10296 9537 10308 9571
rect 10296 9531 10324 9537
rect 10318 9528 10324 9531
rect 10376 9528 10382 9580
rect 11164 9568 11192 9596
rect 10980 9540 11192 9568
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2792 9364 2820 9463
rect 10134 9460 10140 9512
rect 10192 9460 10198 9512
rect 10410 9460 10416 9512
rect 10468 9460 10474 9512
rect 10980 9500 11008 9540
rect 10612 9472 11008 9500
rect 4614 9432 4620 9444
rect 4448 9404 4620 9432
rect 4448 9364 4476 9404
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 2792 9336 4476 9364
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 10612 9364 10640 9472
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11333 9503 11391 9509
rect 11333 9500 11345 9503
rect 11296 9472 11345 9500
rect 11296 9460 11302 9472
rect 11333 9469 11345 9472
rect 11379 9469 11391 9503
rect 11333 9463 11391 9469
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 10962 9432 10968 9444
rect 10735 9404 10968 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 10962 9392 10968 9404
rect 11020 9432 11026 9444
rect 12176 9432 12204 9676
rect 13722 9636 13728 9648
rect 13644 9608 13728 9636
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 13262 9568 13268 9580
rect 12308 9540 13268 9568
rect 12308 9528 12314 9540
rect 13262 9528 13268 9540
rect 13320 9568 13326 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 13320 9540 13369 9568
rect 13320 9528 13326 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13541 9574 13599 9577
rect 13644 9574 13672 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13832 9580 13860 9676
rect 13998 9636 14004 9648
rect 13924 9608 14004 9636
rect 13541 9571 13672 9574
rect 13541 9537 13553 9571
rect 13587 9546 13672 9571
rect 13587 9537 13599 9546
rect 13541 9531 13599 9537
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 13924 9500 13952 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14277 9639 14335 9645
rect 14277 9636 14289 9639
rect 14240 9608 14289 9636
rect 14240 9596 14246 9608
rect 14277 9605 14289 9608
rect 14323 9605 14335 9639
rect 14277 9599 14335 9605
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 17926 9636 17954 9676
rect 18322 9664 18328 9716
rect 18380 9704 18386 9716
rect 20162 9704 20168 9716
rect 18380 9676 20168 9704
rect 18380 9664 18386 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 21324 9676 21864 9704
rect 21324 9664 21330 9676
rect 18046 9636 18052 9648
rect 14700 9608 16160 9636
rect 17926 9608 18052 9636
rect 14700 9596 14706 9608
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9568 14151 9571
rect 14139 9558 14228 9568
rect 14366 9558 14372 9580
rect 14139 9540 14372 9558
rect 14139 9537 14151 9540
rect 14093 9531 14151 9537
rect 14200 9530 14372 9540
rect 14366 9528 14372 9530
rect 14424 9528 14430 9580
rect 16132 9577 16160 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 21542 9596 21548 9648
rect 21600 9596 21606 9648
rect 21836 9645 21864 9676
rect 21910 9664 21916 9716
rect 21968 9704 21974 9716
rect 23201 9707 23259 9713
rect 23201 9704 23213 9707
rect 21968 9676 23213 9704
rect 21968 9664 21974 9676
rect 23201 9673 23213 9676
rect 23247 9673 23259 9707
rect 23201 9667 23259 9673
rect 23569 9707 23627 9713
rect 23569 9673 23581 9707
rect 23615 9704 23627 9707
rect 23934 9704 23940 9716
rect 23615 9676 23940 9704
rect 23615 9673 23627 9676
rect 23569 9667 23627 9673
rect 23934 9664 23940 9676
rect 23992 9704 23998 9716
rect 24305 9707 24363 9713
rect 24305 9704 24317 9707
rect 23992 9676 24317 9704
rect 23992 9664 23998 9676
rect 24305 9673 24317 9676
rect 24351 9673 24363 9707
rect 24305 9667 24363 9673
rect 24670 9664 24676 9716
rect 24728 9704 24734 9716
rect 24765 9707 24823 9713
rect 24765 9704 24777 9707
rect 24728 9676 24777 9704
rect 24728 9664 24734 9676
rect 24765 9673 24777 9676
rect 24811 9673 24823 9707
rect 24765 9667 24823 9673
rect 26237 9707 26295 9713
rect 26237 9673 26249 9707
rect 26283 9704 26295 9707
rect 27338 9704 27344 9716
rect 26283 9676 27344 9704
rect 26283 9673 26295 9676
rect 26237 9667 26295 9673
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 28902 9664 28908 9716
rect 28960 9704 28966 9716
rect 31386 9704 31392 9716
rect 28960 9676 31392 9704
rect 28960 9664 28966 9676
rect 31386 9664 31392 9676
rect 31444 9664 31450 9716
rect 40862 9664 40868 9716
rect 40920 9664 40926 9716
rect 21821 9639 21879 9645
rect 21821 9605 21833 9639
rect 21867 9605 21879 9639
rect 23382 9636 23388 9648
rect 21821 9599 21879 9605
rect 21928 9608 23388 9636
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16574 9568 16580 9580
rect 16255 9540 16580 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16724 9540 16865 9568
rect 16724 9528 16730 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17402 9568 17408 9580
rect 17359 9540 17408 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18598 9568 18604 9580
rect 17644 9540 18604 9568
rect 17644 9528 17650 9540
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 20346 9568 20352 9580
rect 19024 9540 20352 9568
rect 19024 9528 19030 9540
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 21560 9568 21588 9596
rect 21928 9580 21956 9608
rect 23382 9596 23388 9608
rect 23440 9636 23446 9648
rect 32858 9636 32864 9648
rect 23440 9608 23704 9636
rect 23440 9596 23446 9608
rect 21910 9568 21916 9580
rect 21560 9540 21916 9568
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 22060 9540 22109 9568
rect 22060 9528 22066 9540
rect 22097 9537 22109 9540
rect 22143 9568 22155 9571
rect 23676 9568 23704 9608
rect 28644 9608 32864 9636
rect 28644 9577 28672 9608
rect 32858 9596 32864 9608
rect 32916 9596 32922 9648
rect 42518 9596 42524 9648
rect 42576 9596 42582 9648
rect 24673 9571 24731 9577
rect 22143 9540 22692 9568
rect 23676 9540 23796 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 13771 9472 13952 9500
rect 14001 9503 14059 9509
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 15838 9500 15844 9512
rect 14047 9472 15844 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9492 16083 9503
rect 16071 9469 16252 9492
rect 16025 9464 16252 9469
rect 16025 9463 16083 9464
rect 11020 9404 12204 9432
rect 13633 9435 13691 9441
rect 11020 9392 11026 9404
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 14090 9432 14096 9444
rect 13679 9404 14096 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 14090 9392 14096 9404
rect 14148 9392 14154 9444
rect 16224 9432 16252 9464
rect 16298 9460 16304 9512
rect 16356 9460 16362 9512
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 20530 9500 20536 9512
rect 16540 9472 20536 9500
rect 16540 9460 16546 9472
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21450 9500 21456 9512
rect 20772 9472 21456 9500
rect 20772 9460 20778 9472
rect 21450 9460 21456 9472
rect 21508 9500 21514 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21508 9472 21833 9500
rect 21508 9460 21514 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 22664 9444 22692 9540
rect 23658 9460 23664 9512
rect 23716 9460 23722 9512
rect 23768 9509 23796 9540
rect 24673 9537 24685 9571
rect 24719 9568 24731 9571
rect 26145 9571 26203 9577
rect 24719 9540 24808 9568
rect 24719 9537 24731 9540
rect 24673 9531 24731 9537
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9469 23811 9503
rect 23753 9463 23811 9469
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 16224 9404 16681 9432
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 22094 9432 22100 9444
rect 16669 9395 16727 9401
rect 19306 9404 22100 9432
rect 9539 9336 10640 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14240 9336 14473 9364
rect 14240 9324 14246 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 16485 9367 16543 9373
rect 16485 9333 16497 9367
rect 16531 9364 16543 9367
rect 19306 9364 19334 9404
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 22646 9392 22652 9444
rect 22704 9432 22710 9444
rect 22830 9432 22836 9444
rect 22704 9404 22836 9432
rect 22704 9392 22710 9404
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 24780 9376 24808 9540
rect 26145 9537 26157 9571
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9537 28687 9571
rect 28629 9531 28687 9537
rect 28721 9571 28779 9577
rect 28721 9537 28733 9571
rect 28767 9537 28779 9571
rect 28721 9531 28779 9537
rect 24949 9503 25007 9509
rect 24949 9469 24961 9503
rect 24995 9500 25007 9503
rect 25222 9500 25228 9512
rect 24995 9472 25228 9500
rect 24995 9469 25007 9472
rect 24949 9463 25007 9469
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 26160 9376 26188 9531
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9500 26479 9503
rect 26602 9500 26608 9512
rect 26467 9472 26608 9500
rect 26467 9469 26479 9472
rect 26421 9463 26479 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 28534 9460 28540 9512
rect 28592 9460 28598 9512
rect 28736 9500 28764 9531
rect 28902 9528 28908 9580
rect 28960 9528 28966 9580
rect 28997 9571 29055 9577
rect 28997 9537 29009 9571
rect 29043 9537 29055 9571
rect 28997 9531 29055 9537
rect 29181 9571 29239 9577
rect 29181 9537 29193 9571
rect 29227 9537 29239 9571
rect 29181 9531 29239 9537
rect 29012 9500 29040 9531
rect 28736 9472 29040 9500
rect 29196 9500 29224 9531
rect 29270 9528 29276 9580
rect 29328 9528 29334 9580
rect 29457 9571 29515 9577
rect 29457 9537 29469 9571
rect 29503 9568 29515 9571
rect 29546 9568 29552 9580
rect 29503 9540 29552 9568
rect 29503 9537 29515 9540
rect 29457 9531 29515 9537
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 30650 9528 30656 9580
rect 30708 9528 30714 9580
rect 30834 9528 30840 9580
rect 30892 9528 30898 9580
rect 31481 9571 31539 9577
rect 31481 9537 31493 9571
rect 31527 9568 31539 9571
rect 32030 9568 32036 9580
rect 31527 9540 32036 9568
rect 31527 9537 31539 9540
rect 31481 9531 31539 9537
rect 32030 9528 32036 9540
rect 32088 9528 32094 9580
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 30006 9500 30012 9512
rect 29196 9472 30012 9500
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 28261 9435 28319 9441
rect 28261 9432 28273 9435
rect 27396 9404 28273 9432
rect 27396 9392 27402 9404
rect 28261 9401 28273 9404
rect 28307 9401 28319 9435
rect 28966 9432 28994 9472
rect 30006 9460 30012 9472
rect 30064 9500 30070 9512
rect 31297 9503 31355 9509
rect 31297 9500 31309 9503
rect 30064 9472 31309 9500
rect 30064 9460 30070 9472
rect 31297 9469 31309 9472
rect 31343 9469 31355 9503
rect 31297 9463 31355 9469
rect 31662 9460 31668 9512
rect 31720 9460 31726 9512
rect 31754 9460 31760 9512
rect 31812 9460 31818 9512
rect 28966 9404 29592 9432
rect 28261 9395 28319 9401
rect 16531 9336 19334 9364
rect 16531 9333 16543 9336
rect 16485 9327 16543 9333
rect 21726 9324 21732 9376
rect 21784 9364 21790 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21784 9336 22017 9364
rect 21784 9324 21790 9336
rect 22005 9333 22017 9336
rect 22051 9364 22063 9367
rect 24394 9364 24400 9376
rect 22051 9336 24400 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 24762 9324 24768 9376
rect 24820 9324 24826 9376
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25498 9364 25504 9376
rect 24912 9336 25504 9364
rect 24912 9324 24918 9336
rect 25498 9324 25504 9336
rect 25556 9364 25562 9376
rect 25777 9367 25835 9373
rect 25777 9364 25789 9367
rect 25556 9336 25789 9364
rect 25556 9324 25562 9336
rect 25777 9333 25789 9336
rect 25823 9333 25835 9367
rect 25777 9327 25835 9333
rect 26142 9324 26148 9376
rect 26200 9324 26206 9376
rect 28442 9324 28448 9376
rect 28500 9364 28506 9376
rect 28721 9367 28779 9373
rect 28721 9364 28733 9367
rect 28500 9336 28733 9364
rect 28500 9324 28506 9336
rect 28721 9333 28733 9336
rect 28767 9333 28779 9367
rect 28721 9327 28779 9333
rect 28810 9324 28816 9376
rect 28868 9364 28874 9376
rect 29564 9373 29592 9404
rect 30466 9392 30472 9444
rect 30524 9432 30530 9444
rect 30745 9435 30803 9441
rect 30745 9432 30757 9435
rect 30524 9404 30757 9432
rect 30524 9392 30530 9404
rect 30745 9401 30757 9404
rect 30791 9401 30803 9435
rect 32140 9432 32168 9531
rect 32214 9528 32220 9580
rect 32272 9568 32278 9580
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 32272 9540 32321 9568
rect 32272 9528 32278 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 33689 9503 33747 9509
rect 33689 9469 33701 9503
rect 33735 9500 33747 9503
rect 38562 9500 38568 9512
rect 33735 9472 38568 9500
rect 33735 9469 33747 9472
rect 33689 9463 33747 9469
rect 30745 9395 30803 9401
rect 31588 9404 32168 9432
rect 31588 9376 31616 9404
rect 33962 9392 33968 9444
rect 34020 9392 34026 9444
rect 34072 9376 34100 9472
rect 38562 9460 38568 9472
rect 38620 9460 38626 9512
rect 41506 9460 41512 9512
rect 41564 9460 41570 9512
rect 29089 9367 29147 9373
rect 29089 9364 29101 9367
rect 28868 9336 29101 9364
rect 28868 9324 28874 9336
rect 29089 9333 29101 9336
rect 29135 9333 29147 9367
rect 29089 9327 29147 9333
rect 29549 9367 29607 9373
rect 29549 9333 29561 9367
rect 29595 9364 29607 9367
rect 29638 9364 29644 9376
rect 29595 9336 29644 9364
rect 29595 9333 29607 9336
rect 29549 9327 29607 9333
rect 29638 9324 29644 9336
rect 29696 9324 29702 9376
rect 30834 9324 30840 9376
rect 30892 9364 30898 9376
rect 31202 9364 31208 9376
rect 30892 9336 31208 9364
rect 30892 9324 30898 9336
rect 31202 9324 31208 9336
rect 31260 9324 31266 9376
rect 31570 9324 31576 9376
rect 31628 9324 31634 9376
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 31938 9364 31944 9376
rect 31812 9336 31944 9364
rect 31812 9324 31818 9336
rect 31938 9324 31944 9336
rect 31996 9364 32002 9376
rect 32217 9367 32275 9373
rect 32217 9364 32229 9367
rect 31996 9336 32229 9364
rect 31996 9324 32002 9336
rect 32217 9333 32229 9336
rect 32263 9333 32275 9367
rect 32217 9327 32275 9333
rect 34054 9324 34060 9376
rect 34112 9324 34118 9376
rect 34146 9324 34152 9376
rect 34204 9324 34210 9376
rect 43714 9324 43720 9376
rect 43772 9364 43778 9376
rect 43809 9367 43867 9373
rect 43809 9364 43821 9367
rect 43772 9336 43821 9364
rect 43772 9324 43778 9336
rect 43809 9333 43821 9336
rect 43855 9364 43867 9367
rect 44266 9364 44272 9376
rect 43855 9336 44272 9364
rect 43855 9333 43867 9336
rect 43809 9327 43867 9333
rect 44266 9324 44272 9336
rect 44324 9324 44330 9376
rect 1104 9274 44620 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 44620 9274
rect 1104 9200 44620 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2498 9160 2504 9172
rect 2271 9132 2504 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9160 9827 9163
rect 10410 9160 10416 9172
rect 9815 9132 10416 9160
rect 9815 9129 9827 9132
rect 9769 9123 9827 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10594 9120 10600 9172
rect 10652 9120 10658 9172
rect 10686 9120 10692 9172
rect 10744 9120 10750 9172
rect 11238 9120 11244 9172
rect 11296 9120 11302 9172
rect 11514 9120 11520 9172
rect 11572 9120 11578 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 12032 9132 12081 9160
rect 12032 9120 12038 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12710 9160 12716 9172
rect 12584 9132 12716 9160
rect 12584 9120 12590 9132
rect 12710 9120 12716 9132
rect 12768 9160 12774 9172
rect 13630 9160 13636 9172
rect 12768 9132 13636 9160
rect 12768 9120 12774 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 13998 9160 14004 9172
rect 13955 9132 14004 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14090 9120 14096 9172
rect 14148 9120 14154 9172
rect 14366 9160 14372 9172
rect 14200 9132 14372 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2041 9095 2099 9101
rect 2041 9092 2053 9095
rect 1627 9064 2053 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2041 9061 2053 9064
rect 2087 9061 2099 9095
rect 9674 9092 9680 9104
rect 2041 9055 2099 9061
rect 6656 9064 9680 9092
rect 1762 8984 1768 9036
rect 1820 8984 1826 9036
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 6656 8965 6684 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 10042 9052 10048 9104
rect 10100 9052 10106 9104
rect 10612 9092 10640 9120
rect 11532 9092 11560 9120
rect 13170 9092 13176 9104
rect 10612 9064 11560 9092
rect 11624 9064 13176 9092
rect 6730 8984 6736 9036
rect 6788 8984 6794 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7374 9024 7380 9036
rect 7331 8996 7380 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 7024 8956 7052 8987
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 10060 9024 10088 9052
rect 7760 8996 10088 9024
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7024 8928 7481 8956
rect 6641 8919 6699 8925
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7377 8891 7435 8897
rect 7377 8888 7389 8891
rect 7156 8860 7389 8888
rect 7156 8848 7162 8860
rect 7377 8857 7389 8860
rect 7423 8888 7435 8891
rect 7760 8888 7788 8996
rect 9968 8965 9996 8996
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 11624 9024 11652 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 13357 9095 13415 9101
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 14200 9092 14228 9132
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 14476 9132 14657 9160
rect 13403 9064 14228 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 10980 8996 11652 9024
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7423 8860 7788 8888
rect 7852 8928 8125 8956
rect 7423 8857 7435 8860
rect 7377 8851 7435 8857
rect 7852 8829 7880 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10520 8956 10548 8984
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10520 8928 10885 8956
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 10410 8888 10416 8900
rect 10367 8860 10416 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 10502 8848 10508 8900
rect 10560 8848 10566 8900
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 7926 8780 7932 8832
rect 7984 8780 7990 8832
rect 10428 8820 10456 8848
rect 10980 8820 11008 8996
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11103 8928 11376 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11348 8829 11376 8928
rect 11514 8916 11520 8968
rect 11572 8916 11578 8968
rect 11624 8956 11652 8996
rect 12084 8996 12909 9024
rect 11695 8959 11753 8965
rect 11695 8956 11707 8959
rect 11624 8928 11707 8956
rect 11695 8925 11707 8928
rect 11741 8925 11753 8959
rect 11695 8919 11753 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12084 8956 12112 8996
rect 12897 8993 12909 8996
rect 12943 9024 12955 9027
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 12943 8996 13553 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 13541 8993 13553 8996
rect 13587 9024 13599 9027
rect 14476 9024 14504 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 16298 9120 16304 9172
rect 16356 9120 16362 9172
rect 16853 9163 16911 9169
rect 16853 9129 16865 9163
rect 16899 9160 16911 9163
rect 17126 9160 17132 9172
rect 16899 9132 17132 9160
rect 16899 9129 16911 9132
rect 16853 9123 16911 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 18690 9160 18696 9172
rect 17460 9132 17632 9160
rect 17460 9120 17466 9132
rect 15562 9052 15568 9104
rect 15620 9092 15626 9104
rect 16316 9092 16344 9120
rect 17604 9104 17632 9132
rect 17880 9132 18696 9160
rect 16945 9095 17003 9101
rect 16945 9092 16957 9095
rect 15620 9064 16252 9092
rect 16316 9064 16957 9092
rect 15620 9052 15626 9064
rect 16224 9033 16252 9064
rect 16945 9061 16957 9064
rect 16991 9061 17003 9095
rect 16945 9055 17003 9061
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 17276 9064 17540 9092
rect 17276 9052 17282 9064
rect 16209 9027 16267 9033
rect 13587 8996 14504 9024
rect 14936 8996 16160 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 14936 8968 14964 8996
rect 12023 8928 12112 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12084 8832 12112 8928
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 10428 8792 11008 8820
rect 11333 8823 11391 8829
rect 11333 8789 11345 8823
rect 11379 8789 11391 8823
rect 11333 8783 11391 8789
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 13188 8820 13216 8919
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13412 8928 13461 8956
rect 13412 8916 13418 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13688 8928 13737 8956
rect 13688 8916 13694 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 14240 8928 14289 8956
rect 14240 8916 14246 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 14424 8928 14473 8956
rect 14424 8916 14430 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14550 8916 14556 8968
rect 14608 8916 14614 8968
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 14660 8888 14688 8919
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16022 8956 16028 8968
rect 15979 8928 16028 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16132 8965 16160 8996
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 17512 9024 17540 9064
rect 17586 9052 17592 9104
rect 17644 9052 17650 9104
rect 17880 9024 17908 9132
rect 17954 9052 17960 9104
rect 18012 9052 18018 9104
rect 18049 9095 18107 9101
rect 18049 9061 18061 9095
rect 18095 9061 18107 9095
rect 18049 9055 18107 9061
rect 18064 9024 18092 9055
rect 16632 8996 17448 9024
rect 17512 8996 17908 9024
rect 17972 8996 18092 9024
rect 16632 8984 16638 8996
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 16298 8916 16304 8968
rect 16356 8916 16362 8968
rect 16728 8959 16786 8965
rect 16728 8925 16740 8959
rect 16774 8956 16786 8959
rect 17129 8959 17187 8965
rect 16774 8928 17080 8956
rect 16774 8925 16786 8928
rect 16728 8919 16786 8925
rect 16942 8888 16948 8900
rect 13320 8860 14688 8888
rect 15028 8860 16948 8888
rect 13320 8848 13326 8860
rect 13998 8820 14004 8832
rect 13188 8792 14004 8820
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 15028 8829 15056 8860
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 15013 8823 15071 8829
rect 15013 8789 15025 8823
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 16025 8823 16083 8829
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16071 8792 16681 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 17052 8820 17080 8928
rect 17129 8925 17141 8959
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17144 8888 17172 8919
rect 17218 8916 17224 8968
rect 17276 8916 17282 8968
rect 17420 8965 17448 8996
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17586 8956 17592 8968
rect 17543 8928 17592 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 17972 8965 18000 8996
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8956 17739 8959
rect 17957 8959 18015 8965
rect 17727 8928 17908 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 17310 8888 17316 8900
rect 17144 8860 17316 8888
rect 17310 8848 17316 8860
rect 17368 8888 17374 8900
rect 17880 8888 17908 8928
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 18156 8956 18184 9132
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 19334 9120 19340 9172
rect 19392 9120 19398 9172
rect 19889 9163 19947 9169
rect 19889 9129 19901 9163
rect 19935 9160 19947 9163
rect 19978 9160 19984 9172
rect 19935 9132 19984 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20162 9120 20168 9172
rect 20220 9160 20226 9172
rect 20530 9160 20536 9172
rect 20220 9132 20536 9160
rect 20220 9120 20226 9132
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 22189 9163 22247 9169
rect 22189 9129 22201 9163
rect 22235 9160 22247 9163
rect 22278 9160 22284 9172
rect 22235 9132 22284 9160
rect 22235 9129 22247 9132
rect 22189 9123 22247 9129
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22428 9132 22753 9160
rect 22428 9120 22434 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 24394 9120 24400 9172
rect 24452 9120 24458 9172
rect 24670 9120 24676 9172
rect 24728 9160 24734 9172
rect 25685 9163 25743 9169
rect 25685 9160 25697 9163
rect 24728 9132 25697 9160
rect 24728 9120 24734 9132
rect 25685 9129 25697 9132
rect 25731 9129 25743 9163
rect 25685 9123 25743 9129
rect 27798 9120 27804 9172
rect 27856 9160 27862 9172
rect 30377 9163 30435 9169
rect 30377 9160 30389 9163
rect 27856 9132 30389 9160
rect 27856 9120 27862 9132
rect 30377 9129 30389 9132
rect 30423 9129 30435 9163
rect 30377 9123 30435 9129
rect 30650 9120 30656 9172
rect 30708 9160 30714 9172
rect 31478 9160 31484 9172
rect 30708 9132 31484 9160
rect 30708 9120 30714 9132
rect 31478 9120 31484 9132
rect 31536 9120 31542 9172
rect 33032 9163 33090 9169
rect 33032 9129 33044 9163
rect 33078 9160 33090 9163
rect 36906 9160 36912 9172
rect 33078 9132 36912 9160
rect 33078 9129 33090 9132
rect 33032 9123 33090 9129
rect 36906 9120 36912 9132
rect 36964 9120 36970 9172
rect 18230 9052 18236 9104
rect 18288 9052 18294 9104
rect 18248 9024 18276 9052
rect 18248 8996 18460 9024
rect 17957 8919 18015 8925
rect 18064 8928 18184 8956
rect 18064 8897 18092 8928
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18432 8965 18460 8996
rect 18708 8965 18736 9120
rect 18782 9052 18788 9104
rect 18840 9052 18846 9104
rect 19352 9092 19380 9120
rect 20441 9095 20499 9101
rect 20441 9092 20453 9095
rect 19352 9064 20453 9092
rect 20441 9061 20453 9064
rect 20487 9061 20499 9095
rect 20441 9055 20499 9061
rect 22002 9052 22008 9104
rect 22060 9052 22066 9104
rect 22462 9052 22468 9104
rect 22520 9052 22526 9104
rect 22646 9092 22652 9104
rect 22572 9064 22652 9092
rect 18800 9024 18828 9052
rect 18969 9027 19027 9033
rect 18800 8996 18920 9024
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8925 18843 8959
rect 18892 8956 18920 8996
rect 18969 8993 18981 9027
rect 19015 9024 19027 9027
rect 20533 9027 20591 9033
rect 19015 8996 19472 9024
rect 19015 8993 19027 8996
rect 18969 8987 19027 8993
rect 19444 8965 19472 8996
rect 20533 8993 20545 9027
rect 20579 9024 20591 9027
rect 21545 9027 21603 9033
rect 21545 9024 21557 9027
rect 20579 8996 21557 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 21545 8993 21557 8996
rect 21591 8993 21603 9027
rect 22020 9024 22048 9052
rect 22480 9024 22508 9052
rect 22572 9033 22600 9064
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 24762 9052 24768 9104
rect 24820 9092 24826 9104
rect 26513 9095 26571 9101
rect 26513 9092 26525 9095
rect 24820 9064 26525 9092
rect 24820 9052 24826 9064
rect 21545 8987 21603 8993
rect 21836 8996 22048 9024
rect 22112 8996 22508 9024
rect 22557 9027 22615 9033
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18892 8928 19257 8956
rect 18785 8919 18843 8925
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 19978 8956 19984 8968
rect 19659 8928 19984 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 17368 8860 17908 8888
rect 17368 8848 17374 8860
rect 17402 8820 17408 8832
rect 17052 8792 17408 8820
rect 16669 8783 16727 8789
rect 17402 8780 17408 8792
rect 17460 8780 17466 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17644 8792 17785 8820
rect 17644 8780 17650 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17880 8820 17908 8860
rect 18049 8891 18107 8897
rect 18049 8857 18061 8891
rect 18095 8857 18107 8891
rect 18524 8888 18552 8919
rect 18800 8888 18828 8919
rect 18049 8851 18107 8857
rect 18156 8860 18552 8888
rect 18616 8860 18828 8888
rect 18156 8820 18184 8860
rect 18616 8832 18644 8860
rect 17880 8792 18184 8820
rect 18233 8823 18291 8829
rect 17773 8783 17831 8789
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18322 8820 18328 8832
rect 18279 8792 18328 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18598 8780 18604 8832
rect 18656 8780 18662 8832
rect 19260 8820 19288 8919
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19536 8888 19564 8919
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 19392 8860 19564 8888
rect 20272 8888 20300 8919
rect 20346 8916 20352 8968
rect 20404 8916 20410 8968
rect 20622 8916 20628 8968
rect 20680 8916 20686 8968
rect 21726 8916 21732 8968
rect 21784 8916 21790 8968
rect 21836 8965 21864 8996
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 22112 8965 22140 8996
rect 22557 8993 22569 9027
rect 22603 8993 22615 9027
rect 23014 9024 23020 9036
rect 22557 8987 22615 8993
rect 22664 8996 23020 9024
rect 22664 8965 22692 8996
rect 23014 8984 23020 8996
rect 23072 9024 23078 9036
rect 23474 9024 23480 9036
rect 23072 8996 23480 9024
rect 23072 8984 23078 8996
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 24872 9033 24900 9064
rect 26513 9061 26525 9064
rect 26559 9061 26571 9095
rect 26513 9055 26571 9061
rect 30466 9052 30472 9104
rect 30524 9092 30530 9104
rect 30524 9064 30972 9092
rect 30524 9052 30530 9064
rect 24857 9027 24915 9033
rect 24857 8993 24869 9027
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 25041 9027 25099 9033
rect 25041 8993 25053 9027
rect 25087 9024 25099 9027
rect 25222 9024 25228 9036
rect 25087 8996 25228 9024
rect 25087 8993 25099 8996
rect 25041 8987 25099 8993
rect 25222 8984 25228 8996
rect 25280 8984 25286 9036
rect 26329 9027 26387 9033
rect 26329 8993 26341 9027
rect 26375 9024 26387 9027
rect 26602 9024 26608 9036
rect 26375 8996 26608 9024
rect 26375 8993 26387 8996
rect 26329 8987 26387 8993
rect 26602 8984 26608 8996
rect 26660 8984 26666 9036
rect 26970 8984 26976 9036
rect 27028 8984 27034 9036
rect 27157 9027 27215 9033
rect 27157 8993 27169 9027
rect 27203 9024 27215 9027
rect 27246 9024 27252 9036
rect 27203 8996 27252 9024
rect 27203 8993 27215 8996
rect 27157 8987 27215 8993
rect 27246 8984 27252 8996
rect 27304 8984 27310 9036
rect 29730 8984 29736 9036
rect 29788 9024 29794 9036
rect 30944 9024 30972 9064
rect 31018 9052 31024 9104
rect 31076 9092 31082 9104
rect 31570 9092 31576 9104
rect 31076 9064 31576 9092
rect 31076 9052 31082 9064
rect 31570 9052 31576 9064
rect 31628 9052 31634 9104
rect 31113 9027 31171 9033
rect 31113 9024 31125 9027
rect 29788 8996 30788 9024
rect 30944 8996 31125 9024
rect 29788 8984 29794 8996
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22373 8959 22431 8965
rect 22373 8925 22385 8959
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8956 22891 8959
rect 22879 8928 23520 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 20640 8888 20668 8916
rect 20272 8860 20668 8888
rect 22388 8888 22416 8919
rect 22388 8860 22692 8888
rect 19392 8848 19398 8860
rect 22664 8832 22692 8860
rect 23492 8832 23520 8928
rect 26142 8916 26148 8968
rect 26200 8956 26206 8968
rect 27617 8959 27675 8965
rect 27617 8956 27629 8959
rect 26200 8928 27629 8956
rect 26200 8916 26206 8928
rect 27617 8925 27629 8928
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 27706 8916 27712 8968
rect 27764 8956 27770 8968
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27764 8928 27813 8956
rect 27764 8916 27770 8928
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27801 8919 27859 8925
rect 27890 8916 27896 8968
rect 27948 8916 27954 8968
rect 29270 8916 29276 8968
rect 29328 8956 29334 8968
rect 30101 8959 30159 8965
rect 30101 8956 30113 8959
rect 29328 8928 30113 8956
rect 29328 8916 29334 8928
rect 30101 8925 30113 8928
rect 30147 8925 30159 8959
rect 30101 8919 30159 8925
rect 30285 8959 30343 8965
rect 30285 8925 30297 8959
rect 30331 8956 30343 8959
rect 30374 8956 30380 8968
rect 30331 8928 30380 8956
rect 30331 8925 30343 8928
rect 30285 8919 30343 8925
rect 30374 8916 30380 8928
rect 30432 8956 30438 8968
rect 30561 8959 30619 8965
rect 30561 8956 30573 8959
rect 30432 8928 30573 8956
rect 30432 8916 30438 8928
rect 30561 8925 30573 8928
rect 30607 8925 30619 8959
rect 30760 8958 30788 8996
rect 31113 8993 31125 8996
rect 31159 8993 31171 9027
rect 31113 8987 31171 8993
rect 31202 8984 31208 9036
rect 31260 8984 31266 9036
rect 30929 8959 30987 8965
rect 30760 8950 30880 8958
rect 30929 8950 30941 8959
rect 30760 8930 30941 8950
rect 30561 8919 30619 8925
rect 30852 8925 30941 8930
rect 30975 8925 30987 8959
rect 30852 8922 30987 8925
rect 30929 8919 30987 8922
rect 31021 8953 31079 8959
rect 31220 8956 31248 8984
rect 31588 8965 31616 9052
rect 32769 9027 32827 9033
rect 32769 8993 32781 9027
rect 32815 9024 32827 9027
rect 33134 9024 33140 9036
rect 32815 8996 33140 9024
rect 32815 8993 32827 8996
rect 32769 8987 32827 8993
rect 33134 8984 33140 8996
rect 33192 9024 33198 9036
rect 33502 9024 33508 9036
rect 33192 8996 33508 9024
rect 33192 8984 33198 8996
rect 33502 8984 33508 8996
rect 33560 8984 33566 9036
rect 35069 9027 35127 9033
rect 35069 8993 35081 9027
rect 35115 9024 35127 9027
rect 35342 9024 35348 9036
rect 35115 8996 35348 9024
rect 35115 8993 35127 8996
rect 35069 8987 35127 8993
rect 35342 8984 35348 8996
rect 35400 8984 35406 9036
rect 31021 8919 31033 8953
rect 31067 8950 31079 8953
rect 31128 8950 31248 8956
rect 31067 8928 31248 8950
rect 31573 8959 31631 8965
rect 31067 8922 31156 8928
rect 31573 8925 31585 8959
rect 31619 8925 31631 8959
rect 31067 8919 31079 8922
rect 31573 8919 31631 8925
rect 31021 8913 31079 8919
rect 31662 8916 31668 8968
rect 31720 8916 31726 8968
rect 36909 8959 36967 8965
rect 36909 8956 36921 8959
rect 36832 8928 36921 8956
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8888 24823 8891
rect 24946 8888 24952 8900
rect 24811 8860 24952 8888
rect 24811 8857 24823 8860
rect 24765 8851 24823 8857
rect 24946 8848 24952 8860
rect 25004 8888 25010 8900
rect 25004 8860 25912 8888
rect 25004 8848 25010 8860
rect 25884 8832 25912 8860
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 29178 8888 29184 8900
rect 28224 8860 29184 8888
rect 28224 8848 28230 8860
rect 29178 8848 29184 8860
rect 29236 8848 29242 8900
rect 30193 8891 30251 8897
rect 30193 8857 30205 8891
rect 30239 8888 30251 8891
rect 30466 8888 30472 8900
rect 30239 8860 30472 8888
rect 30239 8857 30251 8860
rect 30193 8851 30251 8857
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 30650 8848 30656 8900
rect 30708 8848 30714 8900
rect 30745 8891 30803 8897
rect 30745 8857 30757 8891
rect 30791 8857 30803 8891
rect 30745 8851 30803 8857
rect 20162 8820 20168 8832
rect 19260 8792 20168 8820
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 22646 8780 22652 8832
rect 22704 8780 22710 8832
rect 23474 8780 23480 8832
rect 23532 8780 23538 8832
rect 25866 8780 25872 8832
rect 25924 8780 25930 8832
rect 26053 8823 26111 8829
rect 26053 8789 26065 8823
rect 26099 8820 26111 8823
rect 26326 8820 26332 8832
rect 26099 8792 26332 8820
rect 26099 8789 26111 8792
rect 26053 8783 26111 8789
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26878 8780 26884 8832
rect 26936 8780 26942 8832
rect 27985 8823 28043 8829
rect 27985 8789 27997 8823
rect 28031 8820 28043 8823
rect 29638 8820 29644 8832
rect 28031 8792 29644 8820
rect 28031 8789 28043 8792
rect 27985 8783 28043 8789
rect 29638 8780 29644 8792
rect 29696 8780 29702 8832
rect 30760 8820 30788 8851
rect 31110 8820 31116 8832
rect 30760 8792 31116 8820
rect 31110 8780 31116 8792
rect 31168 8820 31174 8832
rect 31680 8820 31708 8916
rect 34790 8888 34796 8900
rect 34270 8860 34796 8888
rect 34790 8848 34796 8860
rect 34848 8888 34854 8900
rect 35345 8891 35403 8897
rect 34848 8860 35296 8888
rect 34848 8848 34854 8860
rect 31168 8792 31708 8820
rect 31168 8780 31174 8792
rect 34514 8780 34520 8832
rect 34572 8780 34578 8832
rect 35268 8820 35296 8860
rect 35345 8857 35357 8891
rect 35391 8888 35403 8891
rect 35434 8888 35440 8900
rect 35391 8860 35440 8888
rect 35391 8857 35403 8860
rect 35345 8851 35403 8857
rect 35434 8848 35440 8860
rect 35492 8848 35498 8900
rect 35728 8860 35834 8888
rect 35728 8820 35756 8860
rect 35268 8792 35756 8820
rect 36078 8780 36084 8832
rect 36136 8820 36142 8832
rect 36832 8829 36860 8928
rect 36909 8925 36921 8928
rect 36955 8925 36967 8959
rect 36909 8919 36967 8925
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8956 37611 8959
rect 37645 8959 37703 8965
rect 37645 8956 37657 8959
rect 37599 8928 37657 8956
rect 37599 8925 37611 8928
rect 37553 8919 37611 8925
rect 37645 8925 37657 8928
rect 37691 8925 37703 8959
rect 37645 8919 37703 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8956 37887 8959
rect 37918 8956 37924 8968
rect 37875 8928 37924 8956
rect 37875 8925 37887 8928
rect 37829 8919 37887 8925
rect 37918 8916 37924 8928
rect 37976 8916 37982 8968
rect 36817 8823 36875 8829
rect 36817 8820 36829 8823
rect 36136 8792 36829 8820
rect 36136 8780 36142 8792
rect 36817 8789 36829 8792
rect 36863 8789 36875 8823
rect 36817 8783 36875 8789
rect 37734 8780 37740 8832
rect 37792 8780 37798 8832
rect 1104 8730 44620 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 44620 8730
rect 1104 8656 44620 8678
rect 10134 8576 10140 8628
rect 10192 8576 10198 8628
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10284 8588 10425 8616
rect 10284 8576 10290 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 11514 8616 11520 8628
rect 10735 8588 11520 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12952 8588 13093 8616
rect 12952 8576 12958 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13228 8588 13461 8616
rect 13228 8576 13234 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14458 8616 14464 8628
rect 14415 8588 14464 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 17034 8616 17040 8628
rect 14608 8588 17040 8616
rect 14608 8576 14614 8588
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17310 8576 17316 8628
rect 17368 8576 17374 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 20165 8619 20223 8625
rect 18012 8588 20116 8616
rect 18012 8576 18018 8588
rect 10152 8548 10180 8576
rect 10318 8548 10324 8560
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 7926 8480 7932 8492
rect 7883 8452 7932 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7432 8384 7481 8412
rect 7432 8372 7438 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8588 8412 8616 8534
rect 10152 8520 10324 8548
rect 10318 8508 10324 8520
rect 10376 8548 10382 8560
rect 12176 8548 12204 8576
rect 13998 8548 14004 8560
rect 10376 8520 12204 8548
rect 12268 8520 14004 8548
rect 10376 8508 10382 8520
rect 12268 8492 12296 8520
rect 13998 8508 14004 8520
rect 14056 8548 14062 8560
rect 17494 8548 17500 8560
rect 14056 8520 16068 8548
rect 14056 8508 14062 8520
rect 9263 8483 9321 8489
rect 9263 8449 9275 8483
rect 9309 8480 9321 8483
rect 10134 8480 10140 8492
rect 9309 8452 10140 8480
rect 9309 8449 9321 8452
rect 9263 8443 9321 8449
rect 10134 8440 10140 8452
rect 10192 8480 10198 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 10192 8452 10241 8480
rect 10192 8440 10198 8452
rect 10229 8449 10241 8452
rect 10275 8480 10287 8483
rect 10502 8480 10508 8492
rect 10275 8452 10508 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10502 8440 10508 8452
rect 10560 8480 10566 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10560 8452 10609 8480
rect 10560 8440 10566 8452
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 12032 8452 12081 8480
rect 12032 8440 12038 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12250 8440 12256 8492
rect 12308 8440 12314 8492
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13262 8440 13268 8492
rect 13320 8440 13326 8492
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13722 8480 13728 8492
rect 13587 8452 13728 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 13906 8480 13912 8492
rect 13780 8452 13912 8480
rect 13780 8440 13786 8452
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14384 8489 14412 8520
rect 16040 8492 16068 8520
rect 17236 8520 17500 8548
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 8352 8384 8616 8412
rect 8352 8372 8358 8384
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 11900 8412 11928 8440
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11756 8384 12173 8412
rect 11756 8372 11762 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 13188 8412 13216 8440
rect 14108 8412 14136 8443
rect 13188 8384 14136 8412
rect 14292 8412 14320 8443
rect 15654 8440 15660 8492
rect 15712 8440 15718 8492
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 17236 8489 17264 8520
rect 17494 8508 17500 8520
rect 17552 8508 17558 8560
rect 17604 8548 17632 8576
rect 18138 8548 18144 8560
rect 17604 8520 18144 8548
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 18322 8508 18328 8560
rect 18380 8508 18386 8560
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 17368 8452 17417 8480
rect 17368 8440 17374 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17512 8480 17540 8508
rect 18340 8480 18368 8508
rect 17512 8452 18368 8480
rect 17405 8443 17463 8449
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 15672 8412 15700 8440
rect 14292 8384 15700 8412
rect 12345 8375 12403 8381
rect 12360 8344 12388 8375
rect 18046 8372 18052 8424
rect 18104 8372 18110 8424
rect 18322 8372 18328 8424
rect 18380 8372 18386 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18874 8412 18880 8424
rect 18555 8384 18880 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 19245 8415 19303 8421
rect 19245 8412 19257 8415
rect 19076 8384 19257 8412
rect 12526 8344 12532 8356
rect 11440 8316 12532 8344
rect 11440 8288 11468 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 17218 8344 17224 8356
rect 13688 8316 17224 8344
rect 13688 8304 13694 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18064 8344 18092 8372
rect 18782 8344 18788 8356
rect 18064 8316 18788 8344
rect 18782 8304 18788 8316
rect 18840 8344 18846 8356
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 18840 8316 18981 8344
rect 18840 8304 18846 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 18969 8307 19027 8313
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 11422 8276 11428 8288
rect 10008 8248 11428 8276
rect 10008 8236 10014 8248
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 11882 8236 11888 8288
rect 11940 8236 11946 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 13354 8276 13360 8288
rect 12124 8248 13360 8276
rect 12124 8236 12130 8248
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 17586 8276 17592 8288
rect 13504 8248 17592 8276
rect 13504 8236 13510 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18230 8236 18236 8288
rect 18288 8276 18294 8288
rect 19076 8276 19104 8384
rect 19245 8381 19257 8384
rect 19291 8381 19303 8415
rect 19245 8375 19303 8381
rect 19383 8415 19441 8421
rect 19383 8381 19395 8415
rect 19429 8412 19441 8415
rect 20088 8412 20116 8588
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20346 8616 20352 8628
rect 20211 8588 20352 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 23293 8619 23351 8625
rect 23293 8616 23305 8619
rect 22060 8588 23305 8616
rect 22060 8576 22066 8588
rect 23293 8585 23305 8588
rect 23339 8585 23351 8619
rect 23293 8579 23351 8585
rect 23382 8576 23388 8628
rect 23440 8576 23446 8628
rect 23658 8576 23664 8628
rect 23716 8616 23722 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23716 8588 24041 8616
rect 23716 8576 23722 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 24397 8619 24455 8625
rect 24397 8585 24409 8619
rect 24443 8616 24455 8619
rect 24946 8616 24952 8628
rect 24443 8588 24952 8616
rect 24443 8585 24455 8588
rect 24397 8579 24455 8585
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 26053 8619 26111 8625
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26878 8616 26884 8628
rect 26099 8588 26884 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26878 8576 26884 8588
rect 26936 8616 26942 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26936 8588 27353 8616
rect 26936 8576 26942 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27341 8579 27399 8585
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 28997 8619 29055 8625
rect 28997 8616 29009 8619
rect 28592 8588 29009 8616
rect 28592 8576 28598 8588
rect 28997 8585 29009 8588
rect 29043 8585 29055 8619
rect 28997 8579 29055 8585
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 29788 8588 30389 8616
rect 29788 8576 29794 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 30377 8579 30435 8585
rect 30650 8576 30656 8628
rect 30708 8616 30714 8628
rect 30708 8588 31892 8616
rect 30708 8576 30714 8588
rect 22462 8548 22468 8560
rect 21652 8520 22468 8548
rect 21652 8489 21680 8520
rect 22462 8508 22468 8520
rect 22520 8508 22526 8560
rect 23400 8548 23428 8576
rect 23400 8520 23980 8548
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8449 21695 8483
rect 21637 8443 21695 8449
rect 21910 8440 21916 8492
rect 21968 8440 21974 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8480 22155 8483
rect 23474 8480 23480 8492
rect 22143 8452 23480 8480
rect 22143 8449 22155 8452
rect 22097 8443 22155 8449
rect 23474 8440 23480 8452
rect 23532 8440 23538 8492
rect 23569 8483 23627 8489
rect 23569 8449 23581 8483
rect 23615 8449 23627 8483
rect 23569 8443 23627 8449
rect 19429 8384 20116 8412
rect 19429 8381 19441 8384
rect 19383 8375 19441 8381
rect 21358 8372 21364 8424
rect 21416 8372 21422 8424
rect 21928 8412 21956 8440
rect 22186 8412 22192 8424
rect 21928 8384 22192 8412
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 21545 8347 21603 8353
rect 21545 8313 21557 8347
rect 21591 8344 21603 8347
rect 22278 8344 22284 8356
rect 21591 8316 22284 8344
rect 21591 8313 21603 8316
rect 21545 8307 21603 8313
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 18288 8248 19104 8276
rect 18288 8236 18294 8248
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 20162 8276 20168 8288
rect 19576 8248 20168 8276
rect 19576 8236 19582 8248
rect 20162 8236 20168 8248
rect 20220 8236 20226 8288
rect 22094 8236 22100 8288
rect 22152 8236 22158 8288
rect 23584 8276 23612 8443
rect 23658 8440 23664 8492
rect 23716 8440 23722 8492
rect 23952 8489 23980 8520
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 23768 8344 23796 8443
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 28552 8489 28580 8576
rect 28626 8508 28632 8560
rect 28684 8548 28690 8560
rect 28684 8520 28856 8548
rect 28684 8508 28690 8520
rect 28828 8489 28856 8520
rect 24489 8483 24547 8489
rect 24489 8480 24501 8483
rect 24084 8452 24501 8480
rect 24084 8440 24090 8452
rect 24489 8449 24501 8452
rect 24535 8480 24547 8483
rect 27525 8483 27583 8489
rect 24535 8452 25360 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 25332 8424 25360 8452
rect 27525 8449 27537 8483
rect 27571 8480 27583 8483
rect 28537 8483 28595 8489
rect 27571 8452 28304 8480
rect 27571 8449 27583 8452
rect 27525 8443 27583 8449
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 25314 8372 25320 8424
rect 25372 8372 25378 8424
rect 26145 8415 26203 8421
rect 26145 8381 26157 8415
rect 26191 8381 26203 8415
rect 26145 8375 26203 8381
rect 26237 8415 26295 8421
rect 26237 8381 26249 8415
rect 26283 8412 26295 8415
rect 26602 8412 26608 8424
rect 26283 8384 26608 8412
rect 26283 8381 26295 8384
rect 26237 8375 26295 8381
rect 24946 8344 24952 8356
rect 23768 8316 24952 8344
rect 24946 8304 24952 8316
rect 25004 8304 25010 8356
rect 26160 8344 26188 8375
rect 26602 8372 26608 8384
rect 26660 8372 26666 8424
rect 27062 8372 27068 8424
rect 27120 8372 27126 8424
rect 27709 8415 27767 8421
rect 27709 8381 27721 8415
rect 27755 8412 27767 8415
rect 28166 8412 28172 8424
rect 27755 8384 28172 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 28166 8372 28172 8384
rect 28224 8372 28230 8424
rect 28276 8412 28304 8452
rect 28537 8449 28549 8483
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29104 8412 29132 8443
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 30190 8480 30196 8492
rect 29604 8452 30196 8480
rect 29604 8440 29610 8452
rect 30190 8440 30196 8452
rect 30248 8480 30254 8492
rect 30285 8483 30343 8489
rect 30285 8480 30297 8483
rect 30248 8452 30297 8480
rect 30248 8440 30254 8452
rect 30285 8449 30297 8452
rect 30331 8449 30343 8483
rect 30285 8443 30343 8449
rect 30374 8440 30380 8492
rect 30432 8480 30438 8492
rect 30760 8489 30788 8588
rect 30926 8508 30932 8560
rect 30984 8548 30990 8560
rect 31864 8548 31892 8588
rect 32214 8576 32220 8628
rect 32272 8576 32278 8628
rect 34146 8576 34152 8628
rect 34204 8576 34210 8628
rect 34514 8576 34520 8628
rect 34572 8576 34578 8628
rect 35434 8576 35440 8628
rect 35492 8616 35498 8628
rect 35529 8619 35587 8625
rect 35529 8616 35541 8619
rect 35492 8588 35541 8616
rect 35492 8576 35498 8588
rect 35529 8585 35541 8588
rect 35575 8585 35587 8619
rect 35529 8579 35587 8585
rect 37734 8576 37740 8628
rect 37792 8576 37798 8628
rect 41506 8576 41512 8628
rect 41564 8616 41570 8628
rect 42521 8619 42579 8625
rect 42521 8616 42533 8619
rect 41564 8588 42533 8616
rect 41564 8576 41570 8588
rect 42521 8585 42533 8588
rect 42567 8585 42579 8619
rect 42521 8579 42579 8585
rect 32232 8548 32260 8576
rect 30984 8520 31064 8548
rect 30984 8508 30990 8520
rect 31036 8489 31064 8520
rect 31864 8520 32260 8548
rect 30469 8483 30527 8489
rect 30469 8480 30481 8483
rect 30432 8452 30481 8480
rect 30432 8440 30438 8452
rect 30469 8449 30481 8452
rect 30515 8449 30527 8483
rect 30469 8443 30527 8449
rect 30745 8483 30803 8489
rect 30745 8449 30757 8483
rect 30791 8449 30803 8483
rect 30745 8443 30803 8449
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8480 31079 8483
rect 31202 8480 31208 8492
rect 31067 8452 31208 8480
rect 31067 8449 31079 8452
rect 31021 8443 31079 8449
rect 29178 8412 29184 8424
rect 28276 8384 28856 8412
rect 29104 8384 29184 8412
rect 26326 8344 26332 8356
rect 26160 8316 26332 8344
rect 26326 8304 26332 8316
rect 26384 8344 26390 8356
rect 27080 8344 27108 8372
rect 28828 8356 28856 8384
rect 29178 8372 29184 8384
rect 29236 8372 29242 8424
rect 30484 8412 30512 8443
rect 31202 8440 31208 8452
rect 31260 8440 31266 8492
rect 31294 8440 31300 8492
rect 31352 8484 31358 8492
rect 31481 8484 31539 8489
rect 31352 8483 31539 8484
rect 31352 8456 31493 8483
rect 31352 8440 31358 8456
rect 31481 8449 31493 8456
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31768 8483 31826 8489
rect 31768 8449 31780 8483
rect 31814 8480 31826 8483
rect 31864 8480 31892 8520
rect 31814 8452 31892 8480
rect 31814 8449 31826 8452
rect 31768 8443 31826 8449
rect 31938 8440 31944 8492
rect 31996 8480 32002 8492
rect 32125 8483 32183 8489
rect 32125 8480 32137 8483
rect 31996 8452 32137 8480
rect 31996 8440 32002 8452
rect 32125 8449 32137 8452
rect 32171 8449 32183 8483
rect 32232 8480 32260 8520
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 32232 8452 32321 8480
rect 32125 8443 32183 8449
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 33873 8483 33931 8489
rect 33873 8449 33885 8483
rect 33919 8449 33931 8483
rect 34164 8480 34192 8576
rect 34425 8551 34483 8557
rect 34425 8517 34437 8551
rect 34471 8548 34483 8551
rect 34532 8548 34560 8576
rect 37752 8548 37780 8576
rect 34471 8520 34560 8548
rect 35636 8520 37780 8548
rect 34471 8517 34483 8520
rect 34425 8511 34483 8517
rect 35636 8489 35664 8520
rect 43714 8508 43720 8560
rect 43772 8548 43778 8560
rect 43772 8520 44312 8548
rect 43772 8508 43778 8520
rect 34701 8483 34759 8489
rect 34701 8480 34713 8483
rect 34164 8452 34713 8480
rect 33873 8443 33931 8449
rect 34701 8449 34713 8452
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 35437 8483 35495 8489
rect 35437 8449 35449 8483
rect 35483 8449 35495 8483
rect 35437 8443 35495 8449
rect 35621 8483 35679 8489
rect 35621 8449 35633 8483
rect 35667 8449 35679 8483
rect 35621 8443 35679 8449
rect 35897 8483 35955 8489
rect 35897 8449 35909 8483
rect 35943 8449 35955 8483
rect 35897 8443 35955 8449
rect 30484 8384 30696 8412
rect 26384 8316 27108 8344
rect 26384 8304 26390 8316
rect 27154 8304 27160 8356
rect 27212 8344 27218 8356
rect 28261 8347 28319 8353
rect 28261 8344 28273 8347
rect 27212 8316 28273 8344
rect 27212 8304 27218 8316
rect 28261 8313 28273 8316
rect 28307 8313 28319 8347
rect 28261 8307 28319 8313
rect 28810 8304 28816 8356
rect 28868 8304 28874 8356
rect 30561 8347 30619 8353
rect 30561 8344 30573 8347
rect 28920 8316 30573 8344
rect 24578 8276 24584 8288
rect 23584 8248 24584 8276
rect 24578 8236 24584 8248
rect 24636 8236 24642 8288
rect 25682 8236 25688 8288
rect 25740 8236 25746 8288
rect 28721 8279 28779 8285
rect 28721 8245 28733 8279
rect 28767 8276 28779 8279
rect 28920 8276 28948 8316
rect 30561 8313 30573 8316
rect 30607 8313 30619 8347
rect 30668 8344 30696 8384
rect 30834 8372 30840 8424
rect 30892 8372 30898 8424
rect 30929 8415 30987 8421
rect 30929 8381 30941 8415
rect 30975 8412 30987 8415
rect 31110 8412 31116 8424
rect 30975 8384 31116 8412
rect 30975 8381 30987 8384
rect 30929 8375 30987 8381
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 33888 8412 33916 8443
rect 33965 8415 34023 8421
rect 33965 8412 33977 8415
rect 33888 8384 33977 8412
rect 33965 8381 33977 8384
rect 34011 8381 34023 8415
rect 35452 8412 35480 8443
rect 35526 8412 35532 8424
rect 35452 8384 35532 8412
rect 33965 8375 34023 8381
rect 35526 8372 35532 8384
rect 35584 8412 35590 8424
rect 35713 8415 35771 8421
rect 35713 8412 35725 8415
rect 35584 8384 35725 8412
rect 35584 8372 35590 8384
rect 35713 8381 35725 8384
rect 35759 8381 35771 8415
rect 35912 8412 35940 8443
rect 36078 8440 36084 8492
rect 36136 8440 36142 8492
rect 36909 8483 36967 8489
rect 36909 8480 36921 8483
rect 36740 8452 36921 8480
rect 36740 8412 36768 8452
rect 36909 8449 36921 8452
rect 36955 8449 36967 8483
rect 36909 8443 36967 8449
rect 37093 8483 37151 8489
rect 37093 8449 37105 8483
rect 37139 8480 37151 8483
rect 37277 8483 37335 8489
rect 37277 8480 37289 8483
rect 37139 8452 37289 8480
rect 37139 8449 37151 8452
rect 37093 8443 37151 8449
rect 37277 8449 37289 8452
rect 37323 8449 37335 8483
rect 37277 8443 37335 8449
rect 38010 8440 38016 8492
rect 38068 8440 38074 8492
rect 38194 8440 38200 8492
rect 38252 8440 38258 8492
rect 38289 8483 38347 8489
rect 38289 8449 38301 8483
rect 38335 8480 38347 8483
rect 38378 8480 38384 8492
rect 38335 8452 38384 8480
rect 38335 8449 38347 8452
rect 38289 8443 38347 8449
rect 38378 8440 38384 8452
rect 38436 8440 38442 8492
rect 44284 8489 44312 8520
rect 44269 8483 44327 8489
rect 42812 8452 42918 8480
rect 42812 8424 42840 8452
rect 44269 8449 44281 8483
rect 44315 8449 44327 8483
rect 44269 8443 44327 8449
rect 35912 8384 36768 8412
rect 35713 8375 35771 8381
rect 31205 8347 31263 8353
rect 31205 8344 31217 8347
rect 30668 8316 31217 8344
rect 30561 8307 30619 8313
rect 31205 8313 31217 8316
rect 31251 8313 31263 8347
rect 31205 8307 31263 8313
rect 31478 8304 31484 8356
rect 31536 8344 31542 8356
rect 32217 8347 32275 8353
rect 32217 8344 32229 8347
rect 31536 8316 32229 8344
rect 31536 8304 31542 8316
rect 32217 8313 32229 8316
rect 32263 8313 32275 8347
rect 32217 8307 32275 8313
rect 33226 8304 33232 8356
rect 33284 8344 33290 8356
rect 33689 8347 33747 8353
rect 33689 8344 33701 8347
rect 33284 8316 33701 8344
rect 33284 8304 33290 8316
rect 33689 8313 33701 8316
rect 33735 8313 33747 8347
rect 33689 8307 33747 8313
rect 34054 8304 34060 8356
rect 34112 8304 34118 8356
rect 34330 8304 34336 8356
rect 34388 8344 34394 8356
rect 34517 8347 34575 8353
rect 34517 8344 34529 8347
rect 34388 8316 34529 8344
rect 34388 8304 34394 8316
rect 34517 8313 34529 8316
rect 34563 8313 34575 8347
rect 36740 8344 36768 8384
rect 36817 8415 36875 8421
rect 36817 8381 36829 8415
rect 36863 8412 36875 8415
rect 37001 8415 37059 8421
rect 37001 8412 37013 8415
rect 36863 8384 37013 8412
rect 36863 8381 36875 8384
rect 36817 8375 36875 8381
rect 37001 8381 37013 8384
rect 37047 8381 37059 8415
rect 37001 8375 37059 8381
rect 37921 8415 37979 8421
rect 37921 8381 37933 8415
rect 37967 8381 37979 8415
rect 37921 8375 37979 8381
rect 37936 8344 37964 8375
rect 42794 8372 42800 8424
rect 42852 8372 42858 8424
rect 43990 8372 43996 8424
rect 44048 8372 44054 8424
rect 38013 8347 38071 8353
rect 38013 8344 38025 8347
rect 36740 8316 37320 8344
rect 37936 8316 38025 8344
rect 34517 8307 34575 8313
rect 28767 8248 28948 8276
rect 28767 8245 28779 8248
rect 28721 8239 28779 8245
rect 31386 8236 31392 8288
rect 31444 8276 31450 8288
rect 31570 8276 31576 8288
rect 31444 8248 31576 8276
rect 31444 8236 31450 8248
rect 31570 8236 31576 8248
rect 31628 8276 31634 8288
rect 31938 8276 31944 8288
rect 31628 8248 31944 8276
rect 31628 8236 31634 8248
rect 31938 8236 31944 8248
rect 31996 8236 32002 8288
rect 36170 8236 36176 8288
rect 36228 8236 36234 8288
rect 37292 8276 37320 8316
rect 38013 8313 38025 8316
rect 38059 8313 38071 8347
rect 38013 8307 38071 8313
rect 37918 8276 37924 8288
rect 37292 8248 37924 8276
rect 37918 8236 37924 8248
rect 37976 8236 37982 8288
rect 1104 8186 44620 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 44620 8186
rect 1104 8112 44620 8134
rect 6730 8032 6736 8084
rect 6788 8032 6794 8084
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 12250 8072 12256 8084
rect 11195 8044 12256 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 13262 8072 13268 8084
rect 12406 8044 13268 8072
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6748 7936 6776 8032
rect 10781 8007 10839 8013
rect 10781 7973 10793 8007
rect 10827 8004 10839 8007
rect 11054 8004 11060 8016
rect 10827 7976 11060 8004
rect 10827 7973 10839 7976
rect 10781 7967 10839 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 12406 8004 12434 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13446 8072 13452 8084
rect 13403 8044 13452 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 16301 8075 16359 8081
rect 15611 8044 16252 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 11348 7976 12434 8004
rect 6687 7908 6776 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 7098 7896 7104 7948
rect 7156 7896 7162 7948
rect 10152 7908 11008 7936
rect 10152 7880 10180 7908
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 7190 7868 7196 7880
rect 6779 7840 7196 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 10134 7828 10140 7880
rect 10192 7828 10198 7880
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 9950 7692 9956 7744
rect 10008 7692 10014 7744
rect 10336 7732 10364 7828
rect 10428 7800 10456 7831
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 10980 7877 11008 7908
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 10704 7800 10732 7828
rect 10428 7772 10732 7800
rect 10796 7800 10824 7831
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11072 7800 11100 7828
rect 10796 7772 11100 7800
rect 11348 7732 11376 7976
rect 15654 7964 15660 8016
rect 15712 8004 15718 8016
rect 16224 8004 16252 8044
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16390 8072 16396 8084
rect 16347 8044 16396 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 17773 8075 17831 8081
rect 17773 8041 17785 8075
rect 17819 8072 17831 8075
rect 18230 8072 18236 8084
rect 17819 8044 18236 8072
rect 17819 8041 17831 8044
rect 17773 8035 17831 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18380 8044 18613 8072
rect 18380 8032 18386 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18932 8044 19257 8072
rect 18932 8032 18938 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 19978 8032 19984 8084
rect 20036 8032 20042 8084
rect 20622 8032 20628 8084
rect 20680 8032 20686 8084
rect 21453 8075 21511 8081
rect 21453 8041 21465 8075
rect 21499 8072 21511 8075
rect 21542 8072 21548 8084
rect 21499 8044 21548 8072
rect 21499 8041 21511 8044
rect 21453 8035 21511 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 22278 8032 22284 8084
rect 22336 8032 22342 8084
rect 23474 8032 23480 8084
rect 23532 8032 23538 8084
rect 25866 8032 25872 8084
rect 25924 8032 25930 8084
rect 27706 8032 27712 8084
rect 27764 8072 27770 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 27764 8044 28089 8072
rect 27764 8032 27770 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 28258 8032 28264 8084
rect 28316 8072 28322 8084
rect 28810 8072 28816 8084
rect 28316 8044 28816 8072
rect 28316 8032 28322 8044
rect 28810 8032 28816 8044
rect 28868 8032 28874 8084
rect 31113 8075 31171 8081
rect 31113 8041 31125 8075
rect 31159 8041 31171 8075
rect 31113 8035 31171 8041
rect 19061 8007 19119 8013
rect 15712 7976 16160 8004
rect 16224 7976 19012 8004
rect 15712 7964 15718 7976
rect 11882 7896 11888 7948
rect 11940 7896 11946 7948
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7936 12035 7939
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12023 7908 12725 7936
rect 12023 7905 12035 7908
rect 11977 7899 12035 7905
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 14936 7908 15424 7936
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11550 7871 11608 7877
rect 11550 7868 11562 7871
rect 11480 7840 11562 7868
rect 11480 7828 11486 7840
rect 11550 7837 11562 7840
rect 11596 7837 11608 7871
rect 11900 7868 11928 7896
rect 14936 7880 14964 7908
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11900 7840 12081 7868
rect 11550 7831 11608 7837
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 12894 7868 12900 7880
rect 12851 7840 12900 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 12636 7800 12664 7831
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 14918 7828 14924 7880
rect 14976 7828 14982 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15396 7877 15424 7908
rect 15672 7877 15700 7964
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 16132 7936 16160 7976
rect 16853 7939 16911 7945
rect 16132 7908 16528 7936
rect 16500 7880 16528 7908
rect 16853 7905 16865 7939
rect 16899 7936 16911 7939
rect 17678 7936 17684 7948
rect 16899 7908 17684 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17678 7896 17684 7908
rect 17736 7936 17742 7948
rect 18509 7939 18567 7945
rect 17736 7908 18184 7936
rect 17736 7896 17742 7908
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 15068 7840 15117 7868
rect 15068 7828 15074 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7837 15255 7871
rect 15197 7831 15255 7837
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 13078 7800 13084 7812
rect 12636 7772 13084 7800
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 15212 7800 15240 7831
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 15286 7800 15292 7812
rect 13596 7772 15292 7800
rect 13596 7760 13602 7772
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 15396 7772 15761 7800
rect 10336 7704 11376 7732
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 11606 7692 11612 7744
rect 11664 7692 11670 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15396 7732 15424 7772
rect 15749 7769 15761 7772
rect 15795 7800 15807 7803
rect 16408 7800 16436 7831
rect 16482 7828 16488 7880
rect 16540 7868 16546 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 16540 7840 16681 7868
rect 16540 7828 16546 7840
rect 16669 7837 16681 7840
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 16960 7800 16988 7831
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 17092 7840 17141 7868
rect 17092 7828 17098 7840
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17644 7840 17969 7868
rect 17644 7828 17650 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18156 7868 18184 7908
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18598 7936 18604 7948
rect 18555 7908 18604 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18156 7840 18705 7868
rect 18049 7831 18107 7837
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18877 7871 18935 7877
rect 18877 7868 18889 7871
rect 18831 7840 18889 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18877 7837 18889 7840
rect 18923 7837 18935 7871
rect 18984 7868 19012 7976
rect 19061 7973 19073 8007
rect 19107 8004 19119 8007
rect 19996 8004 20024 8032
rect 19107 7976 20024 8004
rect 20640 8004 20668 8032
rect 20640 7976 22048 8004
rect 19107 7973 19119 7976
rect 19061 7967 19119 7973
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 19978 7936 19984 7948
rect 19935 7908 19984 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20254 7896 20260 7948
rect 20312 7896 20318 7948
rect 21910 7896 21916 7948
rect 21968 7896 21974 7948
rect 19061 7871 19119 7877
rect 19061 7868 19073 7871
rect 18984 7840 19073 7868
rect 18877 7831 18935 7837
rect 19061 7837 19073 7840
rect 19107 7868 19119 7871
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19107 7840 19625 7868
rect 19107 7837 19119 7840
rect 19061 7831 19119 7837
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 20272 7868 20300 7896
rect 19751 7840 20300 7868
rect 21637 7871 21695 7877
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 21637 7837 21649 7871
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 21818 7868 21824 7880
rect 21775 7840 21824 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 17773 7803 17831 7809
rect 17773 7800 17785 7803
rect 15795 7772 16436 7800
rect 16500 7772 16988 7800
rect 17052 7772 17785 7800
rect 15795 7769 15807 7772
rect 15749 7763 15807 7769
rect 15252 7704 15424 7732
rect 15252 7692 15258 7704
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 16500 7741 16528 7772
rect 17052 7744 17080 7772
rect 17773 7769 17785 7772
rect 17819 7769 17831 7803
rect 17773 7763 17831 7769
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15712 7704 15853 7732
rect 15712 7692 15718 7704
rect 15841 7701 15853 7704
rect 15887 7732 15899 7735
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 15887 7704 16497 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 16485 7701 16497 7704
rect 16531 7701 16543 7735
rect 16485 7695 16543 7701
rect 17034 7692 17040 7744
rect 17092 7692 17098 7744
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18064 7732 18092 7831
rect 18800 7800 18828 7831
rect 18524 7772 18828 7800
rect 21652 7800 21680 7831
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22020 7877 22048 7976
rect 30190 7964 30196 8016
rect 30248 8004 30254 8016
rect 30834 8004 30840 8016
rect 30248 7976 30840 8004
rect 30248 7964 30254 7976
rect 30834 7964 30840 7976
rect 30892 8004 30898 8016
rect 31128 8004 31156 8035
rect 31294 8032 31300 8084
rect 31352 8032 31358 8084
rect 31570 8032 31576 8084
rect 31628 8032 31634 8084
rect 38010 8032 38016 8084
rect 38068 8072 38074 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 38068 8044 38117 8072
rect 38068 8032 38074 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 38378 8032 38384 8084
rect 38436 8032 38442 8084
rect 43533 8075 43591 8081
rect 43533 8041 43545 8075
rect 43579 8072 43591 8075
rect 43990 8072 43996 8084
rect 43579 8044 43996 8072
rect 43579 8041 43591 8044
rect 43533 8035 43591 8041
rect 43990 8032 43996 8044
rect 44048 8032 44054 8084
rect 30892 7976 31156 8004
rect 30892 7964 30898 7976
rect 22186 7896 22192 7948
rect 22244 7936 22250 7948
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 22244 7908 22845 7936
rect 22244 7896 22250 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 22833 7899 22891 7905
rect 24121 7939 24179 7945
rect 24121 7905 24133 7939
rect 24167 7936 24179 7939
rect 24578 7936 24584 7948
rect 24167 7908 24584 7936
rect 24167 7905 24179 7908
rect 24121 7899 24179 7905
rect 24578 7896 24584 7908
rect 24636 7896 24642 7948
rect 24670 7896 24676 7948
rect 24728 7936 24734 7948
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24728 7908 24961 7936
rect 24728 7896 24734 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 26510 7896 26516 7948
rect 26568 7936 26574 7948
rect 27430 7936 27436 7948
rect 26568 7908 27436 7936
rect 26568 7896 26574 7908
rect 27430 7896 27436 7908
rect 27488 7896 27494 7948
rect 28902 7896 28908 7948
rect 28960 7936 28966 7948
rect 29178 7936 29184 7948
rect 28960 7908 29184 7936
rect 28960 7896 28966 7908
rect 29178 7896 29184 7908
rect 29236 7936 29242 7948
rect 29549 7939 29607 7945
rect 29549 7936 29561 7939
rect 29236 7908 29561 7936
rect 29236 7896 29242 7908
rect 29549 7905 29561 7908
rect 29595 7905 29607 7939
rect 29549 7899 29607 7905
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 31312 7936 31340 8032
rect 37918 7964 37924 8016
rect 37976 8004 37982 8016
rect 38197 8007 38255 8013
rect 38197 8004 38209 8007
rect 37976 7976 38209 8004
rect 37976 7964 37982 7976
rect 38197 7973 38209 7976
rect 38243 7973 38255 8007
rect 38197 7967 38255 7973
rect 31665 7939 31723 7945
rect 31665 7936 31677 7939
rect 31251 7908 31677 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 31665 7905 31677 7908
rect 31711 7905 31723 7939
rect 31665 7899 31723 7905
rect 37274 7896 37280 7948
rect 37332 7936 37338 7948
rect 38396 7936 38424 8032
rect 37332 7908 38424 7936
rect 37332 7896 37338 7908
rect 31757 7881 31815 7887
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7868 23903 7871
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 23891 7840 24777 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 24765 7837 24777 7840
rect 24811 7868 24823 7871
rect 25682 7868 25688 7880
rect 24811 7840 25688 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 26329 7871 26387 7877
rect 26329 7837 26341 7871
rect 26375 7868 26387 7871
rect 26375 7840 27752 7868
rect 26375 7837 26387 7840
rect 26329 7831 26387 7837
rect 22094 7800 22100 7812
rect 21652 7772 22100 7800
rect 18524 7744 18552 7772
rect 22094 7760 22100 7772
rect 22152 7760 22158 7812
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 22704 7772 24440 7800
rect 22704 7760 22710 7772
rect 17736 7704 18092 7732
rect 17736 7692 17742 7704
rect 18506 7692 18512 7744
rect 18564 7692 18570 7744
rect 22738 7692 22744 7744
rect 22796 7692 22802 7744
rect 23937 7735 23995 7741
rect 23937 7701 23949 7735
rect 23983 7732 23995 7735
rect 24302 7732 24308 7744
rect 23983 7704 24308 7732
rect 23983 7701 23995 7704
rect 23937 7695 23995 7701
rect 24302 7692 24308 7704
rect 24360 7692 24366 7744
rect 24412 7741 24440 7772
rect 24854 7760 24860 7812
rect 24912 7760 24918 7812
rect 26237 7803 26295 7809
rect 26237 7769 26249 7803
rect 26283 7800 26295 7803
rect 26283 7772 27568 7800
rect 26283 7769 26295 7772
rect 26237 7763 26295 7769
rect 27540 7744 27568 7772
rect 27724 7744 27752 7840
rect 29270 7828 29276 7880
rect 29328 7868 29334 7880
rect 29822 7868 29828 7880
rect 29328 7840 29828 7868
rect 29328 7828 29334 7840
rect 29822 7828 29828 7840
rect 29880 7828 29886 7880
rect 30009 7871 30067 7877
rect 30009 7837 30021 7871
rect 30055 7868 30067 7871
rect 30098 7868 30104 7880
rect 30055 7840 30104 7868
rect 30055 7837 30067 7840
rect 30009 7831 30067 7837
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 30190 7828 30196 7880
rect 30248 7868 30254 7880
rect 30285 7871 30343 7877
rect 30285 7868 30297 7871
rect 30248 7840 30297 7868
rect 30248 7828 30254 7840
rect 30285 7837 30297 7840
rect 30331 7868 30343 7871
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 30331 7840 31309 7868
rect 30331 7837 30343 7840
rect 30285 7831 30343 7837
rect 31297 7837 31309 7840
rect 31343 7868 31355 7871
rect 31478 7868 31484 7880
rect 31343 7840 31484 7868
rect 31343 7837 31355 7840
rect 31297 7831 31355 7837
rect 31478 7828 31484 7840
rect 31536 7828 31542 7880
rect 31757 7868 31769 7881
rect 31726 7847 31769 7868
rect 31803 7847 31815 7881
rect 31726 7841 31815 7847
rect 34517 7871 34575 7877
rect 31726 7840 31800 7841
rect 31726 7812 31754 7840
rect 34517 7837 34529 7871
rect 34563 7868 34575 7871
rect 37461 7871 37519 7877
rect 37461 7868 37473 7871
rect 34563 7840 35388 7868
rect 34563 7837 34575 7840
rect 34517 7831 34575 7837
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 29914 7800 29920 7812
rect 28500 7772 29920 7800
rect 28500 7760 28506 7772
rect 29914 7760 29920 7772
rect 29972 7800 29978 7812
rect 29972 7772 31432 7800
rect 31726 7772 31760 7812
rect 29972 7760 29978 7772
rect 24397 7735 24455 7741
rect 24397 7701 24409 7735
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 27522 7692 27528 7744
rect 27580 7692 27586 7744
rect 27706 7692 27712 7744
rect 27764 7692 27770 7744
rect 28245 7735 28303 7741
rect 28245 7701 28257 7735
rect 28291 7732 28303 7735
rect 28626 7732 28632 7744
rect 28291 7704 28632 7732
rect 28291 7701 28303 7704
rect 28245 7695 28303 7701
rect 28626 7692 28632 7704
rect 28684 7732 28690 7744
rect 29822 7732 29828 7744
rect 28684 7704 29828 7732
rect 28684 7692 28690 7704
rect 29822 7692 29828 7704
rect 29880 7732 29886 7744
rect 31404 7741 31432 7772
rect 31754 7760 31760 7772
rect 31812 7760 31818 7812
rect 33778 7760 33784 7812
rect 33836 7760 33842 7812
rect 34241 7803 34299 7809
rect 34241 7769 34253 7803
rect 34287 7800 34299 7803
rect 34330 7800 34336 7812
rect 34287 7772 34336 7800
rect 34287 7769 34299 7772
rect 34241 7763 34299 7769
rect 34330 7760 34336 7772
rect 34388 7760 34394 7812
rect 35360 7744 35388 7840
rect 37384 7840 37473 7868
rect 35894 7760 35900 7812
rect 35952 7800 35958 7812
rect 37093 7803 37151 7809
rect 37093 7800 37105 7803
rect 35952 7772 37105 7800
rect 35952 7760 35958 7772
rect 37093 7769 37105 7772
rect 37139 7769 37151 7803
rect 37093 7763 37151 7769
rect 37384 7800 37412 7840
rect 37461 7837 37473 7840
rect 37507 7837 37519 7871
rect 37461 7831 37519 7837
rect 43346 7828 43352 7880
rect 43404 7828 43410 7880
rect 38349 7803 38407 7809
rect 38349 7800 38361 7803
rect 37384 7772 38361 7800
rect 37384 7744 37412 7772
rect 38349 7769 38361 7772
rect 38395 7769 38407 7803
rect 38349 7763 38407 7769
rect 38562 7760 38568 7812
rect 38620 7760 38626 7812
rect 30929 7735 30987 7741
rect 30929 7732 30941 7735
rect 29880 7704 30941 7732
rect 29880 7692 29886 7704
rect 30929 7701 30941 7704
rect 30975 7701 30987 7735
rect 30929 7695 30987 7701
rect 31389 7735 31447 7741
rect 31389 7701 31401 7735
rect 31435 7701 31447 7735
rect 31389 7695 31447 7701
rect 32769 7735 32827 7741
rect 32769 7701 32781 7735
rect 32815 7732 32827 7735
rect 33410 7732 33416 7744
rect 32815 7704 33416 7732
rect 32815 7701 32827 7704
rect 32769 7695 32827 7701
rect 33410 7692 33416 7704
rect 33468 7692 33474 7744
rect 35342 7692 35348 7744
rect 35400 7732 35406 7744
rect 35805 7735 35863 7741
rect 35805 7732 35817 7735
rect 35400 7704 35817 7732
rect 35400 7692 35406 7704
rect 35805 7701 35817 7704
rect 35851 7732 35863 7735
rect 36998 7732 37004 7744
rect 35851 7704 37004 7732
rect 35851 7701 35863 7704
rect 35805 7695 35863 7701
rect 36998 7692 37004 7704
rect 37056 7692 37062 7744
rect 37366 7692 37372 7744
rect 37424 7692 37430 7744
rect 1104 7642 44620 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 44620 7642
rect 1104 7568 44620 7590
rect 7190 7488 7196 7540
rect 7248 7488 7254 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7742 7528 7748 7540
rect 7331 7500 7748 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 9950 7488 9956 7540
rect 10008 7488 10014 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7497 11023 7531
rect 10965 7491 11023 7497
rect 7208 7460 7236 7488
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 7208 7432 7389 7460
rect 7377 7429 7389 7432
rect 7423 7429 7435 7463
rect 7377 7423 7435 7429
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 7282 7392 7288 7404
rect 5859 7364 7288 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 7282 7352 7288 7364
rect 7340 7392 7346 7404
rect 9968 7392 9996 7488
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10980 7460 11008 7491
rect 11146 7488 11152 7540
rect 11204 7488 11210 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 11480 7500 12357 7528
rect 11480 7488 11486 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 12492 7500 12725 7528
rect 12492 7488 12498 7500
rect 12713 7497 12725 7500
rect 12759 7497 12771 7531
rect 12713 7491 12771 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 15378 7528 15384 7540
rect 13412 7500 15384 7528
rect 13412 7488 13418 7500
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 19061 7531 19119 7537
rect 19061 7497 19073 7531
rect 19107 7528 19119 7531
rect 19334 7528 19340 7540
rect 19107 7500 19340 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 21358 7488 21364 7540
rect 21416 7488 21422 7540
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 21876 7500 22569 7528
rect 21876 7488 21882 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23937 7531 23995 7537
rect 23937 7528 23949 7531
rect 22796 7500 23949 7528
rect 22796 7488 22802 7500
rect 23937 7497 23949 7500
rect 23983 7497 23995 7531
rect 23937 7491 23995 7497
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25004 7500 25176 7528
rect 25004 7488 25010 7500
rect 11606 7460 11612 7472
rect 10100 7432 10640 7460
rect 10980 7432 11612 7460
rect 10100 7420 10106 7432
rect 10612 7404 10640 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 15565 7463 15623 7469
rect 15565 7460 15577 7463
rect 12406 7432 15577 7460
rect 12406 7404 12434 7432
rect 15565 7429 15577 7432
rect 15611 7429 15623 7463
rect 15948 7460 15976 7488
rect 16025 7463 16083 7469
rect 16025 7460 16037 7463
rect 15948 7432 16037 7460
rect 15565 7423 15623 7429
rect 16025 7429 16037 7432
rect 16071 7460 16083 7463
rect 18138 7460 18144 7472
rect 16071 7432 18144 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 22373 7463 22431 7469
rect 22373 7429 22385 7463
rect 22419 7460 22431 7463
rect 22462 7460 22468 7472
rect 22419 7432 22468 7460
rect 22419 7429 22431 7432
rect 22373 7423 22431 7429
rect 22462 7420 22468 7432
rect 22520 7420 22526 7472
rect 24397 7463 24455 7469
rect 24397 7429 24409 7463
rect 24443 7460 24455 7463
rect 25038 7460 25044 7472
rect 24443 7432 25044 7460
rect 24443 7429 24455 7432
rect 24397 7423 24455 7429
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 25148 7460 25176 7500
rect 25314 7488 25320 7540
rect 25372 7488 25378 7540
rect 25777 7531 25835 7537
rect 25777 7497 25789 7531
rect 25823 7528 25835 7531
rect 26694 7528 26700 7540
rect 25823 7500 26700 7528
rect 25823 7497 25835 7500
rect 25777 7491 25835 7497
rect 26694 7488 26700 7500
rect 26752 7488 26758 7540
rect 26970 7488 26976 7540
rect 27028 7528 27034 7540
rect 27433 7531 27491 7537
rect 27433 7528 27445 7531
rect 27028 7500 27445 7528
rect 27028 7488 27034 7500
rect 27433 7497 27445 7500
rect 27479 7497 27491 7531
rect 27433 7491 27491 7497
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28077 7531 28135 7537
rect 28077 7528 28089 7531
rect 27948 7500 28089 7528
rect 27948 7488 27954 7500
rect 28077 7497 28089 7500
rect 28123 7497 28135 7531
rect 28077 7491 28135 7497
rect 28258 7488 28264 7540
rect 28316 7488 28322 7540
rect 28902 7488 28908 7540
rect 28960 7488 28966 7540
rect 29270 7488 29276 7540
rect 29328 7488 29334 7540
rect 29641 7531 29699 7537
rect 29641 7528 29653 7531
rect 29472 7500 29653 7528
rect 26237 7463 26295 7469
rect 26237 7460 26249 7463
rect 25148 7432 26249 7460
rect 26237 7429 26249 7432
rect 26283 7429 26295 7463
rect 27154 7460 27160 7472
rect 26237 7423 26295 7429
rect 26436 7432 27160 7460
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 7340 7364 9674 7392
rect 9968 7364 10517 7392
rect 7340 7352 7346 7364
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6730 7324 6736 7336
rect 5951 7296 6736 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7466 7284 7472 7336
rect 7524 7284 7530 7336
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 8202 7256 8208 7268
rect 6227 7228 8208 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 8202 7216 8208 7228
rect 8260 7216 8266 7268
rect 9646 7256 9674 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 10928 7364 11069 7392
rect 10928 7352 10934 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11238 7352 11244 7404
rect 11296 7352 11302 7404
rect 12342 7392 12348 7404
rect 11348 7364 12348 7392
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 11348 7324 11376 7364
rect 12342 7352 12348 7364
rect 12400 7364 12434 7404
rect 12400 7352 12406 7364
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 14936 7364 15393 7392
rect 10827 7296 11376 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 10502 7256 10508 7268
rect 9646 7228 10508 7256
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 10704 7256 10732 7287
rect 12158 7284 12164 7336
rect 12216 7284 12222 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12894 7324 12900 7336
rect 12299 7296 12900 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 11054 7256 11060 7268
rect 10704 7228 11060 7256
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11790 7216 11796 7268
rect 11848 7256 11854 7268
rect 13170 7256 13176 7268
rect 11848 7228 13176 7256
rect 11848 7216 11854 7228
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 13630 7216 13636 7268
rect 13688 7256 13694 7268
rect 14200 7256 14228 7352
rect 14936 7336 14964 7364
rect 15381 7361 15393 7364
rect 15427 7392 15439 7395
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15427 7364 15669 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 15979 7364 16068 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16040 7336 16068 7364
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18012 7364 18613 7392
rect 18012 7352 18018 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18690 7352 18696 7404
rect 18748 7352 18754 7404
rect 18782 7352 18788 7404
rect 18840 7392 18846 7404
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18840 7364 18889 7392
rect 18840 7352 18846 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 20806 7352 20812 7404
rect 20864 7392 20870 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20864 7364 21005 7392
rect 20864 7352 20870 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 14918 7284 14924 7336
rect 14976 7284 14982 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 14642 7256 14648 7268
rect 13688 7228 14648 7256
rect 13688 7216 13694 7228
rect 14642 7216 14648 7228
rect 14700 7256 14706 7268
rect 15212 7256 15240 7287
rect 16022 7284 16028 7336
rect 16080 7284 16086 7336
rect 21192 7324 21220 7355
rect 22830 7352 22836 7404
rect 22888 7392 22894 7404
rect 22888 7364 22932 7392
rect 22888 7352 22894 7364
rect 24302 7352 24308 7404
rect 24360 7352 24366 7404
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 24857 7395 24915 7401
rect 24857 7392 24869 7395
rect 24728 7364 24869 7392
rect 24728 7352 24734 7364
rect 24857 7361 24869 7364
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 25682 7352 25688 7404
rect 25740 7352 25746 7404
rect 26436 7401 26464 7432
rect 27154 7420 27160 7432
rect 27212 7420 27218 7472
rect 26421 7395 26479 7401
rect 26421 7361 26433 7395
rect 26467 7361 26479 7395
rect 26421 7355 26479 7361
rect 26510 7352 26516 7404
rect 26568 7352 26574 7404
rect 26697 7395 26755 7401
rect 26697 7392 26709 7395
rect 26687 7361 26709 7392
rect 26743 7361 26755 7395
rect 26687 7355 26755 7361
rect 21450 7324 21456 7336
rect 21192 7296 21456 7324
rect 21450 7284 21456 7296
rect 21508 7324 21514 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 21508 7296 22569 7324
rect 21508 7284 21514 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 14700 7228 15240 7256
rect 14700 7216 14706 7228
rect 22186 7216 22192 7268
rect 22244 7216 22250 7268
rect 24320 7256 24348 7352
rect 24578 7284 24584 7336
rect 24636 7284 24642 7336
rect 25866 7284 25872 7336
rect 25924 7284 25930 7336
rect 26687 7256 26715 7355
rect 26786 7352 26792 7404
rect 26844 7352 26850 7404
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 27706 7392 27712 7404
rect 27387 7364 27712 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 28169 7395 28227 7401
rect 28169 7361 28181 7395
rect 28215 7392 28227 7395
rect 28276 7392 28304 7488
rect 28613 7463 28671 7469
rect 28613 7429 28625 7463
rect 28659 7460 28671 7463
rect 28718 7460 28724 7472
rect 28659 7432 28724 7460
rect 28659 7429 28671 7432
rect 28613 7423 28671 7429
rect 28718 7420 28724 7432
rect 28776 7420 28782 7472
rect 28813 7463 28871 7469
rect 28813 7429 28825 7463
rect 28859 7460 28871 7463
rect 28920 7460 28948 7488
rect 29288 7460 29316 7488
rect 29472 7472 29500 7500
rect 29641 7497 29653 7500
rect 29687 7497 29699 7531
rect 29641 7491 29699 7497
rect 30098 7488 30104 7540
rect 30156 7528 30162 7540
rect 30156 7500 31248 7528
rect 30156 7488 30162 7500
rect 28859 7432 28948 7460
rect 29104 7432 29316 7460
rect 28859 7429 28871 7432
rect 28813 7423 28871 7429
rect 28215 7364 28304 7392
rect 28828 7392 28856 7423
rect 29104 7401 29132 7432
rect 29454 7420 29460 7472
rect 29512 7420 29518 7472
rect 30190 7460 30196 7472
rect 29564 7432 30196 7460
rect 28893 7395 28951 7401
rect 28893 7392 28905 7395
rect 28828 7364 28905 7392
rect 28215 7361 28227 7364
rect 28169 7355 28227 7361
rect 28893 7361 28905 7364
rect 28939 7361 28951 7395
rect 28893 7355 28951 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29181 7395 29239 7401
rect 29181 7361 29193 7395
rect 29227 7361 29239 7395
rect 29181 7355 29239 7361
rect 29319 7395 29377 7401
rect 29319 7361 29331 7395
rect 29365 7392 29377 7395
rect 29564 7392 29592 7432
rect 30190 7420 30196 7432
rect 30248 7420 30254 7472
rect 31220 7469 31248 7500
rect 33134 7488 33140 7540
rect 33192 7488 33198 7540
rect 33778 7488 33784 7540
rect 33836 7528 33842 7540
rect 35986 7528 35992 7540
rect 33836 7500 35992 7528
rect 33836 7488 33842 7500
rect 35986 7488 35992 7500
rect 36044 7528 36050 7540
rect 37093 7531 37151 7537
rect 36044 7500 36952 7528
rect 36044 7488 36050 7500
rect 31205 7463 31263 7469
rect 31205 7429 31217 7463
rect 31251 7429 31263 7463
rect 31205 7423 31263 7429
rect 31389 7463 31447 7469
rect 31389 7429 31401 7463
rect 31435 7460 31447 7463
rect 31754 7460 31760 7472
rect 31435 7432 31760 7460
rect 31435 7429 31447 7432
rect 31389 7423 31447 7429
rect 31754 7420 31760 7432
rect 31812 7420 31818 7472
rect 31846 7420 31852 7472
rect 31904 7460 31910 7472
rect 34609 7463 34667 7469
rect 34609 7460 34621 7463
rect 31904 7432 34621 7460
rect 31904 7420 31910 7432
rect 34609 7429 34621 7432
rect 34655 7460 34667 7463
rect 35894 7460 35900 7472
rect 34655 7432 35900 7460
rect 34655 7429 34667 7432
rect 34609 7423 34667 7429
rect 35894 7420 35900 7432
rect 35952 7420 35958 7472
rect 36004 7460 36032 7488
rect 36924 7460 36952 7500
rect 37093 7497 37105 7531
rect 37139 7528 37151 7531
rect 37366 7528 37372 7540
rect 37139 7500 37372 7528
rect 37139 7497 37151 7500
rect 37093 7491 37151 7497
rect 37366 7488 37372 7500
rect 37424 7488 37430 7540
rect 37458 7488 37464 7540
rect 37516 7528 37522 7540
rect 38562 7528 38568 7540
rect 37516 7500 38568 7528
rect 37516 7488 37522 7500
rect 38562 7488 38568 7500
rect 38620 7488 38626 7540
rect 42794 7528 42800 7540
rect 41386 7500 42800 7528
rect 36004 7432 36110 7460
rect 36924 7446 37766 7460
rect 36924 7432 37780 7446
rect 29365 7364 29592 7392
rect 29365 7361 29377 7364
rect 29319 7355 29377 7361
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 27488 7296 27537 7324
rect 27488 7284 27494 7296
rect 27525 7293 27537 7296
rect 27571 7324 27583 7327
rect 27816 7324 27844 7355
rect 27571 7296 27844 7324
rect 27985 7327 28043 7333
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 27985 7293 27997 7327
rect 28031 7293 28043 7327
rect 27985 7287 28043 7293
rect 27801 7259 27859 7265
rect 27801 7256 27813 7259
rect 24320 7228 26372 7256
rect 26687 7228 27813 7256
rect 6914 7148 6920 7200
rect 6972 7148 6978 7200
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 11422 7188 11428 7200
rect 10744 7160 11428 7188
rect 10744 7148 10750 7160
rect 11422 7148 11428 7160
rect 11480 7188 11486 7200
rect 19334 7188 19340 7200
rect 11480 7160 19340 7188
rect 11480 7148 11486 7160
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 22741 7191 22799 7197
rect 22741 7157 22753 7191
rect 22787 7188 22799 7191
rect 23474 7188 23480 7200
rect 22787 7160 23480 7188
rect 22787 7157 22799 7160
rect 22741 7151 22799 7157
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 25133 7191 25191 7197
rect 25133 7157 25145 7191
rect 25179 7188 25191 7191
rect 25314 7188 25320 7200
rect 25179 7160 25320 7188
rect 25179 7157 25191 7160
rect 25133 7151 25191 7157
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 25590 7148 25596 7200
rect 25648 7188 25654 7200
rect 25866 7188 25872 7200
rect 25648 7160 25872 7188
rect 25648 7148 25654 7160
rect 25866 7148 25872 7160
rect 25924 7148 25930 7200
rect 26344 7188 26372 7228
rect 27801 7225 27813 7228
rect 27847 7225 27859 7259
rect 28000 7256 28028 7287
rect 28994 7256 29000 7268
rect 28000 7228 29000 7256
rect 27801 7219 27859 7225
rect 28994 7216 29000 7228
rect 29052 7216 29058 7268
rect 29104 7200 29132 7355
rect 29196 7324 29224 7355
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 29914 7352 29920 7404
rect 29972 7392 29978 7404
rect 30101 7395 30159 7401
rect 29972 7364 30017 7392
rect 29972 7352 29978 7364
rect 30101 7361 30113 7395
rect 30147 7392 30159 7395
rect 30929 7395 30987 7401
rect 30929 7392 30941 7395
rect 30147 7364 30941 7392
rect 30147 7361 30159 7364
rect 30101 7355 30159 7361
rect 30929 7361 30941 7364
rect 30975 7392 30987 7395
rect 31018 7392 31024 7404
rect 30975 7364 31024 7392
rect 30975 7361 30987 7364
rect 30929 7355 30987 7361
rect 31018 7352 31024 7364
rect 31076 7352 31082 7404
rect 29454 7324 29460 7336
rect 29196 7296 29460 7324
rect 29454 7284 29460 7296
rect 29512 7324 29518 7336
rect 29656 7324 29684 7352
rect 29512 7296 29684 7324
rect 29512 7284 29518 7296
rect 29178 7216 29184 7268
rect 29236 7256 29242 7268
rect 29546 7256 29552 7268
rect 29236 7228 29552 7256
rect 29236 7216 29242 7228
rect 29546 7216 29552 7228
rect 29604 7216 29610 7268
rect 29656 7256 29684 7296
rect 29822 7284 29828 7336
rect 29880 7284 29886 7336
rect 30009 7327 30067 7333
rect 30009 7293 30021 7327
rect 30055 7293 30067 7327
rect 30009 7287 30067 7293
rect 30024 7256 30052 7287
rect 30742 7284 30748 7336
rect 30800 7324 30806 7336
rect 30837 7327 30895 7333
rect 30837 7324 30849 7327
rect 30800 7296 30849 7324
rect 30800 7284 30806 7296
rect 30837 7293 30849 7296
rect 30883 7293 30895 7327
rect 30837 7287 30895 7293
rect 31110 7284 31116 7336
rect 31168 7324 31174 7336
rect 31570 7324 31576 7336
rect 31168 7296 31576 7324
rect 31168 7284 31174 7296
rect 31570 7284 31576 7296
rect 31628 7284 31634 7336
rect 35342 7284 35348 7336
rect 35400 7284 35406 7336
rect 35621 7327 35679 7333
rect 35621 7293 35633 7327
rect 35667 7324 35679 7327
rect 36170 7324 36176 7336
rect 35667 7296 36176 7324
rect 35667 7293 35679 7296
rect 35621 7287 35679 7293
rect 36170 7284 36176 7296
rect 36228 7284 36234 7336
rect 37752 7324 37780 7432
rect 38470 7420 38476 7472
rect 38528 7460 38534 7472
rect 41386 7460 41414 7500
rect 42794 7488 42800 7500
rect 42852 7488 42858 7540
rect 43346 7488 43352 7540
rect 43404 7488 43410 7540
rect 38528 7432 41414 7460
rect 38528 7420 38534 7432
rect 43806 7420 43812 7472
rect 43864 7420 43870 7472
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7392 39267 7395
rect 43714 7392 43720 7404
rect 39255 7364 43720 7392
rect 39255 7361 39267 7364
rect 39209 7355 39267 7361
rect 43714 7352 43720 7364
rect 43772 7352 43778 7404
rect 44082 7352 44088 7404
rect 44140 7392 44146 7404
rect 44269 7395 44327 7401
rect 44269 7392 44281 7395
rect 44140 7364 44281 7392
rect 44140 7352 44146 7364
rect 44269 7361 44281 7364
rect 44315 7361 44327 7395
rect 44269 7355 44327 7361
rect 38470 7324 38476 7336
rect 37752 7296 38476 7324
rect 38470 7284 38476 7296
rect 38528 7284 38534 7336
rect 38930 7284 38936 7336
rect 38988 7284 38994 7336
rect 30098 7256 30104 7268
rect 29656 7228 30104 7256
rect 30098 7216 30104 7228
rect 30156 7216 30162 7268
rect 43533 7259 43591 7265
rect 30484 7228 30788 7256
rect 30484 7200 30512 7228
rect 26973 7191 27031 7197
rect 26973 7188 26985 7191
rect 26344 7160 26985 7188
rect 26973 7157 26985 7160
rect 27019 7157 27031 7191
rect 26973 7151 27031 7157
rect 27062 7148 27068 7200
rect 27120 7188 27126 7200
rect 28445 7191 28503 7197
rect 28445 7188 28457 7191
rect 27120 7160 28457 7188
rect 27120 7148 27126 7160
rect 28445 7157 28457 7160
rect 28491 7157 28503 7191
rect 28445 7151 28503 7157
rect 28629 7191 28687 7197
rect 28629 7157 28641 7191
rect 28675 7188 28687 7191
rect 29086 7188 29092 7200
rect 28675 7160 29092 7188
rect 28675 7157 28687 7160
rect 28629 7151 28687 7157
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 30466 7148 30472 7200
rect 30524 7148 30530 7200
rect 30558 7148 30564 7200
rect 30616 7148 30622 7200
rect 30760 7197 30788 7228
rect 43533 7225 43545 7259
rect 43579 7256 43591 7259
rect 44085 7259 44143 7265
rect 44085 7256 44097 7259
rect 43579 7228 44097 7256
rect 43579 7225 43591 7228
rect 43533 7219 43591 7225
rect 44085 7225 44097 7228
rect 44131 7225 44143 7259
rect 44085 7219 44143 7225
rect 30745 7191 30803 7197
rect 30745 7157 30757 7191
rect 30791 7157 30803 7191
rect 30745 7151 30803 7157
rect 30834 7148 30840 7200
rect 30892 7188 30898 7200
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 30892 7160 31033 7188
rect 30892 7148 30898 7160
rect 31021 7157 31033 7160
rect 31067 7188 31079 7191
rect 31478 7188 31484 7200
rect 31067 7160 31484 7188
rect 31067 7157 31079 7160
rect 31021 7151 31079 7157
rect 31478 7148 31484 7160
rect 31536 7148 31542 7200
rect 1104 7098 44620 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 44620 7098
rect 1104 7024 44620 7046
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 10965 6987 11023 6993
rect 10965 6984 10977 6987
rect 10928 6956 10977 6984
rect 10928 6944 10934 6956
rect 10965 6953 10977 6956
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 11296 6956 11437 6984
rect 11296 6944 11302 6956
rect 11425 6953 11437 6956
rect 11471 6984 11483 6987
rect 11471 6956 12480 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 2225 6919 2283 6925
rect 2225 6916 2237 6919
rect 2148 6888 2237 6916
rect 1946 6808 1952 6860
rect 2004 6808 2010 6860
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2148 6848 2176 6888
rect 2225 6885 2237 6888
rect 2271 6885 2283 6919
rect 2225 6879 2283 6885
rect 7009 6919 7067 6925
rect 7009 6885 7021 6919
rect 7055 6885 7067 6919
rect 7009 6879 7067 6885
rect 2096 6820 2176 6848
rect 2409 6851 2467 6857
rect 2096 6808 2102 6820
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2455 6820 2774 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2746 6780 2774 6820
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2746 6752 2973 6780
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7024 6780 7052 6879
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7524 6820 7573 6848
rect 7524 6808 7530 6820
rect 7561 6817 7573 6820
rect 7607 6848 7619 6851
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 7607 6820 8401 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8389 6817 8401 6820
rect 8435 6817 8447 6851
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 8389 6811 8447 6817
rect 10244 6820 11345 6848
rect 10244 6792 10272 6820
rect 11333 6817 11345 6820
rect 11379 6817 11391 6851
rect 12452 6848 12480 6956
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 13872 6956 14749 6984
rect 13872 6944 13878 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 14737 6947 14795 6953
rect 14918 6944 14924 6996
rect 14976 6944 14982 6996
rect 18049 6987 18107 6993
rect 18049 6953 18061 6987
rect 18095 6984 18107 6987
rect 18095 6956 18276 6984
rect 18095 6953 18107 6956
rect 18049 6947 18107 6953
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 15010 6916 15016 6928
rect 12584 6888 15016 6916
rect 12584 6876 12590 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6885 18199 6919
rect 18141 6879 18199 6885
rect 11333 6811 11391 6817
rect 11624 6820 12112 6848
rect 12452 6820 13768 6848
rect 6779 6752 7052 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 7156 6752 7389 6780
rect 7156 6740 7162 6752
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 10962 6780 10968 6792
rect 10919 6752 10968 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 7282 6672 7288 6724
rect 7340 6712 7346 6724
rect 7469 6715 7527 6721
rect 7469 6712 7481 6715
rect 7340 6684 7481 6712
rect 7340 6672 7346 6684
rect 7469 6681 7481 6684
rect 7515 6681 7527 6715
rect 7469 6675 7527 6681
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 9766 6712 9772 6724
rect 8343 6684 9772 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 9766 6672 9772 6684
rect 9824 6712 9830 6724
rect 10686 6712 10692 6724
rect 9824 6684 10692 6712
rect 9824 6672 9830 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 11348 6712 11376 6811
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 11624 6789 11652 6820
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11756 6752 11805 6780
rect 11756 6740 11762 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 12084 6780 12112 6820
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12084 6752 12725 6780
rect 11977 6743 12035 6749
rect 12713 6749 12725 6752
rect 12759 6780 12771 6783
rect 13740 6780 13768 6820
rect 15948 6820 17816 6848
rect 15948 6792 15976 6820
rect 12759 6752 13676 6780
rect 13740 6752 14412 6780
rect 12759 6749 12771 6752
rect 12713 6743 12771 6749
rect 11882 6712 11888 6724
rect 11348 6684 11888 6712
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 11992 6712 12020 6743
rect 11992 6684 12112 6712
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7650 6644 7656 6656
rect 6963 6616 7656 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7834 6604 7840 6656
rect 7892 6604 7898 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 12084 6644 12112 6684
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 12526 6672 12532 6724
rect 12584 6672 12590 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 12728 6684 13369 6712
rect 12544 6644 12572 6672
rect 12728 6656 12756 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13648 6712 13676 6752
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 13648 6684 13737 6712
rect 13357 6675 13415 6681
rect 13725 6681 13737 6684
rect 13771 6712 13783 6715
rect 13998 6712 14004 6724
rect 13771 6684 14004 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14384 6712 14412 6752
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14568 6712 14596 6743
rect 14826 6740 14832 6792
rect 14884 6740 14890 6792
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 15194 6780 15200 6792
rect 15059 6752 15200 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 16080 6752 16129 6780
rect 16080 6740 16086 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16390 6780 16396 6792
rect 16347 6752 16396 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 17788 6789 17816 6820
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18156 6780 18184 6879
rect 18248 6848 18276 6956
rect 25038 6944 25044 6996
rect 25096 6944 25102 6996
rect 26694 6944 26700 6996
rect 26752 6984 26758 6996
rect 26752 6956 27292 6984
rect 26752 6944 26758 6956
rect 18874 6876 18880 6928
rect 18932 6916 18938 6928
rect 20070 6916 20076 6928
rect 18932 6888 20076 6916
rect 18932 6876 18938 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 27264 6916 27292 6956
rect 27706 6944 27712 6996
rect 27764 6984 27770 6996
rect 29549 6987 29607 6993
rect 29549 6984 29561 6987
rect 27764 6956 29561 6984
rect 27764 6944 27770 6956
rect 29549 6953 29561 6956
rect 29595 6953 29607 6987
rect 29549 6947 29607 6953
rect 29733 6987 29791 6993
rect 29733 6953 29745 6987
rect 29779 6984 29791 6987
rect 30374 6984 30380 6996
rect 29779 6956 30380 6984
rect 29779 6953 29791 6956
rect 29733 6947 29791 6953
rect 30374 6944 30380 6956
rect 30432 6944 30438 6996
rect 30558 6944 30564 6996
rect 30616 6944 30622 6996
rect 30760 6956 30972 6984
rect 30576 6916 30604 6944
rect 25516 6888 25728 6916
rect 19242 6848 19248 6860
rect 18248 6820 19248 6848
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 24578 6808 24584 6860
rect 24636 6848 24642 6860
rect 25516 6848 25544 6888
rect 24636 6820 25544 6848
rect 24636 6808 24642 6820
rect 25590 6808 25596 6860
rect 25648 6808 25654 6860
rect 25700 6848 25728 6888
rect 26988 6888 27200 6916
rect 27264 6888 30604 6916
rect 26694 6857 26700 6860
rect 26513 6851 26571 6857
rect 26513 6848 26525 6851
rect 25700 6820 26525 6848
rect 26513 6817 26525 6820
rect 26559 6817 26571 6851
rect 26513 6811 26571 6817
rect 26672 6851 26700 6857
rect 26672 6817 26684 6851
rect 26672 6811 26700 6817
rect 26694 6808 26700 6811
rect 26752 6808 26758 6860
rect 26789 6851 26847 6857
rect 26789 6817 26801 6851
rect 26835 6848 26847 6851
rect 26988 6848 27016 6888
rect 27172 6860 27200 6888
rect 26835 6820 27016 6848
rect 26835 6817 26847 6820
rect 26789 6811 26847 6817
rect 27062 6808 27068 6860
rect 27120 6808 27126 6860
rect 27154 6808 27160 6860
rect 27212 6808 27218 6860
rect 27522 6808 27528 6860
rect 27580 6848 27586 6860
rect 28169 6851 28227 6857
rect 28169 6848 28181 6851
rect 27580 6820 28181 6848
rect 27580 6808 27586 6820
rect 28169 6817 28181 6820
rect 28215 6817 28227 6851
rect 28810 6848 28816 6860
rect 28169 6811 28227 6817
rect 28260 6820 28816 6848
rect 18095 6752 18184 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18288 6752 18429 6780
rect 18288 6740 18294 6752
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 23492 6780 23520 6808
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 23492 6752 25881 6780
rect 18417 6743 18475 6749
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 17954 6712 17960 6724
rect 14384 6684 17960 6712
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 18141 6715 18199 6721
rect 18141 6681 18153 6715
rect 18187 6681 18199 6715
rect 18141 6675 18199 6681
rect 11296 6616 12572 6644
rect 11296 6604 11302 6616
rect 12710 6604 12716 6656
rect 12768 6604 12774 6656
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13078 6644 13084 6656
rect 12943 6616 13084 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 15838 6644 15844 6656
rect 15344 6616 15844 6644
rect 15344 6604 15350 6616
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16209 6647 16267 6653
rect 16209 6644 16221 6647
rect 15988 6616 16221 6644
rect 15988 6604 15994 6616
rect 16209 6613 16221 6616
rect 16255 6613 16267 6647
rect 16209 6607 16267 6613
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17865 6647 17923 6653
rect 17865 6644 17877 6647
rect 17276 6616 17877 6644
rect 17276 6604 17282 6616
rect 17865 6613 17877 6616
rect 17911 6613 17923 6647
rect 17865 6607 17923 6613
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18156 6644 18184 6675
rect 18322 6672 18328 6724
rect 18380 6672 18386 6724
rect 25409 6715 25467 6721
rect 25409 6681 25421 6715
rect 25455 6712 25467 6715
rect 25455 6684 26096 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 18598 6644 18604 6656
rect 18104 6616 18604 6644
rect 18104 6604 18110 6616
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 25501 6647 25559 6653
rect 25501 6613 25513 6647
rect 25547 6644 25559 6647
rect 25682 6644 25688 6656
rect 25547 6616 25688 6644
rect 25547 6613 25559 6616
rect 25501 6607 25559 6613
rect 25682 6604 25688 6616
rect 25740 6604 25746 6656
rect 26068 6644 26096 6684
rect 27540 6644 27568 6808
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6780 27767 6783
rect 27798 6780 27804 6792
rect 27755 6752 27804 6780
rect 27755 6749 27767 6752
rect 27709 6743 27767 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 27890 6740 27896 6792
rect 27948 6740 27954 6792
rect 28077 6783 28135 6789
rect 28077 6749 28089 6783
rect 28123 6780 28135 6783
rect 28260 6780 28288 6820
rect 28810 6808 28816 6820
rect 28868 6808 28874 6860
rect 30469 6851 30527 6857
rect 28920 6820 30236 6848
rect 28920 6792 28948 6820
rect 28123 6752 28288 6780
rect 28353 6783 28411 6789
rect 28123 6749 28135 6752
rect 28077 6743 28135 6749
rect 28353 6749 28365 6783
rect 28399 6780 28411 6783
rect 28442 6780 28448 6792
rect 28399 6752 28448 6780
rect 28399 6749 28411 6752
rect 28353 6743 28411 6749
rect 28442 6740 28448 6752
rect 28500 6740 28506 6792
rect 28629 6783 28687 6789
rect 28629 6749 28641 6783
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 26068 6616 27568 6644
rect 27908 6644 27936 6740
rect 28644 6712 28672 6743
rect 28902 6740 28908 6792
rect 28960 6740 28966 6792
rect 28994 6740 29000 6792
rect 29052 6780 29058 6792
rect 29052 6752 30052 6780
rect 29052 6740 29058 6752
rect 29454 6712 29460 6724
rect 28644 6684 29460 6712
rect 29454 6672 29460 6684
rect 29512 6672 29518 6724
rect 29546 6672 29552 6724
rect 29604 6712 29610 6724
rect 29917 6715 29975 6721
rect 29917 6712 29929 6715
rect 29604 6684 29929 6712
rect 29604 6672 29610 6684
rect 29917 6681 29929 6684
rect 29963 6681 29975 6715
rect 30024 6712 30052 6752
rect 30098 6740 30104 6792
rect 30156 6740 30162 6792
rect 30208 6780 30236 6820
rect 30469 6817 30481 6851
rect 30515 6848 30527 6851
rect 30760 6848 30788 6956
rect 30834 6876 30840 6928
rect 30892 6876 30898 6928
rect 30944 6916 30972 6956
rect 31018 6944 31024 6996
rect 31076 6984 31082 6996
rect 31573 6987 31631 6993
rect 31573 6984 31585 6987
rect 31076 6956 31585 6984
rect 31076 6944 31082 6956
rect 31573 6953 31585 6956
rect 31619 6953 31631 6987
rect 35250 6984 35256 6996
rect 31573 6947 31631 6953
rect 34808 6956 35256 6984
rect 33781 6919 33839 6925
rect 30944 6888 31432 6916
rect 30515 6820 30788 6848
rect 31404 6848 31432 6888
rect 33781 6885 33793 6919
rect 33827 6916 33839 6919
rect 34330 6916 34336 6928
rect 33827 6888 34336 6916
rect 33827 6885 33839 6888
rect 33781 6879 33839 6885
rect 34330 6876 34336 6888
rect 34388 6876 34394 6928
rect 31404 6820 31708 6848
rect 30515 6817 30527 6820
rect 30469 6811 30527 6817
rect 30653 6783 30711 6789
rect 30653 6780 30665 6783
rect 30208 6752 30665 6780
rect 30653 6749 30665 6752
rect 30699 6780 30711 6783
rect 30742 6780 30748 6792
rect 30699 6752 30748 6780
rect 30699 6749 30711 6752
rect 30653 6743 30711 6749
rect 30742 6740 30748 6752
rect 30800 6740 30806 6792
rect 31021 6783 31079 6789
rect 31021 6776 31033 6783
rect 30852 6749 31033 6776
rect 31067 6780 31079 6783
rect 31110 6780 31116 6792
rect 31067 6752 31116 6780
rect 31067 6749 31079 6752
rect 30852 6748 31079 6749
rect 30285 6715 30343 6721
rect 30285 6712 30297 6715
rect 30024 6684 30297 6712
rect 29917 6675 29975 6681
rect 30285 6681 30297 6684
rect 30331 6712 30343 6715
rect 30852 6712 30880 6748
rect 31021 6743 31079 6748
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 31404 6789 31432 6820
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6749 31263 6783
rect 31205 6743 31263 6749
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6749 31447 6783
rect 31389 6743 31447 6749
rect 31220 6712 31248 6743
rect 31478 6740 31484 6792
rect 31536 6740 31542 6792
rect 31680 6789 31708 6820
rect 33410 6808 33416 6860
rect 33468 6808 33474 6860
rect 34808 6857 34836 6956
rect 35250 6944 35256 6956
rect 35308 6944 35314 6996
rect 33873 6851 33931 6857
rect 33873 6817 33885 6851
rect 33919 6817 33931 6851
rect 33873 6811 33931 6817
rect 34793 6851 34851 6857
rect 34793 6817 34805 6851
rect 34839 6817 34851 6851
rect 34793 6811 34851 6817
rect 36541 6851 36599 6857
rect 36541 6817 36553 6851
rect 36587 6817 36599 6851
rect 36541 6811 36599 6817
rect 31665 6783 31723 6789
rect 31665 6749 31677 6783
rect 31711 6749 31723 6783
rect 31665 6743 31723 6749
rect 33321 6783 33379 6789
rect 33321 6749 33333 6783
rect 33367 6780 33379 6783
rect 33888 6780 33916 6811
rect 33367 6752 33916 6780
rect 33367 6749 33379 6752
rect 33321 6743 33379 6749
rect 36078 6740 36084 6792
rect 36136 6780 36142 6792
rect 36556 6780 36584 6811
rect 37458 6808 37464 6860
rect 37516 6808 37522 6860
rect 38013 6851 38071 6857
rect 38013 6817 38025 6851
rect 38059 6848 38071 6851
rect 38194 6848 38200 6860
rect 38059 6820 38200 6848
rect 38059 6817 38071 6820
rect 38013 6811 38071 6817
rect 38194 6808 38200 6820
rect 38252 6808 38258 6860
rect 37274 6780 37280 6792
rect 36136 6752 36202 6780
rect 36556 6752 37280 6780
rect 36136 6740 36142 6752
rect 37274 6740 37280 6752
rect 37332 6740 37338 6792
rect 30331 6684 30880 6712
rect 31036 6684 31248 6712
rect 30331 6681 30343 6684
rect 30285 6675 30343 6681
rect 29707 6647 29765 6653
rect 29707 6644 29719 6647
rect 27908 6616 29719 6644
rect 29707 6613 29719 6616
rect 29753 6644 29765 6647
rect 30834 6644 30840 6656
rect 29753 6616 30840 6644
rect 29753 6613 29765 6616
rect 29707 6607 29765 6613
rect 30834 6604 30840 6616
rect 30892 6644 30898 6656
rect 31036 6644 31064 6684
rect 35066 6672 35072 6724
rect 35124 6672 35130 6724
rect 30892 6616 31064 6644
rect 30892 6604 30898 6616
rect 31294 6604 31300 6656
rect 31352 6604 31358 6656
rect 32858 6604 32864 6656
rect 32916 6644 32922 6656
rect 33137 6647 33195 6653
rect 33137 6644 33149 6647
rect 32916 6616 33149 6644
rect 32916 6604 32922 6616
rect 33137 6613 33149 6616
rect 33183 6613 33195 6647
rect 33137 6607 33195 6613
rect 36998 6604 37004 6656
rect 37056 6644 37062 6656
rect 37093 6647 37151 6653
rect 37093 6644 37105 6647
rect 37056 6616 37105 6644
rect 37056 6604 37062 6616
rect 37093 6613 37105 6616
rect 37139 6613 37151 6647
rect 37093 6607 37151 6613
rect 1104 6554 44620 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 44620 6554
rect 1104 6480 44620 6502
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 8036 6412 11928 6440
rect 3160 6372 3188 6400
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3160 6344 3801 6372
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 4798 6332 4804 6384
rect 4856 6332 4862 6384
rect 5276 6372 5304 6403
rect 8036 6372 8064 6412
rect 5276 6344 8064 6372
rect 8202 6332 8208 6384
rect 8260 6332 8266 6384
rect 10505 6375 10563 6381
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 10551 6344 11376 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 11348 6316 11376 6344
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9858 6304 9864 6316
rect 9447 6276 9864 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9858 6264 9864 6276
rect 9916 6304 9922 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 9916 6276 10333 6304
rect 9916 6264 9922 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11146 6304 11152 6316
rect 11011 6276 11152 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11238 6264 11244 6316
rect 11296 6264 11302 6316
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11388 6276 11713 6304
rect 11388 6264 11394 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6236 3571 6239
rect 7374 6236 7380 6248
rect 3559 6208 7380 6236
rect 3559 6205 3571 6208
rect 3513 6199 3571 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10226 6236 10232 6248
rect 10183 6208 10232 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11256 6236 11284 6264
rect 10744 6208 11284 6236
rect 11793 6239 11851 6245
rect 10744 6196 10750 6208
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 11900 6236 11928 6412
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 14550 6440 14556 6452
rect 12676 6412 14556 6440
rect 12676 6400 12682 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14918 6400 14924 6452
rect 14976 6400 14982 6452
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 12636 6372 12664 6400
rect 13630 6372 13636 6384
rect 12216 6344 12664 6372
rect 12728 6344 13636 6372
rect 12216 6332 12222 6344
rect 12250 6264 12256 6316
rect 12308 6264 12314 6316
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12728 6304 12756 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 13998 6372 14004 6384
rect 13955 6344 14004 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 14182 6332 14188 6384
rect 14240 6372 14246 6384
rect 14286 6375 14344 6381
rect 14286 6372 14298 6375
rect 14240 6344 14298 6372
rect 14240 6332 14246 6344
rect 14286 6341 14298 6344
rect 14332 6341 14344 6375
rect 15120 6372 15148 6403
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16301 6443 16359 6449
rect 15436 6412 16160 6440
rect 15436 6400 15442 6412
rect 16132 6372 16160 6412
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 16666 6440 16672 6452
rect 16347 6412 16672 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 17770 6440 17776 6452
rect 16899 6412 17776 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 15120 6344 15884 6372
rect 16132 6344 16804 6372
rect 14286 6335 14344 6341
rect 12483 6276 12756 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14700 6276 14841 6304
rect 14700 6264 14706 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 11900 6208 12909 6236
rect 11793 6199 11851 6205
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 7392 6100 7420 6196
rect 11808 6168 11836 6199
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 15028 6236 15056 6267
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15381 6307 15439 6313
rect 15381 6304 15393 6307
rect 15160 6276 15393 6304
rect 15160 6264 15166 6276
rect 15381 6273 15393 6276
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 15856 6313 15884 6344
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16172 6276 16681 6304
rect 16172 6264 16178 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 13044 6208 15301 6236
rect 13044 6196 13050 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 15930 6236 15936 6248
rect 15611 6208 15936 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 13630 6168 13636 6180
rect 11808 6140 13636 6168
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 14826 6168 14832 6180
rect 14292 6140 14832 6168
rect 8110 6100 8116 6112
rect 7392 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 12618 6100 12624 6112
rect 11204 6072 12624 6100
rect 11204 6060 11210 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 13354 6100 13360 6112
rect 12759 6072 13360 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14292 6109 14320 6140
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15488 6168 15516 6199
rect 15930 6196 15936 6208
rect 15988 6196 15994 6248
rect 16776 6236 16804 6344
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 17052 6313 17080 6412
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 21910 6440 21916 6452
rect 20211 6412 21916 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 22462 6400 22468 6452
rect 22520 6400 22526 6452
rect 25682 6400 25688 6452
rect 25740 6440 25746 6452
rect 27798 6440 27804 6452
rect 25740 6412 27804 6440
rect 25740 6400 25746 6412
rect 27798 6400 27804 6412
rect 27856 6400 27862 6452
rect 28810 6400 28816 6452
rect 28868 6400 28874 6452
rect 35066 6400 35072 6452
rect 35124 6440 35130 6452
rect 35713 6443 35771 6449
rect 35713 6440 35725 6443
rect 35124 6412 35725 6440
rect 35124 6400 35130 6412
rect 35713 6409 35725 6412
rect 35759 6409 35771 6443
rect 35713 6403 35771 6409
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 17543 6344 18368 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 17048 6307 17106 6313
rect 17048 6273 17060 6307
rect 17094 6273 17106 6307
rect 17048 6267 17106 6273
rect 17310 6264 17316 6316
rect 17368 6264 17374 6316
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 17586 6264 17592 6316
rect 17644 6264 17650 6316
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 17954 6304 17960 6316
rect 17911 6276 17960 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 16776 6208 17233 6236
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17420 6236 17448 6264
rect 17788 6236 17816 6267
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18340 6313 18368 6344
rect 22112 6344 22508 6372
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18064 6236 18092 6267
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 22112 6248 22140 6344
rect 22480 6313 22508 6344
rect 27430 6332 27436 6384
rect 27488 6332 27494 6384
rect 28828 6372 28856 6400
rect 28828 6344 29224 6372
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6273 22707 6307
rect 22649 6267 22707 6273
rect 17420 6208 17816 6236
rect 17221 6199 17279 6205
rect 14976 6140 15516 6168
rect 14976 6128 14982 6140
rect 15838 6128 15844 6180
rect 15896 6168 15902 6180
rect 16206 6168 16212 6180
rect 15896 6140 16212 6168
rect 15896 6128 15902 6140
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 17126 6128 17132 6180
rect 17184 6128 17190 6180
rect 14277 6103 14335 6109
rect 14277 6100 14289 6103
rect 13780 6072 14289 6100
rect 13780 6060 13786 6072
rect 14277 6069 14289 6072
rect 14323 6069 14335 6103
rect 14277 6063 14335 6069
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 14424 6072 14473 6100
rect 14424 6060 14430 6072
rect 14461 6069 14473 6072
rect 14507 6100 14519 6103
rect 15102 6100 15108 6112
rect 14507 6072 15108 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17310 6100 17316 6112
rect 17000 6072 17316 6100
rect 17000 6060 17006 6072
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17788 6100 17816 6208
rect 17880 6208 18092 6236
rect 17880 6180 17908 6208
rect 18506 6196 18512 6248
rect 18564 6196 18570 6248
rect 19362 6239 19420 6245
rect 19362 6236 19374 6239
rect 18800 6208 19374 6236
rect 17862 6128 17868 6180
rect 17920 6128 17926 6180
rect 17954 6128 17960 6180
rect 18012 6128 18018 6180
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6168 18291 6171
rect 18800 6168 18828 6208
rect 19362 6205 19374 6208
rect 19408 6205 19420 6239
rect 19362 6199 19420 6205
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 20162 6236 20168 6248
rect 19567 6208 20168 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 22094 6196 22100 6248
rect 22152 6196 22158 6248
rect 22388 6236 22416 6267
rect 22554 6236 22560 6248
rect 22388 6208 22560 6236
rect 22554 6196 22560 6208
rect 22612 6236 22618 6248
rect 22664 6236 22692 6267
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 27065 6307 27123 6313
rect 27065 6304 27077 6307
rect 26568 6276 27077 6304
rect 26568 6264 26574 6276
rect 27065 6273 27077 6276
rect 27111 6273 27123 6307
rect 27065 6267 27123 6273
rect 28812 6307 28870 6313
rect 28812 6273 28824 6307
rect 28858 6273 28870 6307
rect 28812 6267 28870 6273
rect 22612 6208 22692 6236
rect 28827 6236 28855 6267
rect 28902 6264 28908 6316
rect 28960 6264 28966 6316
rect 28997 6307 29055 6313
rect 28997 6273 29009 6307
rect 29043 6304 29055 6307
rect 29086 6304 29092 6316
rect 29043 6276 29092 6304
rect 29043 6273 29055 6276
rect 28997 6267 29055 6273
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 29196 6313 29224 6344
rect 29181 6307 29239 6313
rect 29181 6273 29193 6307
rect 29227 6273 29239 6307
rect 29181 6267 29239 6273
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6273 35863 6307
rect 35805 6267 35863 6273
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6304 37519 6307
rect 38194 6304 38200 6316
rect 37507 6276 38200 6304
rect 37507 6273 37519 6276
rect 37461 6267 37519 6273
rect 35820 6236 35848 6267
rect 38194 6264 38200 6276
rect 38252 6264 38258 6316
rect 36998 6236 37004 6248
rect 28827 6208 28994 6236
rect 35820 6208 37004 6236
rect 22612 6196 22618 6208
rect 28966 6180 28994 6208
rect 36998 6196 37004 6208
rect 37056 6236 37062 6248
rect 37369 6239 37427 6245
rect 37369 6236 37381 6239
rect 37056 6208 37381 6236
rect 37056 6196 37062 6208
rect 37369 6205 37381 6208
rect 37415 6205 37427 6239
rect 37369 6199 37427 6205
rect 37829 6239 37887 6245
rect 37829 6205 37841 6239
rect 37875 6236 37887 6239
rect 38930 6236 38936 6248
rect 37875 6208 38936 6236
rect 37875 6205 37887 6208
rect 37829 6199 37887 6205
rect 38930 6196 38936 6208
rect 38988 6196 38994 6248
rect 18279 6140 18828 6168
rect 18969 6171 19027 6177
rect 18279 6137 18291 6140
rect 18233 6131 18291 6137
rect 18969 6137 18981 6171
rect 19015 6137 19027 6171
rect 18969 6131 19027 6137
rect 18046 6100 18052 6112
rect 17788 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 18984 6100 19012 6131
rect 21174 6128 21180 6180
rect 21232 6168 21238 6180
rect 21821 6171 21879 6177
rect 21821 6168 21833 6171
rect 21232 6140 21833 6168
rect 21232 6128 21238 6140
rect 21821 6137 21833 6140
rect 21867 6137 21879 6171
rect 21821 6131 21879 6137
rect 28537 6171 28595 6177
rect 28537 6137 28549 6171
rect 28583 6137 28595 6171
rect 28966 6140 29000 6180
rect 28537 6131 28595 6137
rect 18840 6072 19012 6100
rect 22281 6103 22339 6109
rect 18840 6060 18846 6072
rect 22281 6069 22293 6103
rect 22327 6100 22339 6103
rect 22922 6100 22928 6112
rect 22327 6072 22928 6100
rect 22327 6069 22339 6072
rect 22281 6063 22339 6069
rect 22922 6060 22928 6072
rect 22980 6100 22986 6112
rect 28552 6100 28580 6131
rect 28994 6128 29000 6140
rect 29052 6128 29058 6180
rect 22980 6072 28580 6100
rect 22980 6060 22986 6072
rect 1104 6010 44620 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 44620 6010
rect 1104 5936 44620 5958
rect 6914 5856 6920 5908
rect 6972 5856 6978 5908
rect 12894 5856 12900 5908
rect 12952 5856 12958 5908
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13412 5868 13584 5896
rect 13412 5856 13418 5868
rect 6932 5760 6960 5856
rect 12529 5831 12587 5837
rect 12529 5797 12541 5831
rect 12575 5828 12587 5831
rect 12575 5800 13446 5828
rect 12575 5797 12587 5800
rect 12529 5791 12587 5797
rect 6748 5732 6960 5760
rect 12544 5732 13308 5760
rect 6748 5701 6776 5732
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12544 5701 12572 5732
rect 13280 5701 13308 5732
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12492 5664 12541 5692
rect 12492 5652 12498 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 12820 5624 12848 5655
rect 12894 5624 12900 5636
rect 12820 5596 12900 5624
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 6546 5516 6552 5568
rect 6604 5516 6610 5568
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 12250 5556 12256 5568
rect 10836 5528 12256 5556
rect 10836 5516 10842 5528
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 12986 5556 12992 5568
rect 12759 5528 12992 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13096 5556 13124 5655
rect 13170 5584 13176 5636
rect 13228 5584 13234 5636
rect 13418 5633 13446 5800
rect 13556 5760 13584 5868
rect 13630 5856 13636 5908
rect 13688 5856 13694 5908
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 15746 5896 15752 5908
rect 14608 5868 15752 5896
rect 14608 5856 14614 5868
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 16080 5868 16221 5896
rect 16080 5856 16086 5868
rect 16209 5865 16221 5868
rect 16255 5865 16267 5899
rect 16209 5859 16267 5865
rect 16393 5899 16451 5905
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 17218 5896 17224 5908
rect 16439 5868 17224 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17862 5856 17868 5908
rect 17920 5856 17926 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 18506 5896 18512 5908
rect 18371 5868 18512 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19334 5856 19340 5908
rect 19392 5856 19398 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 19484 5868 19717 5896
rect 19484 5856 19490 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 19705 5859 19763 5865
rect 21913 5899 21971 5905
rect 21913 5865 21925 5899
rect 21959 5896 21971 5899
rect 23290 5896 23296 5908
rect 21959 5868 23296 5896
rect 21959 5865 21971 5868
rect 21913 5859 21971 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24670 5896 24676 5908
rect 24259 5868 24676 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 32664 5899 32722 5905
rect 32664 5865 32676 5899
rect 32710 5896 32722 5899
rect 32858 5896 32864 5908
rect 32710 5868 32864 5896
rect 32710 5865 32722 5868
rect 32664 5859 32722 5865
rect 32858 5856 32864 5868
rect 32916 5856 32922 5908
rect 13648 5828 13676 5856
rect 15565 5831 15623 5837
rect 13648 5800 13952 5828
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13556 5732 13645 5760
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 13924 5704 13952 5800
rect 15565 5797 15577 5831
rect 15611 5828 15623 5831
rect 18690 5828 18696 5840
rect 15611 5800 18696 5828
rect 15611 5797 15623 5800
rect 15565 5791 15623 5797
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17000 5732 18184 5760
rect 17000 5720 17006 5732
rect 18156 5704 18184 5732
rect 18598 5720 18604 5772
rect 18656 5760 18662 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18656 5732 19257 5760
rect 18656 5720 18662 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19352 5760 19380 5856
rect 24578 5788 24584 5840
rect 24636 5788 24642 5840
rect 20441 5763 20499 5769
rect 20441 5760 20453 5763
rect 19352 5732 20453 5760
rect 19245 5723 19303 5729
rect 20441 5729 20453 5732
rect 20487 5729 20499 5763
rect 20441 5723 20499 5729
rect 22094 5720 22100 5772
rect 22152 5760 22158 5772
rect 25222 5760 25228 5772
rect 22152 5732 23520 5760
rect 22152 5720 22158 5732
rect 23492 5704 23520 5732
rect 23768 5732 25228 5760
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 13814 5652 13820 5704
rect 13872 5652 13878 5704
rect 13906 5652 13912 5704
rect 13964 5652 13970 5704
rect 14090 5652 14096 5704
rect 14148 5652 14154 5704
rect 15010 5652 15016 5704
rect 15068 5692 15074 5704
rect 15473 5695 15531 5701
rect 15473 5692 15485 5695
rect 15068 5664 15485 5692
rect 15068 5652 15074 5664
rect 15473 5661 15485 5664
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 13403 5627 13461 5633
rect 13403 5593 13415 5627
rect 13449 5624 13461 5627
rect 14108 5624 14136 5652
rect 13449 5596 14136 5624
rect 15488 5624 15516 5655
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 15804 5664 16160 5692
rect 15804 5652 15810 5664
rect 15841 5627 15899 5633
rect 15841 5624 15853 5627
rect 15488 5596 15853 5624
rect 13449 5593 13461 5596
rect 13403 5587 13461 5593
rect 15841 5593 15853 5596
rect 15887 5593 15899 5627
rect 15841 5587 15899 5593
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5593 16083 5627
rect 16025 5587 16083 5593
rect 13633 5559 13691 5565
rect 13633 5556 13645 5559
rect 13096 5528 13645 5556
rect 13633 5525 13645 5528
rect 13679 5525 13691 5559
rect 13633 5519 13691 5525
rect 14182 5516 14188 5568
rect 14240 5556 14246 5568
rect 15654 5556 15660 5568
rect 14240 5528 15660 5556
rect 14240 5516 14246 5528
rect 15654 5516 15660 5528
rect 15712 5556 15718 5568
rect 16040 5556 16068 5587
rect 15712 5528 16068 5556
rect 16132 5556 16160 5664
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 16264 5664 16313 5692
rect 16264 5652 16270 5664
rect 16301 5661 16313 5664
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17678 5692 17684 5704
rect 16816 5664 17684 5692
rect 16816 5652 16822 5664
rect 17678 5652 17684 5664
rect 17736 5692 17742 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17736 5664 17785 5692
rect 17736 5652 17742 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18046 5652 18052 5704
rect 18104 5652 18110 5704
rect 18138 5652 18144 5704
rect 18196 5652 18202 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 18340 5664 19349 5692
rect 18230 5624 18236 5636
rect 16592 5596 18236 5624
rect 16592 5556 16620 5596
rect 18230 5584 18236 5596
rect 18288 5584 18294 5636
rect 16132 5528 16620 5556
rect 15712 5516 15718 5528
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 18340 5556 18368 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 19352 5624 19380 5655
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 19521 5695 19579 5701
rect 19521 5692 19533 5695
rect 19484 5664 19533 5692
rect 19484 5652 19490 5664
rect 19521 5661 19533 5664
rect 19567 5661 19579 5695
rect 19521 5655 19579 5661
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 22281 5695 22339 5701
rect 22281 5661 22293 5695
rect 22327 5661 22339 5695
rect 22281 5655 22339 5661
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22557 5695 22615 5701
rect 22557 5692 22569 5695
rect 22511 5664 22569 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22557 5661 22569 5664
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 20438 5624 20444 5636
rect 19352 5596 20444 5624
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 20530 5584 20536 5636
rect 20588 5624 20594 5636
rect 20898 5624 20904 5636
rect 20588 5596 20904 5624
rect 20588 5584 20594 5596
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 22296 5624 22324 5655
rect 23474 5652 23480 5704
rect 23532 5692 23538 5704
rect 23768 5701 23796 5732
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 32401 5763 32459 5769
rect 32401 5729 32413 5763
rect 32447 5760 32459 5763
rect 32766 5760 32772 5772
rect 32447 5732 32772 5760
rect 32447 5729 32459 5732
rect 32401 5723 32459 5729
rect 32766 5720 32772 5732
rect 32824 5760 32830 5772
rect 33134 5760 33140 5772
rect 32824 5732 33140 5760
rect 32824 5720 32830 5732
rect 33134 5720 33140 5732
rect 33192 5720 33198 5772
rect 23753 5695 23811 5701
rect 23753 5692 23765 5695
rect 23532 5664 23765 5692
rect 23532 5652 23538 5664
rect 23753 5661 23765 5664
rect 23799 5661 23811 5695
rect 23753 5655 23811 5661
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 24075 5664 24409 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 24397 5661 24409 5664
rect 24443 5692 24455 5695
rect 24670 5692 24676 5704
rect 24443 5664 24676 5692
rect 24443 5661 24455 5664
rect 24397 5655 24455 5661
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 25133 5695 25191 5701
rect 25133 5661 25145 5695
rect 25179 5692 25191 5695
rect 26050 5692 26056 5704
rect 25179 5664 26056 5692
rect 25179 5661 25191 5664
rect 25133 5655 25191 5661
rect 22296 5596 22600 5624
rect 22572 5568 22600 5596
rect 23382 5584 23388 5636
rect 23440 5624 23446 5636
rect 23845 5627 23903 5633
rect 23845 5624 23857 5627
rect 23440 5596 23857 5624
rect 23440 5584 23446 5596
rect 23845 5593 23857 5596
rect 23891 5624 23903 5627
rect 25148 5624 25176 5655
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 23891 5596 25176 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 33318 5584 33324 5636
rect 33376 5584 33382 5636
rect 16724 5528 18368 5556
rect 16724 5516 16730 5528
rect 22554 5516 22560 5568
rect 22612 5516 22618 5568
rect 22741 5559 22799 5565
rect 22741 5525 22753 5559
rect 22787 5556 22799 5559
rect 22830 5556 22836 5568
rect 22787 5528 22836 5556
rect 22787 5525 22799 5528
rect 22741 5519 22799 5525
rect 22830 5516 22836 5528
rect 22888 5556 22894 5568
rect 23750 5556 23756 5568
rect 22888 5528 23756 5556
rect 22888 5516 22894 5528
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 26418 5516 26424 5568
rect 26476 5556 26482 5568
rect 33042 5556 33048 5568
rect 26476 5528 33048 5556
rect 26476 5516 26482 5528
rect 33042 5516 33048 5528
rect 33100 5516 33106 5568
rect 34146 5516 34152 5568
rect 34204 5516 34210 5568
rect 1104 5466 44620 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 44620 5466
rect 1104 5392 44620 5414
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 8159 5355 8217 5361
rect 7248 5324 8064 5352
rect 7248 5312 7254 5324
rect 8036 5284 8064 5324
rect 8159 5321 8171 5355
rect 8205 5352 8217 5355
rect 8205 5324 9076 5352
rect 8205 5321 8217 5324
rect 8159 5315 8217 5321
rect 9048 5293 9076 5324
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10502 5352 10508 5364
rect 10008 5324 10508 5352
rect 10008 5312 10014 5324
rect 10502 5312 10508 5324
rect 10560 5352 10566 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10560 5324 10609 5352
rect 10560 5312 10566 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 10597 5315 10655 5321
rect 11057 5355 11115 5361
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 12066 5352 12072 5364
rect 11103 5324 12072 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 14366 5352 14372 5364
rect 13280 5324 14372 5352
rect 8665 5287 8723 5293
rect 8665 5284 8677 5287
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 7760 5216 7788 5270
rect 8036 5256 8677 5284
rect 8665 5253 8677 5256
rect 8711 5253 8723 5287
rect 8665 5247 8723 5253
rect 9033 5287 9091 5293
rect 9033 5253 9045 5287
rect 9079 5253 9091 5287
rect 10045 5287 10103 5293
rect 9033 5247 9091 5253
rect 9508 5256 9996 5284
rect 8202 5216 8208 5228
rect 7760 5188 8208 5216
rect 6365 5179 6423 5185
rect 6380 5012 6408 5179
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 6604 5120 6745 5148
rect 6604 5108 6610 5120
rect 6733 5117 6745 5120
rect 6779 5117 6791 5151
rect 8680 5148 8708 5247
rect 9048 5216 9076 5247
rect 9122 5216 9128 5228
rect 9048 5188 9128 5216
rect 9122 5176 9128 5188
rect 9180 5216 9186 5228
rect 9508 5225 9536 5256
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 9180 5188 9505 5216
rect 9180 5176 9186 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 9968 5225 9996 5256
rect 10045 5253 10057 5287
rect 10091 5253 10103 5287
rect 13280 5284 13308 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 14918 5352 14924 5364
rect 14424 5324 14924 5352
rect 14424 5312 14430 5324
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15562 5352 15568 5364
rect 15059 5324 15568 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 31757 5355 31815 5361
rect 31757 5321 31769 5355
rect 31803 5352 31815 5355
rect 32306 5352 32312 5364
rect 31803 5324 32312 5352
rect 31803 5321 31815 5324
rect 31757 5315 31815 5321
rect 32306 5312 32312 5324
rect 32364 5312 32370 5364
rect 10045 5247 10103 5253
rect 11808 5256 13308 5284
rect 13357 5287 13415 5293
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 10060 5216 10088 5247
rect 10226 5216 10232 5228
rect 10060 5188 10232 5216
rect 9953 5179 10011 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10042 5148 10048 5160
rect 8680 5120 10048 5148
rect 6733 5111 6791 5117
rect 10042 5108 10048 5120
rect 10100 5148 10106 5160
rect 10520 5148 10548 5179
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 11054 5176 11060 5228
rect 11112 5176 11118 5228
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 11701 5222 11759 5225
rect 11808 5222 11836 5256
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 13722 5284 13728 5296
rect 13403 5256 13728 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 14550 5284 14556 5296
rect 13964 5256 14556 5284
rect 13964 5244 13970 5256
rect 14550 5244 14556 5256
rect 14608 5284 14614 5296
rect 14608 5256 14964 5284
rect 14608 5244 14614 5256
rect 11701 5219 11836 5222
rect 11701 5185 11713 5219
rect 11747 5194 11836 5219
rect 11879 5219 11937 5225
rect 11747 5185 11759 5194
rect 11701 5179 11759 5185
rect 11879 5185 11891 5219
rect 11925 5185 11937 5219
rect 11879 5179 11937 5185
rect 11072 5148 11100 5176
rect 11900 5148 11928 5179
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 13262 5216 13268 5228
rect 12676 5188 13268 5216
rect 12676 5176 12682 5188
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14182 5216 14188 5228
rect 14016 5188 14188 5216
rect 10100 5120 11008 5148
rect 11072 5120 11928 5148
rect 10100 5108 10106 5120
rect 10980 5080 11008 5120
rect 10980 5052 11836 5080
rect 8110 5012 8116 5024
rect 6380 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 10318 5012 10324 5024
rect 9907 4984 10324 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10318 4972 10324 4984
rect 10376 5012 10382 5024
rect 10962 5012 10968 5024
rect 10376 4984 10968 5012
rect 10376 4972 10382 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11808 5012 11836 5052
rect 11882 5040 11888 5092
rect 11940 5040 11946 5092
rect 12158 5040 12164 5092
rect 12216 5080 12222 5092
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 12216 5052 13001 5080
rect 12216 5040 12222 5052
rect 12989 5049 13001 5052
rect 13035 5080 13047 5083
rect 13906 5080 13912 5092
rect 13035 5052 13912 5080
rect 13035 5049 13047 5052
rect 12989 5043 13047 5049
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14016 5012 14044 5188
rect 14182 5176 14188 5188
rect 14240 5216 14246 5228
rect 14936 5225 14964 5256
rect 15102 5244 15108 5296
rect 15160 5284 15166 5296
rect 16666 5284 16672 5296
rect 15160 5256 16672 5284
rect 15160 5244 15166 5256
rect 16666 5244 16672 5256
rect 16724 5244 16730 5296
rect 26145 5287 26203 5293
rect 26145 5253 26157 5287
rect 26191 5284 26203 5287
rect 26510 5284 26516 5296
rect 26191 5256 26516 5284
rect 26191 5253 26203 5256
rect 26145 5247 26203 5253
rect 26510 5244 26516 5256
rect 26568 5244 26574 5296
rect 32217 5287 32275 5293
rect 32217 5284 32229 5287
rect 31312 5256 32229 5284
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14240 5188 14749 5216
rect 14240 5176 14246 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15194 5216 15200 5228
rect 14967 5188 15200 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5185 22431 5219
rect 22373 5179 22431 5185
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 23382 5216 23388 5228
rect 22603 5188 23388 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15746 5148 15752 5160
rect 14700 5120 15752 5148
rect 14700 5108 14706 5120
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 22388 5148 22416 5179
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 25222 5176 25228 5228
rect 25280 5216 25286 5228
rect 26234 5216 26240 5228
rect 25280 5188 26240 5216
rect 25280 5176 25286 5188
rect 26234 5176 26240 5188
rect 26292 5176 26298 5228
rect 26528 5216 26556 5244
rect 26597 5219 26655 5225
rect 26597 5216 26609 5219
rect 26528 5188 26609 5216
rect 26597 5185 26609 5188
rect 26643 5185 26655 5219
rect 26597 5179 26655 5185
rect 30926 5176 30932 5228
rect 30984 5216 30990 5228
rect 31021 5219 31079 5225
rect 31021 5216 31033 5219
rect 30984 5188 31033 5216
rect 30984 5176 30990 5188
rect 31021 5185 31033 5188
rect 31067 5185 31079 5219
rect 31021 5179 31079 5185
rect 22388 5120 22876 5148
rect 22848 5092 22876 5120
rect 28994 5108 29000 5160
rect 29052 5108 29058 5160
rect 31036 5148 31064 5179
rect 31202 5176 31208 5228
rect 31260 5176 31266 5228
rect 31312 5225 31340 5256
rect 32217 5253 32229 5256
rect 32263 5253 32275 5287
rect 32217 5247 32275 5253
rect 33137 5287 33195 5293
rect 33137 5253 33149 5287
rect 33183 5284 33195 5287
rect 33226 5284 33232 5296
rect 33183 5256 33232 5284
rect 33183 5253 33195 5256
rect 33137 5247 33195 5253
rect 33226 5244 33232 5256
rect 33284 5244 33290 5296
rect 33778 5244 33784 5296
rect 33836 5244 33842 5296
rect 31297 5219 31355 5225
rect 31297 5185 31309 5219
rect 31343 5185 31355 5219
rect 31297 5179 31355 5185
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5185 31447 5219
rect 31573 5219 31631 5225
rect 31573 5216 31585 5219
rect 31389 5179 31447 5185
rect 31496 5188 31585 5216
rect 31404 5148 31432 5179
rect 31036 5120 31432 5148
rect 22830 5040 22836 5092
rect 22888 5040 22894 5092
rect 25777 5083 25835 5089
rect 25777 5049 25789 5083
rect 25823 5080 25835 5083
rect 26050 5080 26056 5092
rect 25823 5052 26056 5080
rect 25823 5049 25835 5052
rect 25777 5043 25835 5049
rect 26050 5040 26056 5052
rect 26108 5040 26114 5092
rect 31021 5083 31079 5089
rect 31021 5049 31033 5083
rect 31067 5080 31079 5083
rect 31110 5080 31116 5092
rect 31067 5052 31116 5080
rect 31067 5049 31079 5052
rect 31021 5043 31079 5049
rect 31110 5040 31116 5052
rect 31168 5040 31174 5092
rect 11808 4984 14044 5012
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 23014 5012 23020 5024
rect 22612 4984 23020 5012
rect 22612 4972 22618 4984
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 23658 4972 23664 5024
rect 23716 5012 23722 5024
rect 25590 5012 25596 5024
rect 23716 4984 25596 5012
rect 23716 4972 23722 4984
rect 25590 4972 25596 4984
rect 25648 5012 25654 5024
rect 26513 5015 26571 5021
rect 26513 5012 26525 5015
rect 25648 4984 26525 5012
rect 25648 4972 25654 4984
rect 26513 4981 26525 4984
rect 26559 5012 26571 5015
rect 27062 5012 27068 5024
rect 26559 4984 27068 5012
rect 26559 4981 26571 4984
rect 26513 4975 26571 4981
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 28350 4972 28356 5024
rect 28408 4972 28414 5024
rect 30650 4972 30656 5024
rect 30708 5012 30714 5024
rect 31496 5012 31524 5188
rect 31573 5185 31585 5188
rect 31619 5216 31631 5219
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 31619 5188 32137 5216
rect 31619 5185 31631 5188
rect 31573 5179 31631 5185
rect 32125 5185 32137 5188
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 32766 5176 32772 5228
rect 32824 5216 32830 5228
rect 32861 5219 32919 5225
rect 32861 5216 32873 5219
rect 32824 5188 32873 5216
rect 32824 5176 32830 5188
rect 32861 5185 32873 5188
rect 32907 5185 32919 5219
rect 32861 5179 32919 5185
rect 31570 5040 31576 5092
rect 31628 5080 31634 5092
rect 32122 5080 32128 5092
rect 31628 5052 32128 5080
rect 31628 5040 31634 5052
rect 32122 5040 32128 5052
rect 32180 5040 32186 5092
rect 30708 4984 31524 5012
rect 30708 4972 30714 4984
rect 32030 4972 32036 5024
rect 32088 5012 32094 5024
rect 33318 5012 33324 5024
rect 32088 4984 33324 5012
rect 32088 4972 32094 4984
rect 33318 4972 33324 4984
rect 33376 4972 33382 5024
rect 34606 4972 34612 5024
rect 34664 4972 34670 5024
rect 1104 4922 44620 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 44620 4922
rect 1104 4848 44620 4870
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4777 11115 4811
rect 11057 4771 11115 4777
rect 10689 4743 10747 4749
rect 10689 4709 10701 4743
rect 10735 4709 10747 4743
rect 11072 4740 11100 4771
rect 11238 4768 11244 4820
rect 11296 4768 11302 4820
rect 11330 4768 11336 4820
rect 11388 4768 11394 4820
rect 11422 4768 11428 4820
rect 11480 4768 11486 4820
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 11790 4808 11796 4820
rect 11747 4780 11796 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13136 4780 13277 4808
rect 13136 4768 13142 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13412 4780 13737 4808
rect 13412 4768 13418 4780
rect 13725 4777 13737 4780
rect 13771 4808 13783 4811
rect 13814 4808 13820 4820
rect 13771 4780 13820 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15620 4780 15853 4808
rect 15620 4768 15626 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 19150 4768 19156 4820
rect 19208 4808 19214 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 19208 4780 19257 4808
rect 19208 4768 19214 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 22741 4811 22799 4817
rect 22741 4777 22753 4811
rect 22787 4808 22799 4811
rect 23382 4808 23388 4820
rect 22787 4780 23388 4808
rect 22787 4777 22799 4780
rect 22741 4771 22799 4777
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 29362 4768 29368 4820
rect 29420 4768 29426 4820
rect 30650 4768 30656 4820
rect 30708 4768 30714 4820
rect 34793 4811 34851 4817
rect 30760 4780 32904 4808
rect 11348 4740 11376 4768
rect 11072 4712 11376 4740
rect 10689 4703 10747 4709
rect 10704 4672 10732 4703
rect 11440 4672 11468 4768
rect 9692 4644 10640 4672
rect 10704 4644 11468 4672
rect 11808 4672 11836 4768
rect 12360 4712 13672 4740
rect 12360 4672 12388 4712
rect 11808 4644 12388 4672
rect 9692 4616 9720 4644
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7834 4604 7840 4616
rect 7055 4576 7840 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 9858 4564 9864 4616
rect 9916 4564 9922 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 10612 4613 10640 4644
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 11606 4604 11612 4616
rect 10643 4576 10916 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 7190 4428 7196 4480
rect 7248 4428 7254 4480
rect 10520 4468 10548 4564
rect 10888 4545 10916 4576
rect 11256 4576 11612 4604
rect 10873 4539 10931 4545
rect 10873 4505 10885 4539
rect 10919 4505 10931 4539
rect 10873 4499 10931 4505
rect 11054 4496 11060 4548
rect 11112 4545 11118 4548
rect 11112 4539 11136 4545
rect 11124 4536 11136 4539
rect 11256 4536 11284 4576
rect 11606 4564 11612 4576
rect 11664 4604 11670 4616
rect 12360 4613 12388 4644
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4672 12495 4675
rect 13446 4672 13452 4684
rect 12483 4644 13452 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11664 4576 12081 4604
rect 11664 4564 11670 4576
rect 12069 4573 12081 4576
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12584 4576 12633 4604
rect 12584 4564 12590 4576
rect 12621 4573 12633 4576
rect 12667 4604 12679 4607
rect 12710 4604 12716 4616
rect 12667 4576 12716 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12820 4613 12848 4644
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13644 4672 13672 4712
rect 13924 4712 15700 4740
rect 13924 4684 13952 4712
rect 13906 4672 13912 4684
rect 13644 4644 13912 4672
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 11124 4508 11284 4536
rect 11124 4505 11136 4508
rect 11112 4499 11136 4505
rect 11112 4496 11118 4499
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11425 4539 11483 4545
rect 11425 4536 11437 4539
rect 11388 4508 11437 4536
rect 11388 4496 11394 4508
rect 11425 4505 11437 4508
rect 11471 4505 11483 4539
rect 13096 4536 13124 4567
rect 13262 4564 13268 4616
rect 13320 4604 13326 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13320 4576 13369 4604
rect 13320 4564 13326 4576
rect 13357 4573 13369 4576
rect 13403 4604 13415 4607
rect 13541 4607 13599 4613
rect 13403 4576 13492 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 13464 4536 13492 4576
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13644 4604 13672 4644
rect 13906 4632 13912 4644
rect 13964 4632 13970 4684
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 15010 4672 15016 4684
rect 14240 4644 15016 4672
rect 14240 4632 14246 4644
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 15672 4681 15700 4712
rect 15746 4700 15752 4752
rect 15804 4700 15810 4752
rect 18966 4700 18972 4752
rect 19024 4740 19030 4752
rect 19521 4743 19579 4749
rect 19521 4740 19533 4743
rect 19024 4712 19533 4740
rect 19024 4700 19030 4712
rect 19521 4709 19533 4712
rect 19567 4709 19579 4743
rect 23934 4740 23940 4752
rect 19521 4703 19579 4709
rect 23400 4712 23940 4740
rect 15657 4675 15715 4681
rect 15120 4644 15608 4672
rect 15120 4613 15148 4644
rect 15580 4616 15608 4644
rect 15657 4641 15669 4675
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 13587 4576 13672 4604
rect 15105 4607 15163 4613
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15470 4564 15476 4616
rect 15528 4564 15534 4616
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 15764 4604 15792 4700
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 18923 4644 19625 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19751 4644 20024 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15764 4576 15945 4604
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 18598 4604 18604 4616
rect 17184 4576 18604 4604
rect 17184 4564 17190 4576
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 15488 4536 15516 4564
rect 11425 4499 11483 4505
rect 11808 4508 13404 4536
rect 13464 4508 15516 4536
rect 15657 4539 15715 4545
rect 11808 4468 11836 4508
rect 10520 4440 11836 4468
rect 13376 4468 13404 4508
rect 15657 4505 15669 4539
rect 15703 4536 15715 4539
rect 17862 4536 17868 4548
rect 15703 4508 17868 4536
rect 15703 4505 15715 4508
rect 15657 4499 15715 4505
rect 17862 4496 17868 4508
rect 17920 4536 17926 4548
rect 18800 4536 18828 4567
rect 17920 4508 18828 4536
rect 17920 4496 17926 4508
rect 16390 4468 16396 4480
rect 13376 4440 16396 4468
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 18984 4468 19012 4567
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4573 19947 4607
rect 19889 4567 19947 4573
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 19904 4536 19932 4567
rect 19392 4508 19932 4536
rect 19392 4496 19398 4508
rect 19996 4468 20024 4644
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22373 4607 22431 4613
rect 22373 4604 22385 4607
rect 22336 4576 22385 4604
rect 22336 4564 22342 4576
rect 22373 4573 22385 4576
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 23014 4564 23020 4616
rect 23072 4564 23078 4616
rect 23400 4613 23428 4712
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 28902 4700 28908 4752
rect 28960 4740 28966 4752
rect 30760 4740 30788 4780
rect 28960 4712 30788 4740
rect 28960 4700 28966 4712
rect 24026 4672 24032 4684
rect 23676 4644 24032 4672
rect 23676 4613 23704 4644
rect 24026 4632 24032 4644
rect 24084 4672 24090 4684
rect 27893 4675 27951 4681
rect 24084 4644 26556 4672
rect 24084 4632 24090 4644
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4573 23259 4607
rect 23201 4567 23259 4573
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 23661 4607 23719 4613
rect 23661 4573 23673 4607
rect 23707 4573 23719 4607
rect 23661 4567 23719 4573
rect 23216 4536 23244 4567
rect 23750 4564 23756 4616
rect 23808 4564 23814 4616
rect 24394 4564 24400 4616
rect 24452 4564 24458 4616
rect 26234 4564 26240 4616
rect 26292 4604 26298 4616
rect 26421 4607 26479 4613
rect 26421 4604 26433 4607
rect 26292 4576 26433 4604
rect 26292 4564 26298 4576
rect 26421 4573 26433 4576
rect 26467 4573 26479 4607
rect 26421 4567 26479 4573
rect 23569 4539 23627 4545
rect 23569 4536 23581 4539
rect 22940 4508 23581 4536
rect 18196 4440 20024 4468
rect 22741 4471 22799 4477
rect 18196 4428 18202 4440
rect 22741 4437 22753 4471
rect 22787 4468 22799 4471
rect 22830 4468 22836 4480
rect 22787 4440 22836 4468
rect 22787 4437 22799 4440
rect 22741 4431 22799 4437
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 22940 4477 22968 4508
rect 23569 4505 23581 4508
rect 23615 4505 23627 4539
rect 24673 4539 24731 4545
rect 24673 4536 24685 4539
rect 23569 4499 23627 4505
rect 23952 4508 24685 4536
rect 22925 4471 22983 4477
rect 22925 4437 22937 4471
rect 22971 4437 22983 4471
rect 22925 4431 22983 4437
rect 23106 4428 23112 4480
rect 23164 4428 23170 4480
rect 23952 4477 23980 4508
rect 24673 4505 24685 4508
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 25406 4496 25412 4548
rect 25464 4496 25470 4548
rect 23937 4471 23995 4477
rect 23937 4437 23949 4471
rect 23983 4437 23995 4471
rect 26528 4468 26556 4644
rect 27893 4641 27905 4675
rect 27939 4672 27951 4675
rect 28350 4672 28356 4684
rect 27939 4644 28356 4672
rect 27939 4641 27951 4644
rect 27893 4635 27951 4641
rect 28350 4632 28356 4644
rect 28408 4632 28414 4684
rect 32030 4672 32036 4684
rect 30944 4644 32036 4672
rect 27614 4564 27620 4616
rect 27672 4564 27678 4616
rect 29178 4536 29184 4548
rect 29118 4508 29184 4536
rect 29178 4496 29184 4508
rect 29236 4536 29242 4548
rect 30944 4536 30972 4644
rect 32030 4632 32036 4644
rect 32088 4632 32094 4684
rect 32401 4675 32459 4681
rect 32401 4641 32413 4675
rect 32447 4672 32459 4675
rect 32766 4672 32772 4684
rect 32447 4644 32772 4672
rect 32447 4641 32459 4644
rect 32401 4635 32459 4641
rect 32766 4632 32772 4644
rect 32824 4632 32830 4684
rect 32876 4672 32904 4780
rect 34793 4777 34805 4811
rect 34839 4777 34851 4811
rect 34793 4771 34851 4777
rect 33229 4743 33287 4749
rect 33229 4740 33241 4743
rect 33060 4712 33241 4740
rect 33060 4672 33088 4712
rect 33229 4709 33241 4712
rect 33275 4709 33287 4743
rect 33229 4703 33287 4709
rect 33413 4743 33471 4749
rect 33413 4709 33425 4743
rect 33459 4740 33471 4743
rect 34606 4740 34612 4752
rect 33459 4712 34612 4740
rect 33459 4709 33471 4712
rect 33413 4703 33471 4709
rect 34606 4700 34612 4712
rect 34664 4740 34670 4752
rect 34808 4740 34836 4771
rect 34664 4712 34836 4740
rect 34664 4700 34670 4712
rect 32876 4644 33088 4672
rect 33689 4607 33747 4613
rect 33689 4573 33701 4607
rect 33735 4604 33747 4607
rect 34146 4604 34152 4616
rect 33735 4576 34152 4604
rect 33735 4573 33747 4576
rect 33689 4567 33747 4573
rect 34146 4564 34152 4576
rect 34204 4564 34210 4616
rect 34425 4607 34483 4613
rect 34425 4573 34437 4607
rect 34471 4604 34483 4607
rect 34606 4604 34612 4616
rect 34471 4576 34612 4604
rect 34471 4573 34483 4576
rect 34425 4567 34483 4573
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34701 4607 34759 4613
rect 34701 4573 34713 4607
rect 34747 4573 34759 4607
rect 34701 4567 34759 4573
rect 29236 4522 30972 4536
rect 32125 4539 32183 4545
rect 29236 4508 30958 4522
rect 29236 4496 29242 4508
rect 32125 4505 32137 4539
rect 32171 4536 32183 4539
rect 33781 4539 33839 4545
rect 33781 4536 33793 4539
rect 32171 4508 33793 4536
rect 32171 4505 32183 4508
rect 32125 4499 32183 4505
rect 33781 4505 33793 4508
rect 33827 4505 33839 4539
rect 34164 4536 34192 4564
rect 34716 4536 34744 4567
rect 34164 4508 34744 4536
rect 33781 4499 33839 4505
rect 35161 4471 35219 4477
rect 35161 4468 35173 4471
rect 26528 4440 35173 4468
rect 23937 4431 23995 4437
rect 35161 4437 35173 4440
rect 35207 4437 35219 4471
rect 35161 4431 35219 4437
rect 1104 4378 44620 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 44620 4378
rect 1104 4304 44620 4326
rect 10796 4236 14136 4264
rect 8202 4156 8208 4208
rect 8260 4156 8266 4208
rect 9309 4199 9367 4205
rect 9309 4165 9321 4199
rect 9355 4196 9367 4199
rect 9858 4196 9864 4208
rect 9355 4168 9864 4196
rect 9355 4165 9367 4168
rect 9309 4159 9367 4165
rect 9858 4156 9864 4168
rect 9916 4196 9922 4208
rect 10045 4199 10103 4205
rect 10045 4196 10057 4199
rect 9916 4168 10057 4196
rect 9916 4156 9922 4168
rect 10045 4165 10057 4168
rect 10091 4165 10103 4199
rect 10045 4159 10103 4165
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7055 4100 7512 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7248 4032 7389 4060
rect 7248 4020 7254 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7484 4060 7512 4100
rect 9122 4088 9128 4140
rect 9180 4088 9186 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 8110 4060 8116 4072
rect 7484 4032 8116 4060
rect 7377 4023 7435 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9416 4060 9444 4091
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10796 4128 10824 4236
rect 12250 4196 12256 4208
rect 12176 4168 12256 4196
rect 10192 4100 10824 4128
rect 10192 4088 10198 4100
rect 9674 4060 9680 4072
rect 8895 4032 9680 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10410 4060 10416 4072
rect 9907 4032 10416 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10796 4060 10824 4100
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4097 11299 4131
rect 11241 4091 11299 4097
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10796 4032 10977 4060
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 11256 4060 11284 4091
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11388 4100 11713 4128
rect 11388 4088 11394 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12176 4128 12204 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 12124 4100 12204 4128
rect 12124 4088 12130 4100
rect 11422 4060 11428 4072
rect 11256 4032 11428 4060
rect 10965 4023 11023 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4060 11575 4063
rect 11606 4060 11612 4072
rect 11563 4032 11612 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 12342 4020 12348 4072
rect 12400 4020 12406 4072
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12710 4060 12716 4072
rect 12575 4032 12716 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12894 4020 12900 4072
rect 12952 4020 12958 4072
rect 13446 4069 13452 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 13096 4032 13277 4060
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 12912 3992 12940 4020
rect 13096 4004 13124 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13403 4063 13452 4069
rect 13403 4029 13415 4063
rect 13449 4029 13452 4063
rect 13403 4023 13452 4029
rect 13446 4020 13452 4023
rect 13504 4020 13510 4072
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 14108 4060 14136 4236
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 17954 4264 17960 4276
rect 14976 4236 17960 4264
rect 14976 4224 14982 4236
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 14737 4199 14795 4205
rect 14737 4196 14749 4199
rect 14424 4168 14749 4196
rect 14424 4156 14430 4168
rect 14737 4165 14749 4168
rect 14783 4165 14795 4199
rect 15197 4199 15255 4205
rect 15197 4196 15209 4199
rect 14737 4159 14795 4165
rect 14936 4168 15209 4196
rect 14936 4140 14964 4168
rect 15197 4165 15209 4168
rect 15243 4165 15255 4199
rect 15197 4159 15255 4165
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4128 14243 4131
rect 14274 4128 14280 4140
rect 14231 4100 14280 4128
rect 14231 4097 14243 4100
rect 14185 4091 14243 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14918 4088 14924 4140
rect 14976 4088 14982 4140
rect 15672 4137 15700 4236
rect 17954 4224 17960 4236
rect 18012 4264 18018 4276
rect 18966 4264 18972 4276
rect 18012 4236 18972 4264
rect 18012 4224 18018 4236
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 22465 4267 22523 4273
rect 22465 4233 22477 4267
rect 22511 4264 22523 4267
rect 23106 4264 23112 4276
rect 22511 4236 23112 4264
rect 22511 4233 22523 4236
rect 22465 4227 22523 4233
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 24670 4224 24676 4276
rect 24728 4224 24734 4276
rect 31846 4264 31852 4276
rect 28736 4236 31852 4264
rect 16206 4156 16212 4208
rect 16264 4196 16270 4208
rect 17773 4199 17831 4205
rect 16264 4168 16344 4196
rect 16264 4156 16270 4168
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15657 4131 15715 4137
rect 15059 4100 15608 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 13587 4032 14136 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 12032 3964 12848 3992
rect 12912 3964 13001 3992
rect 12032 3952 12038 3964
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3924 10379 3927
rect 10594 3924 10600 3936
rect 10367 3896 10600 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 12158 3924 12164 3936
rect 10652 3896 12164 3924
rect 10652 3884 10658 3896
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12820 3924 12848 3964
rect 12989 3961 13001 3964
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 13078 3952 13084 4004
rect 13136 3952 13142 4004
rect 13538 3924 13544 3936
rect 12820 3896 13544 3924
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 14734 3884 14740 3936
rect 14792 3884 14798 3936
rect 15470 3884 15476 3936
rect 15528 3884 15534 3936
rect 15580 3924 15608 4100
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 16114 4128 16120 4140
rect 15804 4100 16120 4128
rect 15804 4088 15810 4100
rect 16114 4088 16120 4100
rect 16172 4128 16178 4140
rect 16316 4137 16344 4168
rect 16500 4168 17172 4196
rect 16301 4131 16359 4137
rect 16172 4100 16252 4128
rect 16172 4088 16178 4100
rect 16224 4060 16252 4100
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16500 4137 16528 4168
rect 17144 4140 17172 4168
rect 17773 4165 17785 4199
rect 17819 4196 17831 4199
rect 17819 4168 18000 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 16485 4131 16543 4137
rect 16485 4128 16497 4131
rect 16448 4100 16497 4128
rect 16448 4088 16454 4100
rect 16485 4097 16497 4100
rect 16531 4097 16543 4131
rect 16485 4091 16543 4097
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17034 4128 17040 4140
rect 16899 4100 17040 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17126 4088 17132 4140
rect 17184 4088 17190 4140
rect 17221 4131 17279 4137
rect 17221 4097 17233 4131
rect 17267 4097 17279 4131
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17221 4091 17279 4097
rect 17328 4100 17509 4128
rect 17236 4060 17264 4091
rect 16224 4032 17264 4060
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 16301 3995 16359 4001
rect 15712 3964 16252 3992
rect 15712 3952 15718 3964
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15580 3896 15761 3924
rect 15749 3893 15761 3896
rect 15795 3924 15807 3927
rect 15930 3924 15936 3936
rect 15795 3896 15936 3924
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16224 3924 16252 3964
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 16482 3992 16488 4004
rect 16347 3964 16488 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 17328 3992 17356 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 17604 4060 17632 4091
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 17460 4032 17632 4060
rect 17460 4020 17466 4032
rect 16868 3964 17356 3992
rect 16868 3924 16896 3964
rect 17494 3952 17500 4004
rect 17552 3952 17558 4004
rect 16224 3896 16896 3924
rect 16942 3884 16948 3936
rect 17000 3884 17006 3936
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17368 3896 17417 3924
rect 17368 3884 17374 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17604 3924 17632 4032
rect 17972 4001 18000 4168
rect 21634 4156 21640 4208
rect 21692 4156 21698 4208
rect 22830 4156 22836 4208
rect 22888 4196 22894 4208
rect 23198 4196 23204 4208
rect 22888 4168 23204 4196
rect 22888 4156 22894 4168
rect 23198 4156 23204 4168
rect 23256 4196 23262 4208
rect 24688 4196 24716 4224
rect 28736 4205 28764 4236
rect 31846 4224 31852 4236
rect 31904 4224 31910 4276
rect 34606 4224 34612 4276
rect 34664 4264 34670 4276
rect 35345 4267 35403 4273
rect 35345 4264 35357 4267
rect 34664 4236 35357 4264
rect 34664 4224 34670 4236
rect 35345 4233 35357 4236
rect 35391 4233 35403 4267
rect 35345 4227 35403 4233
rect 23256 4168 24716 4196
rect 23256 4156 23262 4168
rect 18046 4088 18052 4140
rect 18104 4088 18110 4140
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 18322 4088 18328 4140
rect 18380 4088 18386 4140
rect 18414 4088 18420 4140
rect 18472 4088 18478 4140
rect 18598 4088 18604 4140
rect 18656 4088 18662 4140
rect 18874 4088 18880 4140
rect 18932 4138 18938 4140
rect 18932 4137 19098 4138
rect 18932 4131 19119 4137
rect 18932 4110 19073 4131
rect 18932 4088 18938 4110
rect 19061 4097 19073 4110
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 19426 4128 19432 4140
rect 19208 4100 19432 4128
rect 19208 4088 19214 4100
rect 19426 4088 19432 4100
rect 19484 4128 19490 4140
rect 19978 4128 19984 4140
rect 19484 4100 19984 4128
rect 19484 4088 19490 4100
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20162 4128 20168 4140
rect 20119 4100 20168 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 22554 4088 22560 4140
rect 22612 4088 22618 4140
rect 23492 4137 23520 4168
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4097 23535 4131
rect 23477 4091 23535 4097
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 24121 4131 24179 4137
rect 23799 4100 23980 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4029 18567 4063
rect 18616 4060 18644 4088
rect 18785 4063 18843 4069
rect 18785 4060 18797 4063
rect 18616 4032 18797 4060
rect 18509 4023 18567 4029
rect 18785 4029 18797 4032
rect 18831 4029 18843 4063
rect 19334 4060 19340 4072
rect 18785 4023 18843 4029
rect 18892 4032 19340 4060
rect 17957 3995 18015 4001
rect 17957 3961 17969 3995
rect 18003 3992 18015 3995
rect 18524 3992 18552 4023
rect 18003 3964 18552 3992
rect 18693 3995 18751 4001
rect 18003 3961 18015 3964
rect 17957 3955 18015 3961
rect 18693 3961 18705 3995
rect 18739 3992 18751 3995
rect 18892 3992 18920 4032
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 23842 4060 23848 4072
rect 22419 4032 23848 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 23952 4069 23980 4100
rect 24121 4097 24133 4131
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24351 4100 24532 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 23937 4063 23995 4069
rect 23937 4029 23949 4063
rect 23983 4029 23995 4063
rect 24136 4060 24164 4091
rect 24397 4063 24455 4069
rect 24136 4032 24348 4060
rect 23937 4023 23995 4029
rect 18739 3964 18920 3992
rect 18739 3961 18751 3964
rect 18693 3955 18751 3961
rect 18966 3952 18972 4004
rect 19024 3952 19030 4004
rect 22278 3952 22284 4004
rect 22336 3992 22342 4004
rect 23474 3992 23480 4004
rect 22336 3964 23480 3992
rect 22336 3952 22342 3964
rect 23474 3952 23480 3964
rect 23532 3952 23538 4004
rect 23566 3952 23572 4004
rect 23624 3952 23630 4004
rect 23658 3952 23664 4004
rect 23716 3952 23722 4004
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3961 24271 3995
rect 24213 3955 24271 3961
rect 18414 3924 18420 3936
rect 17604 3896 18420 3924
rect 17405 3887 17463 3893
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18874 3884 18880 3936
rect 18932 3884 18938 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 22925 3927 22983 3933
rect 22925 3924 22937 3927
rect 22520 3896 22937 3924
rect 22520 3884 22526 3896
rect 22925 3893 22937 3896
rect 22971 3893 22983 3927
rect 22925 3887 22983 3893
rect 23290 3884 23296 3936
rect 23348 3884 23354 3936
rect 23492 3924 23520 3952
rect 24228 3924 24256 3955
rect 23492 3896 24256 3924
rect 24320 3924 24348 4032
rect 24397 4029 24409 4063
rect 24443 4029 24455 4063
rect 24504 4060 24532 4100
rect 24578 4088 24584 4140
rect 24636 4088 24642 4140
rect 24688 4137 24716 4168
rect 28721 4199 28779 4205
rect 28721 4165 28733 4199
rect 28767 4165 28779 4199
rect 28721 4159 28779 4165
rect 29178 4156 29184 4208
rect 29236 4196 29242 4208
rect 29236 4168 29946 4196
rect 29236 4156 29242 4168
rect 36078 4156 36084 4208
rect 36136 4156 36142 4208
rect 24673 4131 24731 4137
rect 24673 4097 24685 4131
rect 24719 4097 24731 4131
rect 24673 4091 24731 4097
rect 24857 4131 24915 4137
rect 24857 4097 24869 4131
rect 24903 4128 24915 4131
rect 28902 4128 28908 4140
rect 24903 4100 28908 4128
rect 24903 4097 24915 4100
rect 24857 4091 24915 4097
rect 24765 4063 24823 4069
rect 24765 4060 24777 4063
rect 24504 4032 24777 4060
rect 24397 4023 24455 4029
rect 24765 4029 24777 4032
rect 24811 4029 24823 4063
rect 24765 4023 24823 4029
rect 24412 3992 24440 4023
rect 24486 3992 24492 4004
rect 24412 3964 24492 3992
rect 24486 3952 24492 3964
rect 24544 3992 24550 4004
rect 24872 3992 24900 4091
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 33042 4088 33048 4140
rect 33100 4128 33106 4140
rect 34790 4128 34796 4140
rect 33100 4100 34796 4128
rect 33100 4088 33106 4100
rect 34790 4088 34796 4100
rect 34848 4088 34854 4140
rect 37090 4088 37096 4140
rect 37148 4088 37154 4140
rect 29181 4063 29239 4069
rect 29181 4060 29193 4063
rect 27632 4032 29193 4060
rect 24544 3964 24900 3992
rect 24544 3952 24550 3964
rect 25406 3952 25412 4004
rect 25464 3992 25470 4004
rect 27522 3992 27528 4004
rect 25464 3964 27528 3992
rect 25464 3952 25470 3964
rect 27522 3952 27528 3964
rect 27580 3952 27586 4004
rect 27632 3936 27660 4032
rect 29181 4029 29193 4032
rect 29227 4029 29239 4063
rect 29181 4023 29239 4029
rect 29454 4020 29460 4072
rect 29512 4020 29518 4072
rect 30926 4020 30932 4072
rect 30984 4020 30990 4072
rect 36814 4020 36820 4072
rect 36872 4020 36878 4072
rect 24854 3924 24860 3936
rect 24320 3896 24860 3924
rect 24854 3884 24860 3896
rect 24912 3924 24918 3936
rect 26050 3924 26056 3936
rect 24912 3896 26056 3924
rect 24912 3884 24918 3896
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 27433 3927 27491 3933
rect 27433 3893 27445 3927
rect 27479 3924 27491 3927
rect 27614 3924 27620 3936
rect 27479 3896 27620 3924
rect 27479 3893 27491 3896
rect 27433 3887 27491 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 44620 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 44620 3834
rect 1104 3760 44620 3782
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 9306 3720 9312 3732
rect 8260 3692 9312 3720
rect 8260 3680 8266 3692
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9858 3720 9864 3732
rect 9508 3692 9864 3720
rect 9508 3528 9536 3692
rect 9858 3680 9864 3692
rect 9916 3720 9922 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 9916 3692 10333 3720
rect 9916 3680 9922 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10321 3683 10379 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11020 3692 12572 3720
rect 11020 3680 11026 3692
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3652 9643 3655
rect 11330 3652 11336 3664
rect 9631 3624 11336 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11425 3655 11483 3661
rect 11425 3621 11437 3655
rect 11471 3652 11483 3655
rect 11698 3652 11704 3664
rect 11471 3624 11704 3652
rect 11471 3621 11483 3624
rect 11425 3615 11483 3621
rect 11698 3612 11704 3624
rect 11756 3652 11762 3664
rect 12158 3652 12164 3664
rect 11756 3624 12164 3652
rect 11756 3612 11762 3624
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 12250 3612 12256 3664
rect 12308 3612 12314 3664
rect 12544 3652 12572 3692
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 12768 3692 13185 3720
rect 12768 3680 12774 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 14458 3720 14464 3732
rect 13780 3692 14464 3720
rect 13780 3680 13786 3692
rect 14458 3680 14464 3692
rect 14516 3720 14522 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14516 3692 14841 3720
rect 14516 3680 14522 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 15746 3680 15752 3732
rect 15804 3680 15810 3732
rect 16390 3720 16396 3732
rect 15856 3692 16396 3720
rect 12544 3624 13032 3652
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 10735 3556 12204 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9490 3516 9496 3528
rect 9263 3488 9496 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9732 3488 9781 3516
rect 9732 3476 9738 3488
rect 9769 3485 9781 3488
rect 9815 3516 9827 3519
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9815 3488 10241 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11514 3516 11520 3528
rect 11471 3488 11520 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 12066 3516 12072 3528
rect 11655 3488 12072 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 9401 3451 9459 3457
rect 9401 3417 9413 3451
rect 9447 3417 9459 3451
rect 9401 3411 9459 3417
rect 10137 3451 10195 3457
rect 10137 3417 10149 3451
rect 10183 3448 10195 3451
rect 11149 3451 11207 3457
rect 11149 3448 11161 3451
rect 10183 3420 11161 3448
rect 10183 3417 10195 3420
rect 10137 3411 10195 3417
rect 11149 3417 11161 3420
rect 11195 3448 11207 3451
rect 11624 3448 11652 3479
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 11195 3420 11652 3448
rect 11195 3417 11207 3420
rect 11149 3411 11207 3417
rect 9416 3380 9444 3411
rect 10226 3380 10232 3392
rect 9416 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3380 10290 3392
rect 10962 3380 10968 3392
rect 10284 3352 10968 3380
rect 10284 3340 10290 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11054 3340 11060 3392
rect 11112 3340 11118 3392
rect 12176 3380 12204 3556
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 12621 3587 12679 3593
rect 12621 3584 12633 3587
rect 12400 3556 12633 3584
rect 12400 3544 12406 3556
rect 12621 3553 12633 3556
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 13004 3535 13032 3624
rect 13354 3612 13360 3664
rect 13412 3652 13418 3664
rect 13449 3655 13507 3661
rect 13449 3652 13461 3655
rect 13412 3624 13461 3652
rect 13412 3612 13418 3624
rect 13449 3621 13461 3624
rect 13495 3621 13507 3655
rect 13449 3615 13507 3621
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3652 14703 3655
rect 14918 3652 14924 3664
rect 14691 3624 14924 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 15856 3652 15884 3692
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 18782 3720 18788 3732
rect 18739 3692 18788 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 18874 3680 18880 3732
rect 18932 3680 18938 3732
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22186 3720 22192 3732
rect 22143 3692 22192 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22186 3680 22192 3692
rect 22244 3720 22250 3732
rect 22830 3720 22836 3732
rect 22244 3692 22836 3720
rect 22244 3680 22250 3692
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 22922 3680 22928 3732
rect 22980 3680 22986 3732
rect 23934 3680 23940 3732
rect 23992 3720 23998 3732
rect 24486 3720 24492 3732
rect 23992 3692 24492 3720
rect 23992 3680 23998 3692
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 24854 3680 24860 3732
rect 24912 3680 24918 3732
rect 26145 3723 26203 3729
rect 26145 3689 26157 3723
rect 26191 3720 26203 3723
rect 28721 3723 28779 3729
rect 26191 3692 28304 3720
rect 26191 3689 26203 3692
rect 26145 3683 26203 3689
rect 15028 3624 15884 3652
rect 16301 3655 16359 3661
rect 15028 3584 15056 3624
rect 16301 3621 16313 3655
rect 16347 3652 16359 3655
rect 16347 3624 16436 3652
rect 16347 3621 16359 3624
rect 16301 3615 16359 3621
rect 16408 3593 16436 3624
rect 13376 3556 15056 3584
rect 15197 3587 15255 3593
rect 12994 3529 13052 3535
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12584 3488 12909 3516
rect 12584 3476 12590 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 12994 3495 13006 3529
rect 13040 3495 13052 3529
rect 13376 3528 13404 3556
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 15243 3556 15393 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 15381 3553 15393 3556
rect 15427 3584 15439 3587
rect 16117 3587 16175 3593
rect 16117 3584 16129 3587
rect 15427 3556 16129 3584
rect 15427 3553 15439 3556
rect 15381 3547 15439 3553
rect 16117 3553 16129 3556
rect 16163 3553 16175 3587
rect 16117 3547 16175 3553
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 17037 3587 17095 3593
rect 17037 3584 17049 3587
rect 16540 3556 17049 3584
rect 16540 3544 16546 3556
rect 17037 3553 17049 3556
rect 17083 3553 17095 3587
rect 17037 3547 17095 3553
rect 17310 3544 17316 3596
rect 17368 3544 17374 3596
rect 17451 3587 17509 3593
rect 17451 3553 17463 3587
rect 17497 3584 17509 3587
rect 18892 3584 18920 3680
rect 22462 3612 22468 3664
rect 22520 3612 22526 3664
rect 22741 3655 22799 3661
rect 22741 3621 22753 3655
rect 22787 3652 22799 3655
rect 22940 3652 22968 3680
rect 22787 3624 22968 3652
rect 22787 3621 22799 3624
rect 22741 3615 22799 3621
rect 23566 3612 23572 3664
rect 23624 3612 23630 3664
rect 24872 3652 24900 3680
rect 23952 3624 24900 3652
rect 28276 3652 28304 3692
rect 28721 3689 28733 3723
rect 28767 3720 28779 3723
rect 28994 3720 29000 3732
rect 28767 3692 29000 3720
rect 28767 3689 28779 3692
rect 28721 3683 28779 3689
rect 28994 3680 29000 3692
rect 29052 3680 29058 3732
rect 29454 3680 29460 3732
rect 29512 3680 29518 3732
rect 36265 3723 36323 3729
rect 36265 3689 36277 3723
rect 36311 3720 36323 3723
rect 36814 3720 36820 3732
rect 36311 3692 36820 3720
rect 36311 3689 36323 3692
rect 36265 3683 36323 3689
rect 36814 3680 36820 3692
rect 36872 3680 36878 3732
rect 29472 3652 29500 3680
rect 28276 3624 29500 3652
rect 17497 3556 18920 3584
rect 17497 3553 17509 3556
rect 17451 3547 17509 3553
rect 20162 3544 20168 3596
rect 20220 3584 20226 3596
rect 20349 3587 20407 3593
rect 20349 3584 20361 3587
rect 20220 3556 20361 3584
rect 20220 3544 20226 3556
rect 20349 3553 20361 3556
rect 20395 3553 20407 3587
rect 20349 3547 20407 3553
rect 20717 3587 20775 3593
rect 20717 3553 20729 3587
rect 20763 3584 20775 3587
rect 22281 3587 22339 3593
rect 22281 3584 22293 3587
rect 20763 3556 22293 3584
rect 20763 3553 20775 3556
rect 20717 3547 20775 3553
rect 22281 3553 22293 3556
rect 22327 3553 22339 3587
rect 22480 3584 22508 3612
rect 23584 3584 23612 3612
rect 22480 3556 22600 3584
rect 22281 3547 22339 3553
rect 13354 3503 13360 3528
rect 12994 3489 13052 3495
rect 13345 3497 13360 3503
rect 12897 3479 12955 3485
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 12621 3451 12679 3457
rect 12621 3448 12633 3451
rect 12308 3420 12633 3448
rect 12308 3408 12314 3420
rect 12621 3417 12633 3420
rect 12667 3417 12679 3451
rect 12621 3411 12679 3417
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12768 3420 12817 3448
rect 12768 3408 12774 3420
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 12912 3448 12940 3479
rect 13345 3463 13357 3497
rect 13412 3476 13418 3528
rect 13538 3476 13544 3528
rect 13596 3476 13602 3528
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13722 3516 13728 3528
rect 13679 3488 13728 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 14182 3516 14188 3528
rect 13863 3488 14188 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14608 3488 14749 3516
rect 14608 3476 14614 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 14884 3488 15577 3516
rect 14884 3476 14890 3488
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15565 3479 15623 3485
rect 15672 3488 15945 3516
rect 13391 3463 13403 3476
rect 13170 3448 13176 3460
rect 12912 3420 13176 3448
rect 12805 3411 12863 3417
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 13345 3457 13403 3463
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 13964 3420 14289 3448
rect 13964 3408 13970 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 14458 3408 14464 3460
rect 14516 3408 14522 3460
rect 15672 3380 15700 3488
rect 15933 3485 15945 3488
rect 15979 3516 15991 3519
rect 16206 3516 16212 3528
rect 15979 3488 16212 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 16316 3392 16344 3479
rect 16574 3476 16580 3528
rect 16632 3476 16638 3528
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18288 3488 18337 3516
rect 18288 3476 18294 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 18524 3448 18552 3479
rect 19242 3476 19248 3528
rect 19300 3476 19306 3528
rect 20806 3516 20812 3528
rect 19628 3488 20812 3516
rect 19628 3448 19656 3488
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 22462 3476 22468 3528
rect 22520 3476 22526 3528
rect 22572 3525 22600 3556
rect 22847 3556 23612 3584
rect 22847 3525 22875 3556
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3485 23167 3519
rect 23109 3479 23167 3485
rect 18064 3420 18552 3448
rect 18616 3420 19656 3448
rect 15746 3380 15752 3392
rect 12176 3352 15752 3380
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 16022 3340 16028 3392
rect 16080 3340 16086 3392
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 18064 3380 18092 3420
rect 16356 3352 18092 3380
rect 18233 3383 18291 3389
rect 16356 3340 16362 3352
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18616 3380 18644 3420
rect 20990 3408 20996 3460
rect 21048 3448 21054 3460
rect 21048 3420 21114 3448
rect 21048 3408 21054 3420
rect 22278 3408 22284 3460
rect 22336 3448 22342 3460
rect 23124 3448 23152 3479
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 23293 3519 23351 3525
rect 23293 3516 23305 3519
rect 23256 3488 23305 3516
rect 23256 3476 23262 3488
rect 23293 3485 23305 3488
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3516 23443 3519
rect 23952 3516 23980 3624
rect 24394 3544 24400 3596
rect 24452 3584 24458 3596
rect 26973 3587 27031 3593
rect 26973 3584 26985 3587
rect 24452 3556 26985 3584
rect 24452 3544 24458 3556
rect 26973 3553 26985 3556
rect 27019 3584 27031 3587
rect 27614 3584 27620 3596
rect 27019 3556 27620 3584
rect 27019 3553 27031 3556
rect 26973 3547 27031 3553
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 23431 3488 23980 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 22336 3420 23152 3448
rect 22336 3408 22342 3420
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 25516 3448 25544 3479
rect 26694 3476 26700 3528
rect 26752 3476 26758 3528
rect 36081 3519 36139 3525
rect 36081 3485 36093 3519
rect 36127 3516 36139 3519
rect 36538 3516 36544 3528
rect 36127 3488 36544 3516
rect 36127 3485 36139 3488
rect 36081 3479 36139 3485
rect 36538 3476 36544 3488
rect 36596 3476 36602 3528
rect 27249 3451 27307 3457
rect 27249 3448 27261 3451
rect 23532 3420 25544 3448
rect 26896 3420 27261 3448
rect 23532 3408 23538 3420
rect 18279 3352 18644 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 19426 3340 19432 3392
rect 19484 3340 19490 3392
rect 22554 3340 22560 3392
rect 22612 3380 22618 3392
rect 26896 3389 26924 3420
rect 27249 3417 27261 3420
rect 27295 3417 27307 3451
rect 27249 3411 27307 3417
rect 27522 3408 27528 3460
rect 27580 3448 27586 3460
rect 27580 3420 27738 3448
rect 27580 3408 27586 3420
rect 22925 3383 22983 3389
rect 22925 3380 22937 3383
rect 22612 3352 22937 3380
rect 22612 3340 22618 3352
rect 22925 3349 22937 3352
rect 22971 3349 22983 3383
rect 22925 3343 22983 3349
rect 26881 3383 26939 3389
rect 26881 3349 26893 3383
rect 26927 3349 26939 3383
rect 27632 3380 27660 3420
rect 29178 3380 29184 3392
rect 27632 3352 29184 3380
rect 26881 3343 26939 3349
rect 29178 3340 29184 3352
rect 29236 3340 29242 3392
rect 1104 3290 44620 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 44620 3290
rect 1104 3216 44620 3238
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 8251 3148 9260 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8754 3068 8760 3120
rect 8812 3068 8818 3120
rect 9232 3117 9260 3148
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 11514 3176 11520 3188
rect 9548 3148 10824 3176
rect 9548 3136 9554 3148
rect 9217 3111 9275 3117
rect 9217 3077 9229 3111
rect 9263 3077 9275 3111
rect 9217 3071 9275 3077
rect 9306 3068 9312 3120
rect 9364 3108 9370 3120
rect 9364 3080 9706 3108
rect 9364 3068 9370 3080
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 8036 2972 8064 3003
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 10796 3049 10824 3148
rect 11164 3148 11520 3176
rect 11164 3117 11192 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12710 3136 12716 3188
rect 12768 3136 12774 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 13906 3136 13912 3188
rect 13964 3136 13970 3188
rect 14734 3136 14740 3188
rect 14792 3136 14798 3188
rect 15657 3179 15715 3185
rect 15657 3145 15669 3179
rect 15703 3176 15715 3179
rect 16298 3176 16304 3188
rect 15703 3148 16304 3176
rect 15703 3145 15715 3148
rect 15657 3139 15715 3145
rect 11149 3111 11207 3117
rect 11149 3077 11161 3111
rect 11195 3077 11207 3111
rect 12986 3108 12992 3120
rect 11149 3071 11207 3077
rect 12728 3080 12992 3108
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8168 3012 8953 3040
rect 8168 3000 8174 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 10962 3000 10968 3052
rect 11020 3000 11026 3052
rect 12728 3049 12756 3080
rect 12986 3068 12992 3080
rect 13044 3108 13050 3120
rect 13372 3108 13400 3136
rect 13044 3080 13400 3108
rect 13044 3068 13050 3080
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3040 12955 3043
rect 13924 3040 13952 3136
rect 14752 3108 14780 3136
rect 14829 3111 14887 3117
rect 14829 3108 14841 3111
rect 14752 3080 14841 3108
rect 14829 3077 14841 3080
rect 14875 3077 14887 3111
rect 14829 3071 14887 3077
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 15672 3108 15700 3139
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16632 3148 16865 3176
rect 16632 3136 16638 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 19153 3179 19211 3185
rect 19153 3145 19165 3179
rect 19199 3176 19211 3179
rect 19242 3176 19248 3188
rect 19199 3148 19248 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 19334 3136 19340 3188
rect 19392 3136 19398 3188
rect 19426 3136 19432 3188
rect 19484 3136 19490 3188
rect 20162 3136 20168 3188
rect 20220 3136 20226 3188
rect 21453 3179 21511 3185
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 23474 3176 23480 3188
rect 21499 3148 22784 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 15059 3080 15700 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 16022 3068 16028 3120
rect 16080 3108 16086 3120
rect 19352 3108 19380 3136
rect 16080 3080 17356 3108
rect 16080 3068 16086 3080
rect 12943 3012 13952 3040
rect 15565 3043 15623 3049
rect 12943 3009 12955 3012
rect 12897 3003 12955 3009
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 15654 3040 15660 3052
rect 15611 3012 15660 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15746 3000 15752 3052
rect 15804 3000 15810 3052
rect 15930 3000 15936 3052
rect 15988 3040 15994 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 15988 3012 17049 3040
rect 15988 3000 15994 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17218 3000 17224 3052
rect 17276 3000 17282 3052
rect 17328 3049 17356 3080
rect 17420 3080 19380 3108
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8036 2944 8309 2972
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 13446 2932 13452 2984
rect 13504 2972 13510 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 13504 2944 15209 2972
rect 13504 2932 13510 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 17126 2972 17132 2984
rect 15528 2944 17132 2972
rect 15528 2932 15534 2944
rect 17126 2932 17132 2944
rect 17184 2932 17190 2984
rect 8481 2907 8539 2913
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 8662 2904 8668 2916
rect 8527 2876 8668 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 13170 2864 13176 2916
rect 13228 2904 13234 2916
rect 17420 2904 17448 3080
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 13228 2876 17448 2904
rect 13228 2864 13234 2876
rect 10686 2796 10692 2848
rect 10744 2796 10750 2848
rect 18708 2836 18736 3000
rect 19444 2972 19472 3136
rect 20180 3108 20208 3136
rect 19720 3080 20208 3108
rect 19720 3049 19748 3080
rect 20990 3068 20996 3120
rect 21048 3068 21054 3120
rect 22462 3068 22468 3120
rect 22520 3068 22526 3120
rect 22756 3108 22784 3148
rect 22940 3148 23480 3176
rect 22940 3108 22968 3148
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 23566 3136 23572 3188
rect 23624 3136 23630 3188
rect 24854 3136 24860 3188
rect 24912 3176 24918 3188
rect 30285 3179 30343 3185
rect 24912 3148 30144 3176
rect 24912 3136 24918 3148
rect 22756 3080 22968 3108
rect 23017 3111 23075 3117
rect 23017 3077 23029 3111
rect 23063 3108 23075 3111
rect 23584 3108 23612 3136
rect 23063 3080 23612 3108
rect 23063 3077 23075 3080
rect 23017 3071 23075 3077
rect 25406 3068 25412 3120
rect 25464 3068 25470 3120
rect 26050 3068 26056 3120
rect 26108 3108 26114 3120
rect 26513 3111 26571 3117
rect 26513 3108 26525 3111
rect 26108 3080 26525 3108
rect 26108 3068 26114 3080
rect 26513 3077 26525 3080
rect 26559 3077 26571 3111
rect 26513 3071 26571 3077
rect 29270 3068 29276 3120
rect 29328 3068 29334 3120
rect 30116 3108 30144 3148
rect 30285 3145 30297 3179
rect 30331 3176 30343 3179
rect 31202 3176 31208 3188
rect 30331 3148 31208 3176
rect 30331 3145 30343 3148
rect 30285 3139 30343 3145
rect 31202 3136 31208 3148
rect 31260 3136 31266 3188
rect 31726 3148 36124 3176
rect 31726 3108 31754 3148
rect 36096 3117 36124 3148
rect 36538 3136 36544 3188
rect 36596 3136 36602 3188
rect 30116 3080 31754 3108
rect 36081 3111 36139 3117
rect 36081 3077 36093 3111
rect 36127 3077 36139 3111
rect 36081 3071 36139 3077
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 22186 3000 22192 3052
rect 22244 3038 22250 3052
rect 22244 3010 22287 3038
rect 22244 3000 22250 3010
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 19444 2944 19993 2972
rect 19981 2941 19993 2944
rect 20027 2941 20039 2975
rect 19981 2935 20039 2941
rect 18966 2864 18972 2916
rect 19024 2864 19030 2916
rect 22480 2904 22508 3068
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22664 3012 22753 3040
rect 22664 2981 22692 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 22922 3040 22928 3052
rect 22879 3012 22928 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 23308 3012 23397 3040
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23017 2907 23075 2913
rect 23017 2904 23029 2907
rect 22066 2876 22416 2904
rect 22480 2876 23029 2904
rect 22066 2836 22094 2876
rect 18708 2808 22094 2836
rect 22278 2796 22284 2848
rect 22336 2796 22342 2848
rect 22388 2836 22416 2876
rect 23017 2873 23029 2876
rect 23063 2904 23075 2907
rect 23308 2904 23336 3012
rect 23385 3009 23397 3012
rect 23431 3009 23443 3043
rect 23385 3003 23443 3009
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 24452 3012 24501 3040
rect 24452 3000 24458 3012
rect 24489 3009 24501 3012
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 28537 3043 28595 3049
rect 28537 3040 28549 3043
rect 27672 3012 28549 3040
rect 27672 3000 27678 3012
rect 28537 3009 28549 3012
rect 28583 3009 28595 3043
rect 28537 3003 28595 3009
rect 23474 2932 23480 2984
rect 23532 2932 23538 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 23768 2944 24777 2972
rect 23768 2913 23796 2944
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 24765 2935 24823 2941
rect 28810 2932 28816 2984
rect 28868 2932 28874 2984
rect 23063 2876 23336 2904
rect 23753 2907 23811 2913
rect 23063 2873 23075 2876
rect 23017 2867 23075 2873
rect 23753 2873 23765 2907
rect 23799 2873 23811 2907
rect 23753 2867 23811 2873
rect 36449 2907 36507 2913
rect 36449 2873 36461 2907
rect 36495 2904 36507 2907
rect 43254 2904 43260 2916
rect 36495 2876 43260 2904
rect 36495 2873 36507 2876
rect 36449 2867 36507 2873
rect 43254 2864 43260 2876
rect 43312 2864 43318 2916
rect 24854 2836 24860 2848
rect 22388 2808 24860 2836
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 1104 2746 44620 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 44620 2746
rect 1104 2672 44620 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2038 2632 2044 2644
rect 1627 2604 2044 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 18966 2632 18972 2644
rect 17727 2604 18972 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 26053 2635 26111 2641
rect 26053 2601 26065 2635
rect 26099 2632 26111 2635
rect 26694 2632 26700 2644
rect 26099 2604 26700 2632
rect 26099 2601 26111 2604
rect 26053 2595 26111 2601
rect 26694 2592 26700 2604
rect 26752 2592 26758 2644
rect 43254 2592 43260 2644
rect 43312 2592 43318 2644
rect 25961 2567 26019 2573
rect 25961 2533 25973 2567
rect 26007 2564 26019 2567
rect 26145 2567 26203 2573
rect 26145 2564 26157 2567
rect 26007 2536 26157 2564
rect 26007 2533 26019 2536
rect 25961 2527 26019 2533
rect 26145 2533 26157 2536
rect 26191 2533 26203 2567
rect 26145 2527 26203 2533
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 19797 2499 19855 2505
rect 19797 2496 19809 2499
rect 10744 2468 19809 2496
rect 10744 2456 10750 2468
rect 19797 2465 19809 2468
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 20441 2499 20499 2505
rect 20441 2465 20453 2499
rect 20487 2496 20499 2499
rect 28810 2496 28816 2508
rect 20487 2468 28816 2496
rect 20487 2465 20499 2468
rect 20441 2459 20499 2465
rect 28810 2456 28816 2468
rect 28868 2456 28874 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 24912 2400 25605 2428
rect 24912 2388 24918 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26142 2388 26148 2440
rect 26200 2428 26206 2440
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 26200 2400 26341 2428
rect 26200 2388 26206 2400
rect 26329 2397 26341 2400
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 43220 2400 43453 2428
rect 43220 2388 43226 2400
rect 43441 2397 43453 2400
rect 43487 2397 43499 2431
rect 43441 2391 43499 2397
rect 1104 2202 44620 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 44620 2202
rect 1104 2128 44620 2150
<< via1 >>
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 14832 45500 14884 45552
rect 32220 45500 32272 45552
rect 1400 45475 1452 45484
rect 1400 45441 1409 45475
rect 1409 45441 1443 45475
rect 1443 45441 1452 45475
rect 1400 45432 1452 45441
rect 6460 45432 6512 45484
rect 23940 45475 23992 45484
rect 23940 45441 23949 45475
rect 23949 45441 23983 45475
rect 23983 45441 23992 45475
rect 23940 45432 23992 45441
rect 41236 45432 41288 45484
rect 5908 45228 5960 45280
rect 7288 45228 7340 45280
rect 15108 45271 15160 45280
rect 15108 45237 15117 45271
rect 15117 45237 15151 45271
rect 15151 45237 15160 45271
rect 15108 45228 15160 45237
rect 24308 45228 24360 45280
rect 32312 45271 32364 45280
rect 32312 45237 32321 45271
rect 32321 45237 32355 45271
rect 32355 45237 32364 45271
rect 32312 45228 32364 45237
rect 41328 45271 41380 45280
rect 41328 45237 41337 45271
rect 41337 45237 41371 45271
rect 41371 45237 41380 45271
rect 41328 45228 41380 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 15108 45024 15160 45076
rect 5908 44999 5960 45008
rect 5908 44965 5917 44999
rect 5917 44965 5951 44999
rect 5951 44965 5960 44999
rect 5908 44956 5960 44965
rect 6644 44888 6696 44940
rect 16120 44956 16172 45008
rect 32312 45024 32364 45076
rect 41328 45024 41380 45076
rect 16488 44888 16540 44940
rect 9864 44820 9916 44872
rect 12440 44820 12492 44872
rect 14096 44820 14148 44872
rect 15844 44863 15896 44872
rect 15844 44829 15853 44863
rect 15853 44829 15887 44863
rect 15887 44829 15896 44863
rect 15844 44820 15896 44829
rect 16028 44820 16080 44872
rect 16120 44863 16172 44872
rect 16120 44829 16129 44863
rect 16129 44829 16163 44863
rect 16163 44829 16172 44863
rect 16120 44820 16172 44829
rect 10508 44795 10560 44804
rect 10508 44761 10517 44795
rect 10517 44761 10551 44795
rect 10551 44761 10560 44795
rect 10508 44752 10560 44761
rect 11796 44752 11848 44804
rect 6092 44727 6144 44736
rect 6092 44693 6101 44727
rect 6101 44693 6135 44727
rect 6135 44693 6144 44727
rect 6092 44684 6144 44693
rect 12072 44727 12124 44736
rect 12072 44693 12081 44727
rect 12081 44693 12115 44727
rect 12115 44693 12124 44727
rect 12072 44684 12124 44693
rect 13452 44727 13504 44736
rect 13452 44693 13461 44727
rect 13461 44693 13495 44727
rect 13495 44693 13504 44727
rect 13452 44684 13504 44693
rect 14648 44684 14700 44736
rect 16028 44727 16080 44736
rect 16028 44693 16037 44727
rect 16037 44693 16071 44727
rect 16071 44693 16080 44727
rect 16028 44684 16080 44693
rect 16856 44752 16908 44804
rect 17868 44727 17920 44736
rect 17868 44693 17877 44727
rect 17877 44693 17911 44727
rect 17911 44693 17920 44727
rect 17868 44684 17920 44693
rect 37004 44752 37056 44804
rect 19156 44684 19208 44736
rect 19984 44684 20036 44736
rect 32036 44727 32088 44736
rect 32036 44693 32045 44727
rect 32045 44693 32079 44727
rect 32079 44693 32088 44727
rect 32036 44684 32088 44693
rect 36912 44727 36964 44736
rect 36912 44693 36921 44727
rect 36921 44693 36955 44727
rect 36955 44693 36964 44727
rect 36912 44684 36964 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 6092 44480 6144 44532
rect 10508 44480 10560 44532
rect 12072 44480 12124 44532
rect 13452 44480 13504 44532
rect 15844 44480 15896 44532
rect 19984 44480 20036 44532
rect 7288 44344 7340 44396
rect 6920 44140 6972 44192
rect 8208 44183 8260 44192
rect 8208 44149 8217 44183
rect 8217 44149 8251 44183
rect 8251 44149 8260 44183
rect 8208 44140 8260 44149
rect 11796 44140 11848 44192
rect 20076 44412 20128 44464
rect 32036 44480 32088 44532
rect 36912 44480 36964 44532
rect 20628 44412 20680 44464
rect 14648 44344 14700 44396
rect 17868 44344 17920 44396
rect 18512 44344 18564 44396
rect 11980 44319 12032 44328
rect 11980 44285 11989 44319
rect 11989 44285 12023 44319
rect 12023 44285 12032 44319
rect 11980 44276 12032 44285
rect 12072 44319 12124 44328
rect 12072 44285 12081 44319
rect 12081 44285 12115 44319
rect 12115 44285 12124 44319
rect 12072 44276 12124 44285
rect 12900 44319 12952 44328
rect 12900 44285 12909 44319
rect 12909 44285 12943 44319
rect 12943 44285 12952 44319
rect 12900 44276 12952 44285
rect 13084 44319 13136 44328
rect 13084 44285 13093 44319
rect 13093 44285 13127 44319
rect 13127 44285 13136 44319
rect 13084 44276 13136 44285
rect 14924 44276 14976 44328
rect 17132 44319 17184 44328
rect 17132 44285 17141 44319
rect 17141 44285 17175 44319
rect 17175 44285 17184 44319
rect 17132 44276 17184 44285
rect 17316 44319 17368 44328
rect 17316 44285 17325 44319
rect 17325 44285 17359 44319
rect 17359 44285 17368 44319
rect 17316 44276 17368 44285
rect 17960 44276 18012 44328
rect 19156 44344 19208 44396
rect 19432 44276 19484 44328
rect 27344 44276 27396 44328
rect 14464 44140 14516 44192
rect 18604 44183 18656 44192
rect 18604 44149 18613 44183
rect 18613 44149 18647 44183
rect 18647 44149 18656 44183
rect 18604 44140 18656 44149
rect 20628 44140 20680 44192
rect 25412 44140 25464 44192
rect 31668 44183 31720 44192
rect 31668 44149 31677 44183
rect 31677 44149 31711 44183
rect 31711 44149 31720 44183
rect 31668 44140 31720 44149
rect 36360 44140 36412 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 12900 43936 12952 43988
rect 14096 43979 14148 43988
rect 14096 43945 14105 43979
rect 14105 43945 14139 43979
rect 14139 43945 14148 43979
rect 14096 43936 14148 43945
rect 14188 43868 14240 43920
rect 7012 43800 7064 43852
rect 8208 43800 8260 43852
rect 6920 43664 6972 43716
rect 12072 43800 12124 43852
rect 17132 43936 17184 43988
rect 17776 43979 17828 43988
rect 17776 43945 17785 43979
rect 17785 43945 17819 43979
rect 17819 43945 17828 43979
rect 17776 43936 17828 43945
rect 17316 43868 17368 43920
rect 20536 43936 20588 43988
rect 16120 43800 16172 43852
rect 18604 43800 18656 43852
rect 20076 43800 20128 43852
rect 25412 43843 25464 43852
rect 25412 43809 25421 43843
rect 25421 43809 25455 43843
rect 25455 43809 25464 43843
rect 25412 43800 25464 43809
rect 31668 43800 31720 43852
rect 36360 43843 36412 43852
rect 36360 43809 36369 43843
rect 36369 43809 36403 43843
rect 36403 43809 36412 43843
rect 36360 43800 36412 43809
rect 9864 43732 9916 43784
rect 13176 43775 13228 43784
rect 13176 43741 13185 43775
rect 13185 43741 13219 43775
rect 13219 43741 13228 43775
rect 13176 43732 13228 43741
rect 13912 43775 13964 43784
rect 13912 43741 13921 43775
rect 13921 43741 13955 43775
rect 13955 43741 13964 43775
rect 13912 43732 13964 43741
rect 14464 43775 14516 43784
rect 14464 43741 14473 43775
rect 14473 43741 14507 43775
rect 14507 43741 14516 43775
rect 14464 43732 14516 43741
rect 14924 43775 14976 43784
rect 14924 43741 14933 43775
rect 14933 43741 14967 43775
rect 14967 43741 14976 43775
rect 14924 43732 14976 43741
rect 16856 43732 16908 43784
rect 19064 43732 19116 43784
rect 19248 43775 19300 43784
rect 19248 43741 19257 43775
rect 19257 43741 19291 43775
rect 19291 43741 19300 43775
rect 19248 43732 19300 43741
rect 20628 43732 20680 43784
rect 20812 43732 20864 43784
rect 31208 43732 31260 43784
rect 36084 43775 36136 43784
rect 36084 43741 36093 43775
rect 36093 43741 36127 43775
rect 36127 43741 36136 43775
rect 36084 43732 36136 43741
rect 8484 43639 8536 43648
rect 8484 43605 8493 43639
rect 8493 43605 8527 43639
rect 8527 43605 8536 43639
rect 8484 43596 8536 43605
rect 10876 43707 10928 43716
rect 10876 43673 10885 43707
rect 10885 43673 10919 43707
rect 10919 43673 10928 43707
rect 10876 43664 10928 43673
rect 15568 43707 15620 43716
rect 15568 43673 15577 43707
rect 15577 43673 15611 43707
rect 15611 43673 15620 43707
rect 15568 43664 15620 43673
rect 10968 43596 11020 43648
rect 12532 43639 12584 43648
rect 12532 43605 12541 43639
rect 12541 43605 12575 43639
rect 12575 43605 12584 43639
rect 12532 43596 12584 43605
rect 13820 43596 13872 43648
rect 32588 43664 32640 43716
rect 36820 43664 36872 43716
rect 43444 43707 43496 43716
rect 43444 43673 43453 43707
rect 43453 43673 43487 43707
rect 43487 43673 43496 43707
rect 43444 43664 43496 43673
rect 44640 43664 44692 43716
rect 18420 43639 18472 43648
rect 18420 43605 18429 43639
rect 18429 43605 18463 43639
rect 18463 43605 18472 43639
rect 18420 43596 18472 43605
rect 20996 43639 21048 43648
rect 20996 43605 21005 43639
rect 21005 43605 21039 43639
rect 21039 43605 21048 43639
rect 20996 43596 21048 43605
rect 29184 43596 29236 43648
rect 33048 43639 33100 43648
rect 33048 43605 33057 43639
rect 33057 43605 33091 43639
rect 33091 43605 33100 43639
rect 33048 43596 33100 43605
rect 37832 43639 37884 43648
rect 37832 43605 37841 43639
rect 37841 43605 37875 43639
rect 37875 43605 37884 43639
rect 37832 43596 37884 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 10876 43392 10928 43444
rect 12532 43392 12584 43444
rect 13912 43392 13964 43444
rect 15568 43392 15620 43444
rect 17776 43392 17828 43444
rect 11980 43324 12032 43376
rect 20996 43392 21048 43444
rect 20812 43324 20864 43376
rect 10876 43299 10928 43308
rect 10876 43265 10885 43299
rect 10885 43265 10919 43299
rect 10919 43265 10928 43299
rect 10876 43256 10928 43265
rect 12440 43299 12492 43308
rect 12440 43265 12449 43299
rect 12449 43265 12483 43299
rect 12483 43265 12492 43299
rect 12440 43256 12492 43265
rect 14648 43256 14700 43308
rect 16120 43256 16172 43308
rect 12624 43188 12676 43240
rect 12532 43095 12584 43104
rect 12532 43061 12541 43095
rect 12541 43061 12575 43095
rect 12575 43061 12584 43095
rect 12532 43052 12584 43061
rect 14832 43188 14884 43240
rect 17316 43231 17368 43240
rect 17316 43197 17325 43231
rect 17325 43197 17359 43231
rect 17359 43197 17368 43231
rect 17316 43188 17368 43197
rect 17684 43299 17736 43308
rect 17684 43265 17693 43299
rect 17693 43265 17727 43299
rect 17727 43265 17736 43299
rect 17684 43256 17736 43265
rect 17960 43299 18012 43308
rect 17960 43265 17969 43299
rect 17969 43265 18003 43299
rect 18003 43265 18012 43299
rect 17960 43256 18012 43265
rect 20628 43256 20680 43308
rect 31208 43392 31260 43444
rect 33048 43392 33100 43444
rect 29184 43367 29236 43376
rect 29184 43333 29193 43367
rect 29193 43333 29227 43367
rect 29227 43333 29236 43367
rect 29184 43324 29236 43333
rect 18144 43231 18196 43240
rect 18144 43197 18153 43231
rect 18153 43197 18187 43231
rect 18187 43197 18196 43231
rect 18144 43188 18196 43197
rect 18420 43231 18472 43240
rect 18420 43197 18429 43231
rect 18429 43197 18463 43231
rect 18463 43197 18472 43231
rect 18420 43188 18472 43197
rect 19064 43188 19116 43240
rect 20076 43188 20128 43240
rect 20536 43231 20588 43240
rect 20536 43197 20545 43231
rect 20545 43197 20579 43231
rect 20579 43197 20588 43231
rect 20536 43188 20588 43197
rect 24032 43231 24084 43240
rect 24032 43197 24041 43231
rect 24041 43197 24075 43231
rect 24075 43197 24084 43231
rect 24032 43188 24084 43197
rect 27160 43188 27212 43240
rect 32588 43256 32640 43308
rect 40592 43324 40644 43376
rect 36452 43188 36504 43240
rect 38660 43188 38712 43240
rect 39212 43231 39264 43240
rect 39212 43197 39221 43231
rect 39221 43197 39255 43231
rect 39255 43197 39264 43231
rect 39212 43188 39264 43197
rect 13084 43052 13136 43104
rect 15016 43095 15068 43104
rect 15016 43061 15025 43095
rect 15025 43061 15059 43095
rect 15059 43061 15068 43095
rect 15016 43052 15068 43061
rect 16764 43095 16816 43104
rect 16764 43061 16773 43095
rect 16773 43061 16807 43095
rect 16807 43061 16816 43095
rect 16764 43052 16816 43061
rect 17224 43052 17276 43104
rect 24308 43163 24360 43172
rect 24308 43129 24317 43163
rect 24317 43129 24351 43163
rect 24351 43129 24360 43163
rect 24308 43120 24360 43129
rect 21456 43052 21508 43104
rect 24860 43052 24912 43104
rect 31300 43052 31352 43104
rect 34060 43095 34112 43104
rect 34060 43061 34069 43095
rect 34069 43061 34103 43095
rect 34103 43061 34112 43095
rect 34060 43052 34112 43061
rect 35532 43095 35584 43104
rect 35532 43061 35541 43095
rect 35541 43061 35575 43095
rect 35575 43061 35584 43095
rect 35532 43052 35584 43061
rect 40684 43095 40736 43104
rect 40684 43061 40693 43095
rect 40693 43061 40727 43095
rect 40727 43061 40736 43095
rect 40684 43052 40736 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 12624 42848 12676 42900
rect 13176 42848 13228 42900
rect 17316 42848 17368 42900
rect 18144 42848 18196 42900
rect 6644 42755 6696 42764
rect 6644 42721 6653 42755
rect 6653 42721 6687 42755
rect 6687 42721 6696 42755
rect 6644 42712 6696 42721
rect 5540 42644 5592 42696
rect 17224 42780 17276 42832
rect 24032 42848 24084 42900
rect 39212 42848 39264 42900
rect 43444 42848 43496 42900
rect 8852 42576 8904 42628
rect 10140 42644 10192 42696
rect 10968 42687 11020 42696
rect 10968 42653 10977 42687
rect 10977 42653 11011 42687
rect 11011 42653 11020 42687
rect 10968 42644 11020 42653
rect 11980 42644 12032 42696
rect 14556 42712 14608 42764
rect 14648 42712 14700 42764
rect 8944 42551 8996 42560
rect 8944 42517 8953 42551
rect 8953 42517 8987 42551
rect 8987 42517 8996 42551
rect 8944 42508 8996 42517
rect 9496 42508 9548 42560
rect 10048 42508 10100 42560
rect 13820 42687 13872 42696
rect 13820 42653 13829 42687
rect 13829 42653 13863 42687
rect 13863 42653 13872 42687
rect 13820 42644 13872 42653
rect 13912 42687 13964 42696
rect 13912 42653 13921 42687
rect 13921 42653 13955 42687
rect 13955 42653 13964 42687
rect 13912 42644 13964 42653
rect 14004 42644 14056 42696
rect 15200 42619 15252 42628
rect 15200 42585 15209 42619
rect 15209 42585 15243 42619
rect 15243 42585 15252 42619
rect 15200 42576 15252 42585
rect 18604 42755 18656 42764
rect 18604 42721 18613 42755
rect 18613 42721 18647 42755
rect 18647 42721 18656 42755
rect 19248 42755 19300 42764
rect 18604 42712 18656 42721
rect 19248 42721 19257 42755
rect 19257 42721 19291 42755
rect 19291 42721 19300 42755
rect 19248 42712 19300 42721
rect 38844 42755 38896 42764
rect 38844 42721 38853 42755
rect 38853 42721 38887 42755
rect 38887 42721 38896 42755
rect 38844 42712 38896 42721
rect 40684 42712 40736 42764
rect 16856 42644 16908 42696
rect 18328 42619 18380 42628
rect 18328 42585 18337 42619
rect 18337 42585 18371 42619
rect 18371 42585 18380 42619
rect 18328 42576 18380 42585
rect 14096 42508 14148 42560
rect 14924 42508 14976 42560
rect 17040 42508 17092 42560
rect 24860 42644 24912 42696
rect 20996 42619 21048 42628
rect 20996 42585 21005 42619
rect 21005 42585 21039 42619
rect 21039 42585 21048 42619
rect 20996 42576 21048 42585
rect 36820 42644 36872 42696
rect 37096 42644 37148 42696
rect 40776 42687 40828 42696
rect 40776 42653 40785 42687
rect 40785 42653 40819 42687
rect 40819 42653 40828 42687
rect 40776 42644 40828 42653
rect 34980 42619 35032 42628
rect 34980 42585 34989 42619
rect 34989 42585 35023 42619
rect 35023 42585 35032 42619
rect 34980 42576 35032 42585
rect 19156 42508 19208 42560
rect 25136 42551 25188 42560
rect 25136 42517 25145 42551
rect 25145 42517 25179 42551
rect 25179 42517 25188 42551
rect 25136 42508 25188 42517
rect 34796 42508 34848 42560
rect 36452 42551 36504 42560
rect 36452 42517 36461 42551
rect 36461 42517 36495 42551
rect 36495 42517 36504 42551
rect 36452 42508 36504 42517
rect 36912 42508 36964 42560
rect 40316 42508 40368 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 7012 42168 7064 42220
rect 8852 42236 8904 42288
rect 7380 42143 7432 42152
rect 7380 42109 7389 42143
rect 7389 42109 7423 42143
rect 7423 42109 7432 42143
rect 7380 42100 7432 42109
rect 9864 42304 9916 42356
rect 10968 42304 11020 42356
rect 9496 42236 9548 42288
rect 11796 42236 11848 42288
rect 13268 42236 13320 42288
rect 14648 42236 14700 42288
rect 14832 42347 14884 42356
rect 14832 42313 14841 42347
rect 14841 42313 14875 42347
rect 14875 42313 14884 42347
rect 14832 42304 14884 42313
rect 15200 42304 15252 42356
rect 16672 42304 16724 42356
rect 17684 42304 17736 42356
rect 18328 42304 18380 42356
rect 18420 42304 18472 42356
rect 14924 42211 14976 42220
rect 14924 42177 14933 42211
rect 14933 42177 14967 42211
rect 14967 42177 14976 42211
rect 14924 42168 14976 42177
rect 15016 42211 15068 42220
rect 15016 42177 15026 42211
rect 15026 42177 15060 42211
rect 15060 42177 15068 42211
rect 16764 42236 16816 42288
rect 15016 42168 15068 42177
rect 15568 42168 15620 42220
rect 11244 42100 11296 42152
rect 12164 42143 12216 42152
rect 12164 42109 12173 42143
rect 12173 42109 12207 42143
rect 12207 42109 12216 42143
rect 12164 42100 12216 42109
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 11980 41964 12032 42016
rect 13084 42143 13136 42152
rect 13084 42109 13093 42143
rect 13093 42109 13127 42143
rect 13127 42109 13136 42143
rect 13084 42100 13136 42109
rect 13360 42143 13412 42152
rect 13360 42109 13369 42143
rect 13369 42109 13403 42143
rect 13403 42109 13412 42143
rect 13360 42100 13412 42109
rect 14096 42100 14148 42152
rect 14464 42032 14516 42084
rect 14556 42032 14608 42084
rect 17408 42168 17460 42220
rect 19156 42304 19208 42356
rect 19248 42304 19300 42356
rect 20352 42304 20404 42356
rect 17316 42143 17368 42152
rect 17316 42109 17325 42143
rect 17325 42109 17359 42143
rect 17359 42109 17368 42143
rect 17316 42100 17368 42109
rect 18788 42211 18840 42220
rect 18788 42177 18802 42211
rect 18802 42177 18836 42211
rect 18836 42177 18840 42211
rect 18788 42168 18840 42177
rect 20628 42168 20680 42220
rect 25136 42304 25188 42356
rect 22376 42236 22428 42288
rect 27160 42347 27212 42356
rect 27160 42313 27169 42347
rect 27169 42313 27203 42347
rect 27203 42313 27212 42347
rect 27160 42304 27212 42313
rect 27436 42236 27488 42288
rect 34060 42304 34112 42356
rect 18144 42032 18196 42084
rect 14004 41964 14056 42016
rect 17960 41964 18012 42016
rect 18972 42007 19024 42016
rect 18972 41973 18981 42007
rect 18981 41973 19015 42007
rect 19015 41973 19024 42007
rect 18972 41964 19024 41973
rect 19340 42143 19392 42152
rect 19340 42109 19349 42143
rect 19349 42109 19383 42143
rect 19383 42109 19392 42143
rect 19340 42100 19392 42109
rect 22100 42143 22152 42152
rect 22100 42109 22109 42143
rect 22109 42109 22143 42143
rect 22143 42109 22152 42143
rect 22100 42100 22152 42109
rect 24400 42100 24452 42152
rect 26884 42100 26936 42152
rect 27344 42211 27396 42220
rect 27344 42177 27353 42211
rect 27353 42177 27387 42211
rect 27387 42177 27396 42211
rect 27344 42168 27396 42177
rect 32588 42168 32640 42220
rect 34796 42236 34848 42288
rect 35532 42304 35584 42356
rect 38844 42347 38896 42356
rect 38844 42313 38853 42347
rect 38853 42313 38887 42347
rect 38887 42313 38896 42347
rect 38844 42304 38896 42313
rect 36176 42236 36228 42288
rect 36912 42279 36964 42288
rect 36912 42245 36921 42279
rect 36921 42245 36955 42279
rect 36955 42245 36964 42279
rect 36912 42236 36964 42245
rect 40316 42304 40368 42356
rect 40592 42236 40644 42288
rect 34704 42143 34756 42152
rect 34704 42109 34713 42143
rect 34713 42109 34747 42143
rect 34747 42109 34756 42143
rect 34704 42100 34756 42109
rect 34980 42143 35032 42152
rect 34980 42109 34989 42143
rect 34989 42109 35023 42143
rect 35023 42109 35032 42143
rect 34980 42100 35032 42109
rect 35716 42168 35768 42220
rect 35532 42100 35584 42152
rect 35624 42032 35676 42084
rect 20904 42007 20956 42016
rect 20904 41973 20913 42007
rect 20913 41973 20947 42007
rect 20947 41973 20956 42007
rect 20904 41964 20956 41973
rect 23572 42007 23624 42016
rect 23572 41973 23581 42007
rect 23581 41973 23615 42007
rect 23615 41973 23624 42007
rect 23572 41964 23624 41973
rect 27068 41964 27120 42016
rect 30932 41964 30984 42016
rect 36452 42007 36504 42016
rect 36452 41973 36461 42007
rect 36461 41973 36495 42007
rect 36495 41973 36504 42007
rect 36452 41964 36504 41973
rect 36544 42007 36596 42016
rect 36544 41973 36553 42007
rect 36553 41973 36587 42007
rect 36587 41973 36596 42007
rect 36544 41964 36596 41973
rect 36728 42007 36780 42016
rect 36728 41973 36737 42007
rect 36737 41973 36771 42007
rect 36771 41973 36780 42007
rect 36728 41964 36780 41973
rect 38844 42211 38896 42220
rect 38844 42177 38853 42211
rect 38853 42177 38887 42211
rect 38887 42177 38896 42211
rect 38844 42168 38896 42177
rect 39396 42168 39448 42220
rect 42248 42168 42300 42220
rect 38476 42100 38528 42152
rect 40592 42100 40644 42152
rect 41144 42100 41196 42152
rect 42432 42143 42484 42152
rect 42432 42109 42441 42143
rect 42441 42109 42475 42143
rect 42475 42109 42484 42143
rect 42432 42100 42484 42109
rect 41236 41964 41288 42016
rect 41604 42007 41656 42016
rect 41604 41973 41613 42007
rect 41613 41973 41647 42007
rect 41647 41973 41656 42007
rect 41604 41964 41656 41973
rect 42340 41964 42392 42016
rect 44180 42007 44232 42016
rect 44180 41973 44189 42007
rect 44189 41973 44223 42007
rect 44223 41973 44232 42007
rect 44180 41964 44232 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 7380 41760 7432 41812
rect 8944 41760 8996 41812
rect 10140 41803 10192 41812
rect 10140 41769 10149 41803
rect 10149 41769 10183 41803
rect 10183 41769 10192 41803
rect 10140 41760 10192 41769
rect 11980 41803 12032 41812
rect 11980 41769 11989 41803
rect 11989 41769 12023 41803
rect 12023 41769 12032 41803
rect 11980 41760 12032 41769
rect 12164 41760 12216 41812
rect 9588 41667 9640 41676
rect 9588 41633 9597 41667
rect 9597 41633 9631 41667
rect 9631 41633 9640 41667
rect 9588 41624 9640 41633
rect 9864 41624 9916 41676
rect 13360 41760 13412 41812
rect 15568 41760 15620 41812
rect 17316 41803 17368 41812
rect 17316 41769 17325 41803
rect 17325 41769 17359 41803
rect 17359 41769 17368 41803
rect 17316 41760 17368 41769
rect 18420 41760 18472 41812
rect 18972 41760 19024 41812
rect 19340 41760 19392 41812
rect 20904 41760 20956 41812
rect 22100 41760 22152 41812
rect 23572 41760 23624 41812
rect 31208 41760 31260 41812
rect 12900 41624 12952 41676
rect 10048 41556 10100 41608
rect 11796 41556 11848 41608
rect 11888 41556 11940 41608
rect 12624 41556 12676 41608
rect 8484 41463 8536 41472
rect 8484 41429 8493 41463
rect 8493 41429 8527 41463
rect 8527 41429 8536 41463
rect 8484 41420 8536 41429
rect 9680 41463 9732 41472
rect 9680 41429 9689 41463
rect 9689 41429 9723 41463
rect 9723 41429 9732 41463
rect 9680 41420 9732 41429
rect 10508 41531 10560 41540
rect 10508 41497 10517 41531
rect 10517 41497 10551 41531
rect 10551 41497 10560 41531
rect 10508 41488 10560 41497
rect 12532 41488 12584 41540
rect 15476 41556 15528 41608
rect 16672 41599 16724 41608
rect 16672 41565 16681 41599
rect 16681 41565 16715 41599
rect 16715 41565 16724 41599
rect 16672 41556 16724 41565
rect 16764 41599 16816 41608
rect 16764 41565 16774 41599
rect 16774 41565 16808 41599
rect 16808 41565 16816 41599
rect 16764 41556 16816 41565
rect 17040 41599 17092 41608
rect 17040 41565 17049 41599
rect 17049 41565 17083 41599
rect 17083 41565 17092 41599
rect 17040 41556 17092 41565
rect 18788 41624 18840 41676
rect 17592 41599 17644 41608
rect 17592 41565 17601 41599
rect 17601 41565 17635 41599
rect 17635 41565 17644 41599
rect 17592 41556 17644 41565
rect 13268 41531 13320 41540
rect 13268 41497 13277 41531
rect 13277 41497 13311 41531
rect 13311 41497 13320 41531
rect 13268 41488 13320 41497
rect 15016 41488 15068 41540
rect 18144 41488 18196 41540
rect 20812 41599 20864 41608
rect 20812 41565 20821 41599
rect 20821 41565 20855 41599
rect 20855 41565 20864 41599
rect 20812 41556 20864 41565
rect 24216 41556 24268 41608
rect 17316 41420 17368 41472
rect 17960 41420 18012 41472
rect 19432 41420 19484 41472
rect 23572 41488 23624 41540
rect 34704 41760 34756 41812
rect 35348 41760 35400 41812
rect 36084 41760 36136 41812
rect 37280 41760 37332 41812
rect 38476 41760 38528 41812
rect 38936 41760 38988 41812
rect 32036 41556 32088 41608
rect 33140 41556 33192 41608
rect 34520 41556 34572 41608
rect 35624 41556 35676 41608
rect 36084 41599 36136 41608
rect 36084 41565 36093 41599
rect 36093 41565 36127 41599
rect 36127 41565 36136 41599
rect 36084 41556 36136 41565
rect 34888 41488 34940 41540
rect 35900 41488 35952 41540
rect 36452 41556 36504 41608
rect 36544 41556 36596 41608
rect 38200 41599 38252 41608
rect 38200 41565 38209 41599
rect 38209 41565 38243 41599
rect 38243 41565 38252 41599
rect 38200 41556 38252 41565
rect 39948 41556 40000 41608
rect 40868 41760 40920 41812
rect 41236 41760 41288 41812
rect 40960 41692 41012 41744
rect 41604 41624 41656 41676
rect 42248 41803 42300 41812
rect 42248 41769 42257 41803
rect 42257 41769 42291 41803
rect 42291 41769 42300 41803
rect 42248 41760 42300 41769
rect 40868 41599 40920 41608
rect 40868 41565 40877 41599
rect 40877 41565 40911 41599
rect 40911 41565 40920 41599
rect 40868 41556 40920 41565
rect 40960 41599 41012 41608
rect 40960 41565 40969 41599
rect 40969 41565 41003 41599
rect 41003 41565 41012 41599
rect 40960 41556 41012 41565
rect 39488 41531 39540 41540
rect 39488 41497 39497 41531
rect 39497 41497 39531 41531
rect 39531 41497 39540 41531
rect 39488 41488 39540 41497
rect 22284 41420 22336 41472
rect 35440 41463 35492 41472
rect 35440 41429 35449 41463
rect 35449 41429 35483 41463
rect 35483 41429 35492 41463
rect 35440 41420 35492 41429
rect 36268 41463 36320 41472
rect 36268 41429 36277 41463
rect 36277 41429 36311 41463
rect 36311 41429 36320 41463
rect 36268 41420 36320 41429
rect 39120 41463 39172 41472
rect 39120 41429 39129 41463
rect 39129 41429 39163 41463
rect 39163 41429 39172 41463
rect 39120 41420 39172 41429
rect 39304 41463 39356 41472
rect 39304 41429 39331 41463
rect 39331 41429 39356 41463
rect 39304 41420 39356 41429
rect 39396 41420 39448 41472
rect 39948 41420 40000 41472
rect 40040 41463 40092 41472
rect 40040 41429 40049 41463
rect 40049 41429 40083 41463
rect 40083 41429 40092 41463
rect 40040 41420 40092 41429
rect 40316 41531 40368 41540
rect 40316 41497 40325 41531
rect 40325 41497 40359 41531
rect 40359 41497 40368 41531
rect 40316 41488 40368 41497
rect 40408 41531 40460 41540
rect 40408 41497 40417 41531
rect 40417 41497 40451 41531
rect 40451 41497 40460 41531
rect 40408 41488 40460 41497
rect 40684 41488 40736 41540
rect 41328 41488 41380 41540
rect 41788 41488 41840 41540
rect 42432 41624 42484 41676
rect 43352 41624 43404 41676
rect 43076 41488 43128 41540
rect 42064 41463 42116 41472
rect 42064 41429 42089 41463
rect 42089 41429 42116 41463
rect 42064 41420 42116 41429
rect 44088 41420 44140 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 10508 41216 10560 41268
rect 11888 41259 11940 41268
rect 11888 41225 11897 41259
rect 11897 41225 11931 41259
rect 11931 41225 11940 41259
rect 11888 41216 11940 41225
rect 10876 41080 10928 41132
rect 11520 41080 11572 41132
rect 14004 41012 14056 41064
rect 14280 41055 14332 41064
rect 14280 41021 14289 41055
rect 14289 41021 14323 41055
rect 14323 41021 14332 41055
rect 14280 41012 14332 41021
rect 15476 41055 15528 41064
rect 15476 41021 15485 41055
rect 15485 41021 15519 41055
rect 15519 41021 15528 41055
rect 15476 41012 15528 41021
rect 15568 41055 15620 41064
rect 15568 41021 15577 41055
rect 15577 41021 15611 41055
rect 15611 41021 15620 41055
rect 15568 41012 15620 41021
rect 17592 41080 17644 41132
rect 18144 41123 18196 41132
rect 18144 41089 18153 41123
rect 18153 41089 18187 41123
rect 18187 41089 18196 41123
rect 18144 41080 18196 41089
rect 20812 41216 20864 41268
rect 33140 41216 33192 41268
rect 34888 41216 34940 41268
rect 19432 41148 19484 41200
rect 22192 41148 22244 41200
rect 35716 41216 35768 41268
rect 36268 41216 36320 41268
rect 37096 41216 37148 41268
rect 17960 41055 18012 41064
rect 17960 41021 17969 41055
rect 17969 41021 18003 41055
rect 18003 41021 18012 41055
rect 17960 41012 18012 41021
rect 9864 40876 9916 40928
rect 13728 40876 13780 40928
rect 16120 40919 16172 40928
rect 16120 40885 16129 40919
rect 16129 40885 16163 40919
rect 16163 40885 16172 40919
rect 16120 40876 16172 40885
rect 19156 40919 19208 40928
rect 19156 40885 19165 40919
rect 19165 40885 19199 40919
rect 19199 40885 19208 40919
rect 19156 40876 19208 40885
rect 20444 41055 20496 41064
rect 20444 41021 20453 41055
rect 20453 41021 20487 41055
rect 20487 41021 20496 41055
rect 20444 41012 20496 41021
rect 22008 41080 22060 41132
rect 34612 41080 34664 41132
rect 22560 41012 22612 41064
rect 22928 41055 22980 41064
rect 22928 41021 22937 41055
rect 22937 41021 22971 41055
rect 22971 41021 22980 41055
rect 22928 41012 22980 41021
rect 34796 41012 34848 41064
rect 35348 41055 35400 41064
rect 35348 41021 35357 41055
rect 35357 41021 35391 41055
rect 35391 41021 35400 41055
rect 35348 41012 35400 41021
rect 36176 41012 36228 41064
rect 20076 40876 20128 40928
rect 23940 40919 23992 40928
rect 23940 40885 23949 40919
rect 23949 40885 23983 40919
rect 23983 40885 23992 40919
rect 23940 40876 23992 40885
rect 34888 40876 34940 40928
rect 36084 40876 36136 40928
rect 37280 41123 37332 41132
rect 37280 41089 37289 41123
rect 37289 41089 37323 41123
rect 37323 41089 37332 41123
rect 37280 41080 37332 41089
rect 37556 41055 37608 41064
rect 37556 41021 37565 41055
rect 37565 41021 37599 41055
rect 37599 41021 37608 41055
rect 37556 41012 37608 41021
rect 38844 41216 38896 41268
rect 39304 41216 39356 41268
rect 40776 41216 40828 41268
rect 42064 41259 42116 41268
rect 42064 41225 42073 41259
rect 42073 41225 42107 41259
rect 42107 41225 42116 41259
rect 42064 41216 42116 41225
rect 39396 41148 39448 41200
rect 40408 41148 40460 41200
rect 40960 41148 41012 41200
rect 40040 41123 40092 41132
rect 40040 41089 40049 41123
rect 40049 41089 40083 41123
rect 40083 41089 40092 41123
rect 40040 41080 40092 41089
rect 41328 41080 41380 41132
rect 42708 41148 42760 41200
rect 41144 41012 41196 41064
rect 41788 41012 41840 41064
rect 42340 41080 42392 41132
rect 42524 41012 42576 41064
rect 44180 41080 44232 41132
rect 41052 40944 41104 40996
rect 41880 40876 41932 40928
rect 42800 40919 42852 40928
rect 42800 40885 42809 40919
rect 42809 40885 42843 40919
rect 42843 40885 42852 40919
rect 42800 40876 42852 40885
rect 43168 40919 43220 40928
rect 43168 40885 43177 40919
rect 43177 40885 43211 40919
rect 43211 40885 43220 40919
rect 43168 40876 43220 40885
rect 43260 40876 43312 40928
rect 44088 40919 44140 40928
rect 44088 40885 44097 40919
rect 44097 40885 44131 40919
rect 44131 40885 44140 40919
rect 44088 40876 44140 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 14280 40672 14332 40724
rect 17592 40672 17644 40724
rect 17960 40672 18012 40724
rect 19156 40672 19208 40724
rect 21088 40672 21140 40724
rect 22928 40672 22980 40724
rect 23940 40672 23992 40724
rect 35532 40672 35584 40724
rect 36728 40715 36780 40724
rect 36728 40681 36737 40715
rect 36737 40681 36771 40715
rect 36771 40681 36780 40715
rect 36728 40672 36780 40681
rect 37556 40672 37608 40724
rect 40408 40672 40460 40724
rect 40684 40672 40736 40724
rect 42708 40672 42760 40724
rect 43168 40672 43220 40724
rect 43352 40715 43404 40724
rect 43352 40681 43361 40715
rect 43361 40681 43395 40715
rect 43395 40681 43404 40715
rect 43352 40672 43404 40681
rect 8484 40468 8536 40520
rect 9864 40536 9916 40588
rect 12256 40511 12308 40520
rect 12256 40477 12265 40511
rect 12265 40477 12299 40511
rect 12299 40477 12308 40511
rect 12256 40468 12308 40477
rect 16120 40536 16172 40588
rect 12900 40468 12952 40520
rect 13544 40511 13596 40520
rect 13544 40477 13553 40511
rect 13553 40477 13587 40511
rect 13587 40477 13596 40511
rect 13544 40468 13596 40477
rect 15108 40468 15160 40520
rect 16672 40468 16724 40520
rect 17408 40468 17460 40520
rect 17684 40511 17736 40520
rect 17684 40477 17693 40511
rect 17693 40477 17727 40511
rect 17727 40477 17736 40511
rect 17684 40468 17736 40477
rect 17960 40468 18012 40520
rect 18788 40511 18840 40520
rect 18788 40477 18797 40511
rect 18797 40477 18831 40511
rect 18831 40477 18840 40511
rect 18788 40468 18840 40477
rect 9404 40443 9456 40452
rect 9404 40409 9413 40443
rect 9413 40409 9447 40443
rect 9447 40409 9456 40443
rect 9404 40400 9456 40409
rect 10876 40400 10928 40452
rect 12532 40443 12584 40452
rect 12532 40409 12541 40443
rect 12541 40409 12575 40443
rect 12575 40409 12584 40443
rect 12532 40400 12584 40409
rect 8576 40332 8628 40384
rect 8760 40375 8812 40384
rect 8760 40341 8769 40375
rect 8769 40341 8803 40375
rect 8803 40341 8812 40375
rect 8760 40332 8812 40341
rect 9680 40332 9732 40384
rect 10784 40332 10836 40384
rect 10968 40332 11020 40384
rect 11888 40332 11940 40384
rect 16028 40400 16080 40452
rect 16856 40400 16908 40452
rect 20168 40400 20220 40452
rect 20352 40579 20404 40588
rect 20352 40545 20361 40579
rect 20361 40545 20395 40579
rect 20395 40545 20404 40579
rect 20352 40536 20404 40545
rect 20628 40536 20680 40588
rect 24400 40604 24452 40656
rect 22376 40468 22428 40520
rect 24124 40468 24176 40520
rect 34520 40468 34572 40520
rect 35256 40443 35308 40452
rect 35256 40409 35265 40443
rect 35265 40409 35299 40443
rect 35299 40409 35308 40443
rect 35256 40400 35308 40409
rect 35900 40468 35952 40520
rect 17224 40332 17276 40384
rect 19064 40332 19116 40384
rect 22100 40375 22152 40384
rect 22100 40341 22109 40375
rect 22109 40341 22143 40375
rect 22143 40341 22152 40375
rect 22100 40332 22152 40341
rect 24952 40332 25004 40384
rect 34612 40332 34664 40384
rect 35532 40332 35584 40384
rect 35992 40400 36044 40452
rect 36176 40400 36228 40452
rect 36912 40468 36964 40520
rect 39120 40468 39172 40520
rect 40592 40511 40644 40520
rect 40592 40477 40601 40511
rect 40601 40477 40635 40511
rect 40635 40477 40644 40511
rect 40592 40468 40644 40477
rect 42524 40468 42576 40520
rect 43260 40468 43312 40520
rect 37372 40332 37424 40384
rect 40132 40332 40184 40384
rect 40776 40375 40828 40384
rect 40776 40341 40785 40375
rect 40785 40341 40819 40375
rect 40819 40341 40828 40375
rect 40776 40332 40828 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 8576 40171 8628 40180
rect 8576 40137 8585 40171
rect 8585 40137 8619 40171
rect 8619 40137 8628 40171
rect 8576 40128 8628 40137
rect 8760 40128 8812 40180
rect 9404 40128 9456 40180
rect 12256 40128 12308 40180
rect 13728 40128 13780 40180
rect 19156 40128 19208 40180
rect 21088 40171 21140 40180
rect 21088 40137 21097 40171
rect 21097 40137 21131 40171
rect 21131 40137 21140 40171
rect 21088 40128 21140 40137
rect 9220 39992 9272 40044
rect 9680 40035 9732 40044
rect 9680 40001 9689 40035
rect 9689 40001 9723 40035
rect 9723 40001 9732 40035
rect 9680 39992 9732 40001
rect 7104 39967 7156 39976
rect 7104 39933 7113 39967
rect 7113 39933 7147 39967
rect 7147 39933 7156 39967
rect 7104 39924 7156 39933
rect 9128 39967 9180 39976
rect 9128 39933 9137 39967
rect 9137 39933 9171 39967
rect 9171 39933 9180 39967
rect 9128 39924 9180 39933
rect 9496 39924 9548 39976
rect 16856 40060 16908 40112
rect 17224 40060 17276 40112
rect 17408 40060 17460 40112
rect 19064 40060 19116 40112
rect 20168 40060 20220 40112
rect 8484 39788 8536 39840
rect 8668 39831 8720 39840
rect 8668 39797 8677 39831
rect 8677 39797 8711 39831
rect 8711 39797 8720 39831
rect 8668 39788 8720 39797
rect 15476 39992 15528 40044
rect 12072 39924 12124 39976
rect 12808 39967 12860 39976
rect 12808 39933 12817 39967
rect 12817 39933 12851 39967
rect 12851 39933 12860 39967
rect 12808 39924 12860 39933
rect 16120 39924 16172 39976
rect 16212 39967 16264 39976
rect 16212 39933 16221 39967
rect 16221 39933 16255 39967
rect 16255 39933 16264 39967
rect 16212 39924 16264 39933
rect 18512 40035 18564 40044
rect 18512 40001 18521 40035
rect 18521 40001 18555 40035
rect 18555 40001 18564 40035
rect 18512 39992 18564 40001
rect 10968 39856 11020 39908
rect 11060 39856 11112 39908
rect 11888 39788 11940 39840
rect 13360 39831 13412 39840
rect 13360 39797 13369 39831
rect 13369 39797 13403 39831
rect 13403 39797 13412 39831
rect 13360 39788 13412 39797
rect 14004 39788 14056 39840
rect 15108 39788 15160 39840
rect 18420 39899 18472 39908
rect 18420 39865 18429 39899
rect 18429 39865 18463 39899
rect 18463 39865 18472 39899
rect 18788 39924 18840 39976
rect 20444 40060 20496 40112
rect 20996 40060 21048 40112
rect 22192 40128 22244 40180
rect 24032 40128 24084 40180
rect 24124 40171 24176 40180
rect 24124 40137 24133 40171
rect 24133 40137 24167 40171
rect 24167 40137 24176 40171
rect 24124 40128 24176 40137
rect 35992 40171 36044 40180
rect 35992 40137 36001 40171
rect 36001 40137 36035 40171
rect 36035 40137 36044 40171
rect 35992 40128 36044 40137
rect 22192 40035 22244 40044
rect 22192 40001 22201 40035
rect 22201 40001 22235 40035
rect 22235 40001 22244 40035
rect 22192 39992 22244 40001
rect 36084 40060 36136 40112
rect 41144 40060 41196 40112
rect 23572 40035 23624 40044
rect 23572 40001 23609 40035
rect 23609 40001 23624 40035
rect 23572 39992 23624 40001
rect 20720 39924 20772 39976
rect 22008 39924 22060 39976
rect 18420 39856 18472 39865
rect 15752 39831 15804 39840
rect 15752 39797 15761 39831
rect 15761 39797 15795 39831
rect 15795 39797 15804 39831
rect 15752 39788 15804 39797
rect 20260 39788 20312 39840
rect 22376 39788 22428 39840
rect 25872 40035 25924 40044
rect 25872 40001 25881 40035
rect 25881 40001 25915 40035
rect 25915 40001 25924 40035
rect 25872 39992 25924 40001
rect 26976 39992 27028 40044
rect 40592 40035 40644 40044
rect 40592 40001 40601 40035
rect 40601 40001 40635 40035
rect 40635 40001 40644 40035
rect 40592 39992 40644 40001
rect 40776 39992 40828 40044
rect 41880 39992 41932 40044
rect 43260 39992 43312 40044
rect 24584 39967 24636 39976
rect 24584 39933 24593 39967
rect 24593 39933 24627 39967
rect 24627 39933 24636 39967
rect 24584 39924 24636 39933
rect 32312 39924 32364 39976
rect 24216 39856 24268 39908
rect 25228 39831 25280 39840
rect 25228 39797 25237 39831
rect 25237 39797 25271 39831
rect 25271 39797 25280 39831
rect 25228 39788 25280 39797
rect 25320 39831 25372 39840
rect 25320 39797 25329 39831
rect 25329 39797 25363 39831
rect 25363 39797 25372 39831
rect 25320 39788 25372 39797
rect 26700 39788 26752 39840
rect 26792 39788 26844 39840
rect 32772 39788 32824 39840
rect 34520 39967 34572 39976
rect 34520 39933 34529 39967
rect 34529 39933 34563 39967
rect 34563 39933 34572 39967
rect 34520 39924 34572 39933
rect 38476 39967 38528 39976
rect 38476 39933 38485 39967
rect 38485 39933 38519 39967
rect 38519 39933 38528 39967
rect 38476 39924 38528 39933
rect 38752 39967 38804 39976
rect 38752 39933 38761 39967
rect 38761 39933 38795 39967
rect 38795 39933 38804 39967
rect 38752 39924 38804 39933
rect 42800 39924 42852 39976
rect 34704 39788 34756 39840
rect 41144 39831 41196 39840
rect 41144 39797 41153 39831
rect 41153 39797 41187 39831
rect 41187 39797 41196 39831
rect 41144 39788 41196 39797
rect 41236 39831 41288 39840
rect 41236 39797 41245 39831
rect 41245 39797 41279 39831
rect 41279 39797 41288 39831
rect 41236 39788 41288 39797
rect 42892 39788 42944 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 7104 39584 7156 39636
rect 13544 39584 13596 39636
rect 8484 39448 8536 39500
rect 9404 39448 9456 39500
rect 11888 39448 11940 39500
rect 8668 39380 8720 39432
rect 15752 39584 15804 39636
rect 17960 39584 18012 39636
rect 16120 39448 16172 39500
rect 20720 39584 20772 39636
rect 25872 39584 25924 39636
rect 34520 39584 34572 39636
rect 38752 39584 38804 39636
rect 39948 39584 40000 39636
rect 40132 39584 40184 39636
rect 42800 39584 42852 39636
rect 42892 39584 42944 39636
rect 17684 39448 17736 39500
rect 18420 39448 18472 39500
rect 18512 39448 18564 39500
rect 24400 39491 24452 39500
rect 24400 39457 24409 39491
rect 24409 39457 24443 39491
rect 24443 39457 24452 39491
rect 24400 39448 24452 39457
rect 26148 39448 26200 39500
rect 26792 39448 26844 39500
rect 27436 39448 27488 39500
rect 14004 39380 14056 39432
rect 9864 39355 9916 39364
rect 9864 39321 9873 39355
rect 9873 39321 9907 39355
rect 9907 39321 9916 39355
rect 9864 39312 9916 39321
rect 10876 39312 10928 39364
rect 9588 39244 9640 39296
rect 11520 39244 11572 39296
rect 12624 39244 12676 39296
rect 16028 39312 16080 39364
rect 18880 39423 18932 39432
rect 18880 39389 18889 39423
rect 18889 39389 18923 39423
rect 18923 39389 18932 39423
rect 18880 39380 18932 39389
rect 20628 39380 20680 39432
rect 20812 39380 20864 39432
rect 16580 39287 16632 39296
rect 16580 39253 16589 39287
rect 16589 39253 16623 39287
rect 16623 39253 16632 39287
rect 16580 39244 16632 39253
rect 18144 39244 18196 39296
rect 22560 39423 22612 39432
rect 22560 39389 22569 39423
rect 22569 39389 22603 39423
rect 22603 39389 22612 39423
rect 22560 39380 22612 39389
rect 22928 39380 22980 39432
rect 24952 39312 25004 39364
rect 20352 39244 20404 39296
rect 21272 39244 21324 39296
rect 22100 39287 22152 39296
rect 22100 39253 22109 39287
rect 22109 39253 22143 39287
rect 22143 39253 22152 39287
rect 22100 39244 22152 39253
rect 22284 39244 22336 39296
rect 23756 39244 23808 39296
rect 24308 39244 24360 39296
rect 26332 39244 26384 39296
rect 27896 39448 27948 39500
rect 28908 39448 28960 39500
rect 29460 39312 29512 39364
rect 28540 39244 28592 39296
rect 28724 39244 28776 39296
rect 30380 39312 30432 39364
rect 31668 39448 31720 39500
rect 31760 39491 31812 39500
rect 31760 39457 31769 39491
rect 31769 39457 31803 39491
rect 31803 39457 31812 39491
rect 31760 39448 31812 39457
rect 32036 39491 32088 39500
rect 32036 39457 32045 39491
rect 32045 39457 32079 39491
rect 32079 39457 32088 39491
rect 32036 39448 32088 39457
rect 32496 39448 32548 39500
rect 34612 39380 34664 39432
rect 35532 39380 35584 39432
rect 31668 39312 31720 39364
rect 38752 39380 38804 39432
rect 40224 39380 40276 39432
rect 41144 39380 41196 39432
rect 42156 39423 42208 39432
rect 42156 39389 42165 39423
rect 42165 39389 42199 39423
rect 42199 39389 42208 39423
rect 42156 39380 42208 39389
rect 42432 39448 42484 39500
rect 44180 39491 44232 39500
rect 44180 39457 44189 39491
rect 44189 39457 44223 39491
rect 44223 39457 44232 39491
rect 44180 39448 44232 39457
rect 42524 39380 42576 39432
rect 32220 39244 32272 39296
rect 33876 39287 33928 39296
rect 33876 39253 33885 39287
rect 33885 39253 33919 39287
rect 33919 39253 33928 39287
rect 33876 39244 33928 39253
rect 38108 39287 38160 39296
rect 38108 39253 38117 39287
rect 38117 39253 38151 39287
rect 38151 39253 38160 39287
rect 38108 39244 38160 39253
rect 38200 39244 38252 39296
rect 40592 39312 40644 39364
rect 40316 39244 40368 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 9588 39083 9640 39092
rect 9588 39049 9597 39083
rect 9597 39049 9631 39083
rect 9631 39049 9640 39083
rect 9588 39040 9640 39049
rect 9864 39040 9916 39092
rect 9220 38904 9272 38956
rect 7840 38836 7892 38888
rect 8208 38768 8260 38820
rect 9036 38879 9088 38888
rect 9036 38845 9045 38879
rect 9045 38845 9079 38879
rect 9079 38845 9088 38879
rect 9036 38836 9088 38845
rect 9496 38836 9548 38888
rect 10968 39083 11020 39092
rect 10968 39049 10977 39083
rect 10977 39049 11011 39083
rect 11011 39049 11020 39083
rect 10968 39040 11020 39049
rect 12072 39083 12124 39092
rect 12072 39049 12081 39083
rect 12081 39049 12115 39083
rect 12115 39049 12124 39083
rect 12072 39040 12124 39049
rect 12808 39083 12860 39092
rect 12808 39049 12817 39083
rect 12817 39049 12851 39083
rect 12851 39049 12860 39083
rect 12808 39040 12860 39049
rect 12532 38972 12584 39024
rect 13360 39040 13412 39092
rect 15292 39040 15344 39092
rect 18880 39040 18932 39092
rect 20076 39040 20128 39092
rect 20812 39040 20864 39092
rect 24308 39040 24360 39092
rect 24584 39040 24636 39092
rect 31760 39040 31812 39092
rect 11520 38904 11572 38956
rect 14004 38972 14056 39024
rect 10968 38836 11020 38888
rect 11336 38836 11388 38888
rect 11980 38836 12032 38888
rect 12716 38947 12768 38956
rect 12716 38913 12725 38947
rect 12725 38913 12759 38947
rect 12759 38913 12768 38947
rect 12716 38904 12768 38913
rect 13544 38836 13596 38888
rect 14740 38836 14792 38888
rect 7012 38700 7064 38752
rect 12900 38700 12952 38752
rect 13728 38700 13780 38752
rect 17500 38836 17552 38888
rect 20352 38904 20404 38956
rect 20260 38836 20312 38888
rect 18144 38768 18196 38820
rect 18972 38700 19024 38752
rect 23756 38947 23808 38956
rect 23756 38913 23765 38947
rect 23765 38913 23799 38947
rect 23799 38913 23808 38947
rect 23756 38904 23808 38913
rect 21640 38836 21692 38888
rect 22284 38836 22336 38888
rect 23572 38879 23624 38888
rect 23572 38845 23581 38879
rect 23581 38845 23615 38879
rect 23615 38845 23624 38879
rect 23572 38836 23624 38845
rect 20628 38700 20680 38752
rect 22652 38743 22704 38752
rect 22652 38709 22661 38743
rect 22661 38709 22695 38743
rect 22695 38709 22704 38743
rect 22652 38700 22704 38709
rect 24032 38947 24084 38956
rect 24032 38913 24041 38947
rect 24041 38913 24075 38947
rect 24075 38913 24084 38947
rect 24032 38904 24084 38913
rect 24216 38947 24268 38956
rect 24216 38913 24230 38947
rect 24230 38913 24264 38947
rect 24264 38913 24268 38947
rect 24216 38904 24268 38913
rect 24400 38904 24452 38956
rect 25044 38972 25096 39024
rect 26884 38972 26936 39024
rect 26792 38904 26844 38956
rect 28724 38972 28776 39024
rect 32956 39040 33008 39092
rect 32864 38972 32916 39024
rect 27528 38904 27580 38956
rect 25228 38836 25280 38888
rect 26148 38836 26200 38888
rect 26700 38836 26752 38888
rect 27896 38836 27948 38888
rect 24492 38768 24544 38820
rect 28264 38879 28316 38888
rect 28264 38845 28273 38879
rect 28273 38845 28307 38879
rect 28307 38845 28316 38879
rect 28264 38836 28316 38845
rect 29460 38836 29512 38888
rect 25320 38700 25372 38752
rect 26332 38700 26384 38752
rect 26976 38743 27028 38752
rect 26976 38709 26985 38743
rect 26985 38709 27019 38743
rect 27019 38709 27028 38743
rect 26976 38700 27028 38709
rect 29368 38768 29420 38820
rect 29552 38700 29604 38752
rect 32404 38947 32456 38956
rect 32404 38913 32413 38947
rect 32413 38913 32447 38947
rect 32447 38913 32456 38947
rect 32404 38904 32456 38913
rect 32772 38879 32824 38888
rect 32772 38845 32781 38879
rect 32781 38845 32815 38879
rect 32815 38845 32824 38879
rect 32772 38836 32824 38845
rect 32496 38768 32548 38820
rect 33232 39015 33284 39024
rect 33232 38981 33254 39015
rect 33254 38981 33284 39015
rect 33232 38972 33284 38981
rect 38384 39040 38436 39092
rect 44180 39040 44232 39092
rect 35900 38972 35952 39024
rect 38292 38972 38344 39024
rect 33876 38904 33928 38956
rect 34152 38904 34204 38956
rect 40316 38947 40368 38956
rect 40316 38913 40325 38947
rect 40325 38913 40359 38947
rect 40359 38913 40368 38947
rect 40316 38904 40368 38913
rect 33140 38836 33192 38888
rect 36728 38836 36780 38888
rect 38108 38836 38160 38888
rect 39856 38836 39908 38888
rect 40132 38879 40184 38888
rect 40132 38845 40141 38879
rect 40141 38845 40175 38879
rect 40175 38845 40184 38879
rect 40868 38904 40920 38956
rect 40132 38836 40184 38845
rect 33600 38768 33652 38820
rect 36912 38768 36964 38820
rect 33232 38700 33284 38752
rect 35900 38743 35952 38752
rect 35900 38709 35909 38743
rect 35909 38709 35943 38743
rect 35943 38709 35952 38743
rect 35900 38700 35952 38709
rect 37280 38743 37332 38752
rect 37280 38709 37289 38743
rect 37289 38709 37323 38743
rect 37323 38709 37332 38743
rect 37280 38700 37332 38709
rect 40316 38768 40368 38820
rect 38292 38700 38344 38752
rect 40224 38700 40276 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 6736 38360 6788 38412
rect 8392 38496 8444 38548
rect 9588 38496 9640 38548
rect 14740 38496 14792 38548
rect 23572 38539 23624 38548
rect 23572 38505 23581 38539
rect 23581 38505 23615 38539
rect 23615 38505 23624 38539
rect 23572 38496 23624 38505
rect 28264 38496 28316 38548
rect 29368 38496 29420 38548
rect 32404 38496 32456 38548
rect 33232 38539 33284 38548
rect 33232 38505 33241 38539
rect 33241 38505 33275 38539
rect 33275 38505 33284 38539
rect 33232 38496 33284 38505
rect 33600 38496 33652 38548
rect 40868 38496 40920 38548
rect 42524 38496 42576 38548
rect 9036 38360 9088 38412
rect 12716 38428 12768 38480
rect 25044 38428 25096 38480
rect 9680 38292 9732 38344
rect 11428 38335 11480 38344
rect 11428 38301 11437 38335
rect 11437 38301 11471 38335
rect 11471 38301 11480 38335
rect 11428 38292 11480 38301
rect 12532 38292 12584 38344
rect 12900 38292 12952 38344
rect 20720 38360 20772 38412
rect 22100 38403 22152 38412
rect 22100 38369 22109 38403
rect 22109 38369 22143 38403
rect 22143 38369 22152 38403
rect 22100 38360 22152 38369
rect 25412 38403 25464 38412
rect 25412 38369 25421 38403
rect 25421 38369 25455 38403
rect 25455 38369 25464 38403
rect 25412 38360 25464 38369
rect 28908 38360 28960 38412
rect 29552 38360 29604 38412
rect 31576 38360 31628 38412
rect 7012 38224 7064 38276
rect 9220 38224 9272 38276
rect 10876 38267 10928 38276
rect 10876 38233 10885 38267
rect 10885 38233 10919 38267
rect 10919 38233 10928 38267
rect 10876 38224 10928 38233
rect 9956 38199 10008 38208
rect 9956 38165 9965 38199
rect 9965 38165 9999 38199
rect 9999 38165 10008 38199
rect 9956 38156 10008 38165
rect 13360 38335 13412 38344
rect 13360 38301 13369 38335
rect 13369 38301 13403 38335
rect 13403 38301 13412 38335
rect 13360 38292 13412 38301
rect 13728 38292 13780 38344
rect 16948 38292 17000 38344
rect 18880 38335 18932 38344
rect 18880 38301 18889 38335
rect 18889 38301 18923 38335
rect 18923 38301 18932 38335
rect 18880 38292 18932 38301
rect 28540 38335 28592 38344
rect 28540 38301 28549 38335
rect 28549 38301 28583 38335
rect 28583 38301 28592 38335
rect 28540 38292 28592 38301
rect 29460 38292 29512 38344
rect 33140 38428 33192 38480
rect 15292 38224 15344 38276
rect 16488 38224 16540 38276
rect 17960 38267 18012 38276
rect 17960 38233 17969 38267
rect 17969 38233 18003 38267
rect 18003 38233 18012 38267
rect 17960 38224 18012 38233
rect 20260 38267 20312 38276
rect 20260 38233 20269 38267
rect 20269 38233 20303 38267
rect 20303 38233 20312 38267
rect 20260 38224 20312 38233
rect 22560 38224 22612 38276
rect 27160 38267 27212 38276
rect 27160 38233 27169 38267
rect 27169 38233 27203 38267
rect 27203 38233 27212 38267
rect 27160 38224 27212 38233
rect 28632 38267 28684 38276
rect 28632 38233 28641 38267
rect 28641 38233 28675 38267
rect 28675 38233 28684 38267
rect 28632 38224 28684 38233
rect 17316 38156 17368 38208
rect 17776 38156 17828 38208
rect 20628 38156 20680 38208
rect 21640 38156 21692 38208
rect 29920 38267 29972 38276
rect 29920 38233 29929 38267
rect 29929 38233 29963 38267
rect 29963 38233 29972 38267
rect 29920 38224 29972 38233
rect 30380 38224 30432 38276
rect 33232 38335 33284 38344
rect 33232 38301 33241 38335
rect 33241 38301 33275 38335
rect 33275 38301 33284 38335
rect 33232 38292 33284 38301
rect 33508 38360 33560 38412
rect 33416 38292 33468 38344
rect 38292 38360 38344 38412
rect 34796 38292 34848 38344
rect 36912 38292 36964 38344
rect 37280 38292 37332 38344
rect 37372 38292 37424 38344
rect 37924 38335 37976 38344
rect 37924 38301 37933 38335
rect 37933 38301 37967 38335
rect 37967 38301 37976 38335
rect 37924 38292 37976 38301
rect 39856 38335 39908 38344
rect 39856 38301 39865 38335
rect 39865 38301 39899 38335
rect 39899 38301 39908 38335
rect 39856 38292 39908 38301
rect 42708 38403 42760 38412
rect 42708 38369 42717 38403
rect 42717 38369 42751 38403
rect 42751 38369 42760 38403
rect 42708 38360 42760 38369
rect 42800 38360 42852 38412
rect 42616 38335 42668 38344
rect 42616 38301 42625 38335
rect 42625 38301 42659 38335
rect 42659 38301 42668 38335
rect 42616 38292 42668 38301
rect 43260 38335 43312 38344
rect 43260 38301 43269 38335
rect 43269 38301 43303 38335
rect 43303 38301 43312 38335
rect 43260 38292 43312 38301
rect 33876 38224 33928 38276
rect 35256 38267 35308 38276
rect 35256 38233 35265 38267
rect 35265 38233 35299 38267
rect 35299 38233 35308 38267
rect 35256 38224 35308 38233
rect 40040 38224 40092 38276
rect 40132 38267 40184 38276
rect 40132 38233 40141 38267
rect 40141 38233 40175 38267
rect 40175 38233 40184 38267
rect 40132 38224 40184 38233
rect 30104 38156 30156 38208
rect 31484 38199 31536 38208
rect 31484 38165 31493 38199
rect 31493 38165 31527 38199
rect 31527 38165 31536 38199
rect 31484 38156 31536 38165
rect 33232 38156 33284 38208
rect 36728 38199 36780 38208
rect 36728 38165 36737 38199
rect 36737 38165 36771 38199
rect 36771 38165 36780 38199
rect 36728 38156 36780 38165
rect 38660 38199 38712 38208
rect 38660 38165 38669 38199
rect 38669 38165 38703 38199
rect 38703 38165 38712 38199
rect 38660 38156 38712 38165
rect 42156 38156 42208 38208
rect 42984 38199 43036 38208
rect 42984 38165 42993 38199
rect 42993 38165 43027 38199
rect 43027 38165 43036 38199
rect 42984 38156 43036 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 6736 37884 6788 37936
rect 8392 37884 8444 37936
rect 9956 37952 10008 38004
rect 11428 37952 11480 38004
rect 13728 37952 13780 38004
rect 15292 37884 15344 37936
rect 9404 37859 9456 37868
rect 9404 37825 9413 37859
rect 9413 37825 9447 37859
rect 9447 37825 9456 37859
rect 9404 37816 9456 37825
rect 10968 37816 11020 37868
rect 12900 37816 12952 37868
rect 13360 37859 13412 37868
rect 13360 37825 13369 37859
rect 13369 37825 13403 37859
rect 13403 37825 13412 37859
rect 13360 37816 13412 37825
rect 6920 37748 6972 37800
rect 8944 37791 8996 37800
rect 8944 37757 8953 37791
rect 8953 37757 8987 37791
rect 8987 37757 8996 37791
rect 8944 37748 8996 37757
rect 8392 37655 8444 37664
rect 8392 37621 8401 37655
rect 8401 37621 8435 37655
rect 8435 37621 8444 37655
rect 8392 37612 8444 37621
rect 12992 37655 13044 37664
rect 12992 37621 13001 37655
rect 13001 37621 13035 37655
rect 13035 37621 13044 37655
rect 12992 37612 13044 37621
rect 14004 37748 14056 37800
rect 15292 37748 15344 37800
rect 17776 37952 17828 38004
rect 17960 37952 18012 38004
rect 19248 37952 19300 38004
rect 20260 37952 20312 38004
rect 17040 37859 17092 37868
rect 17040 37825 17049 37859
rect 17049 37825 17083 37859
rect 17083 37825 17092 37859
rect 17040 37816 17092 37825
rect 17316 37859 17368 37868
rect 17316 37825 17325 37859
rect 17325 37825 17359 37859
rect 17359 37825 17368 37859
rect 17316 37816 17368 37825
rect 17408 37859 17460 37868
rect 17408 37825 17417 37859
rect 17417 37825 17451 37859
rect 17451 37825 17460 37859
rect 17408 37816 17460 37825
rect 18512 37816 18564 37868
rect 16672 37680 16724 37732
rect 16028 37655 16080 37664
rect 16028 37621 16037 37655
rect 16037 37621 16071 37655
rect 16071 37621 16080 37655
rect 16028 37612 16080 37621
rect 18880 37612 18932 37664
rect 20720 37816 20772 37868
rect 22652 37952 22704 38004
rect 24860 37952 24912 38004
rect 27528 37952 27580 38004
rect 22284 37927 22336 37936
rect 22284 37893 22293 37927
rect 22293 37893 22327 37927
rect 22327 37893 22336 37927
rect 22284 37884 22336 37893
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 27712 37884 27764 37936
rect 20996 37791 21048 37800
rect 20996 37757 21005 37791
rect 21005 37757 21039 37791
rect 21039 37757 21048 37791
rect 20996 37748 21048 37757
rect 22376 37791 22428 37800
rect 22376 37757 22385 37791
rect 22385 37757 22419 37791
rect 22419 37757 22428 37791
rect 22376 37748 22428 37757
rect 24768 37680 24820 37732
rect 27436 37859 27488 37868
rect 28724 37884 28776 37936
rect 29920 37952 29972 38004
rect 33140 37995 33192 38004
rect 33140 37961 33149 37995
rect 33149 37961 33183 37995
rect 33183 37961 33192 37995
rect 33140 37952 33192 37961
rect 35532 37952 35584 38004
rect 27436 37825 27471 37859
rect 27471 37825 27488 37859
rect 27436 37816 27488 37825
rect 27804 37748 27856 37800
rect 32956 37884 33008 37936
rect 37924 37952 37976 38004
rect 38660 37952 38712 38004
rect 38752 37952 38804 38004
rect 40132 37952 40184 38004
rect 42616 37995 42668 38004
rect 42616 37961 42625 37995
rect 42625 37961 42659 37995
rect 42659 37961 42668 37995
rect 42616 37952 42668 37961
rect 42984 37952 43036 38004
rect 30104 37816 30156 37868
rect 22560 37612 22612 37664
rect 26976 37655 27028 37664
rect 26976 37621 26985 37655
rect 26985 37621 27019 37655
rect 27019 37621 27028 37655
rect 26976 37612 27028 37621
rect 27896 37680 27948 37732
rect 28632 37680 28684 37732
rect 29000 37655 29052 37664
rect 29000 37621 29009 37655
rect 29009 37621 29043 37655
rect 29043 37621 29052 37655
rect 29000 37612 29052 37621
rect 29460 37612 29512 37664
rect 31484 37816 31536 37868
rect 33416 37816 33468 37868
rect 33508 37859 33560 37868
rect 33508 37825 33517 37859
rect 33517 37825 33551 37859
rect 33551 37825 33560 37859
rect 33508 37816 33560 37825
rect 36728 37884 36780 37936
rect 32864 37748 32916 37800
rect 31208 37680 31260 37732
rect 36820 37816 36872 37868
rect 35256 37748 35308 37800
rect 35900 37748 35952 37800
rect 32956 37612 33008 37664
rect 35808 37655 35860 37664
rect 35808 37621 35817 37655
rect 35817 37621 35851 37655
rect 35851 37621 35860 37655
rect 35808 37612 35860 37621
rect 35992 37612 36044 37664
rect 37280 37748 37332 37800
rect 38016 37748 38068 37800
rect 40224 37859 40276 37868
rect 40224 37825 40233 37859
rect 40233 37825 40267 37859
rect 40267 37825 40276 37859
rect 40224 37816 40276 37825
rect 40316 37816 40368 37868
rect 39488 37748 39540 37800
rect 39948 37791 40000 37800
rect 39948 37757 39957 37791
rect 39957 37757 39991 37791
rect 39991 37757 40000 37791
rect 39948 37748 40000 37757
rect 43168 37791 43220 37800
rect 43168 37757 43177 37791
rect 43177 37757 43211 37791
rect 43211 37757 43220 37791
rect 43168 37748 43220 37757
rect 37832 37655 37884 37664
rect 37832 37621 37841 37655
rect 37841 37621 37875 37655
rect 37875 37621 37884 37655
rect 37832 37612 37884 37621
rect 38200 37612 38252 37664
rect 38660 37655 38712 37664
rect 38660 37621 38669 37655
rect 38669 37621 38703 37655
rect 38703 37621 38712 37655
rect 38660 37612 38712 37621
rect 38844 37612 38896 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 6920 37408 6972 37460
rect 8944 37408 8996 37460
rect 17040 37408 17092 37460
rect 20720 37451 20772 37460
rect 20720 37417 20729 37451
rect 20729 37417 20763 37451
rect 20763 37417 20772 37451
rect 20720 37408 20772 37417
rect 8208 37315 8260 37324
rect 8208 37281 8217 37315
rect 8217 37281 8251 37315
rect 8251 37281 8260 37315
rect 8208 37272 8260 37281
rect 940 37204 992 37256
rect 1768 37204 1820 37256
rect 5540 37204 5592 37256
rect 2136 37068 2188 37120
rect 8392 37204 8444 37256
rect 9220 37340 9272 37392
rect 11060 37340 11112 37392
rect 10876 37272 10928 37324
rect 11428 37272 11480 37324
rect 12992 37272 13044 37324
rect 12256 37204 12308 37256
rect 13360 37204 13412 37256
rect 16028 37315 16080 37324
rect 16028 37281 16037 37315
rect 16037 37281 16071 37315
rect 16071 37281 16080 37315
rect 16028 37272 16080 37281
rect 16488 37340 16540 37392
rect 16856 37204 16908 37256
rect 16948 37204 17000 37256
rect 18512 37272 18564 37324
rect 22468 37408 22520 37460
rect 27804 37451 27856 37460
rect 27804 37417 27813 37451
rect 27813 37417 27847 37451
rect 27847 37417 27856 37451
rect 27804 37408 27856 37417
rect 36820 37451 36872 37460
rect 36820 37417 36829 37451
rect 36829 37417 36863 37451
rect 36863 37417 36872 37451
rect 36820 37408 36872 37417
rect 39488 37408 39540 37460
rect 28632 37340 28684 37392
rect 30012 37340 30064 37392
rect 19156 37204 19208 37256
rect 12900 37136 12952 37188
rect 16028 37136 16080 37188
rect 17316 37179 17368 37188
rect 17316 37145 17325 37179
rect 17325 37145 17359 37179
rect 17359 37145 17368 37179
rect 17316 37136 17368 37145
rect 19064 37136 19116 37188
rect 25412 37272 25464 37324
rect 26976 37272 27028 37324
rect 27528 37272 27580 37324
rect 32772 37272 32824 37324
rect 34796 37272 34848 37324
rect 35992 37272 36044 37324
rect 21732 37204 21784 37256
rect 23848 37247 23900 37256
rect 23848 37213 23857 37247
rect 23857 37213 23891 37247
rect 23891 37213 23900 37247
rect 23848 37204 23900 37213
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 25320 37204 25372 37256
rect 25688 37247 25740 37256
rect 25688 37213 25697 37247
rect 25697 37213 25731 37247
rect 25731 37213 25740 37247
rect 25688 37204 25740 37213
rect 7748 37068 7800 37120
rect 10692 37111 10744 37120
rect 10692 37077 10701 37111
rect 10701 37077 10735 37111
rect 10735 37077 10744 37111
rect 10692 37068 10744 37077
rect 11060 37111 11112 37120
rect 11060 37077 11069 37111
rect 11069 37077 11103 37111
rect 11103 37077 11112 37111
rect 11060 37068 11112 37077
rect 13452 37068 13504 37120
rect 13636 37068 13688 37120
rect 15200 37111 15252 37120
rect 15200 37077 15209 37111
rect 15209 37077 15243 37111
rect 15243 37077 15252 37111
rect 15200 37068 15252 37077
rect 18788 37111 18840 37120
rect 18788 37077 18797 37111
rect 18797 37077 18831 37111
rect 18831 37077 18840 37111
rect 18788 37068 18840 37077
rect 18972 37068 19024 37120
rect 23756 37068 23808 37120
rect 23940 37068 23992 37120
rect 25044 37111 25096 37120
rect 25044 37077 25053 37111
rect 25053 37077 25087 37111
rect 25087 37077 25096 37111
rect 25044 37068 25096 37077
rect 33508 37204 33560 37256
rect 36912 37204 36964 37256
rect 37832 37315 37884 37324
rect 37832 37281 37841 37315
rect 37841 37281 37875 37315
rect 37875 37281 37884 37315
rect 37832 37272 37884 37281
rect 38016 37247 38068 37256
rect 38016 37213 38025 37247
rect 38025 37213 38059 37247
rect 38059 37213 38068 37247
rect 38016 37204 38068 37213
rect 38660 37204 38712 37256
rect 38844 37204 38896 37256
rect 40040 37204 40092 37256
rect 41236 37272 41288 37324
rect 26792 37136 26844 37188
rect 33876 37136 33928 37188
rect 34060 37136 34112 37188
rect 35348 37179 35400 37188
rect 35348 37145 35357 37179
rect 35357 37145 35391 37179
rect 35391 37145 35400 37179
rect 35348 37136 35400 37145
rect 27620 37068 27672 37120
rect 33324 37068 33376 37120
rect 42248 37451 42300 37460
rect 42248 37417 42257 37451
rect 42257 37417 42291 37451
rect 42291 37417 42300 37451
rect 42248 37408 42300 37417
rect 42984 37204 43036 37256
rect 44272 37247 44324 37256
rect 44272 37213 44281 37247
rect 44281 37213 44315 37247
rect 44315 37213 44324 37247
rect 44272 37204 44324 37213
rect 42616 37136 42668 37188
rect 41144 37068 41196 37120
rect 41236 37111 41288 37120
rect 41236 37077 41245 37111
rect 41245 37077 41279 37111
rect 41279 37077 41288 37111
rect 41236 37068 41288 37077
rect 41420 37111 41472 37120
rect 41420 37077 41429 37111
rect 41429 37077 41463 37111
rect 41463 37077 41472 37111
rect 41420 37068 41472 37077
rect 41604 37111 41656 37120
rect 41604 37077 41613 37111
rect 41613 37077 41647 37111
rect 41647 37077 41656 37111
rect 41604 37068 41656 37077
rect 41788 37068 41840 37120
rect 43168 37068 43220 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 12256 36907 12308 36916
rect 12256 36873 12265 36907
rect 12265 36873 12299 36907
rect 12299 36873 12308 36907
rect 12256 36864 12308 36873
rect 13452 36864 13504 36916
rect 6736 36796 6788 36848
rect 15200 36864 15252 36916
rect 15292 36907 15344 36916
rect 15292 36873 15301 36907
rect 15301 36873 15335 36907
rect 15335 36873 15344 36907
rect 15292 36864 15344 36873
rect 16672 36864 16724 36916
rect 17316 36907 17368 36916
rect 17316 36873 17325 36907
rect 17325 36873 17359 36907
rect 17359 36873 17368 36907
rect 17316 36864 17368 36873
rect 18788 36864 18840 36916
rect 18880 36864 18932 36916
rect 1768 36703 1820 36712
rect 1768 36669 1777 36703
rect 1777 36669 1811 36703
rect 1811 36669 1820 36703
rect 1768 36660 1820 36669
rect 4620 36703 4672 36712
rect 4620 36669 4629 36703
rect 4629 36669 4663 36703
rect 4663 36669 4672 36703
rect 4620 36660 4672 36669
rect 2136 36635 2188 36644
rect 2136 36601 2145 36635
rect 2145 36601 2179 36635
rect 2179 36601 2188 36635
rect 2136 36592 2188 36601
rect 8208 36728 8260 36780
rect 10968 36728 11020 36780
rect 12624 36728 12676 36780
rect 14004 36771 14056 36780
rect 14004 36737 14013 36771
rect 14013 36737 14047 36771
rect 14047 36737 14056 36771
rect 14004 36728 14056 36737
rect 16028 36839 16080 36848
rect 16028 36805 16037 36839
rect 16037 36805 16071 36839
rect 16071 36805 16080 36839
rect 16028 36796 16080 36805
rect 16672 36728 16724 36780
rect 17132 36796 17184 36848
rect 17224 36796 17276 36848
rect 20996 36864 21048 36916
rect 23848 36907 23900 36916
rect 23848 36873 23857 36907
rect 23857 36873 23891 36907
rect 23891 36873 23900 36907
rect 23848 36864 23900 36873
rect 25044 36864 25096 36916
rect 25412 36864 25464 36916
rect 27712 36864 27764 36916
rect 31208 36864 31260 36916
rect 31668 36864 31720 36916
rect 6368 36660 6420 36712
rect 8300 36660 8352 36712
rect 9404 36660 9456 36712
rect 9864 36703 9916 36712
rect 9864 36669 9873 36703
rect 9873 36669 9907 36703
rect 9907 36669 9916 36703
rect 9864 36660 9916 36669
rect 12164 36660 12216 36712
rect 17040 36771 17092 36780
rect 17040 36737 17049 36771
rect 17049 36737 17083 36771
rect 17083 36737 17092 36771
rect 17040 36728 17092 36737
rect 18788 36771 18840 36780
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 18972 36771 19024 36780
rect 18972 36737 18979 36771
rect 18979 36737 19024 36771
rect 18972 36728 19024 36737
rect 19064 36771 19116 36780
rect 19064 36737 19073 36771
rect 19073 36737 19107 36771
rect 19107 36737 19116 36771
rect 19064 36728 19116 36737
rect 19248 36771 19300 36780
rect 19248 36737 19262 36771
rect 19262 36737 19296 36771
rect 19296 36737 19300 36771
rect 19248 36728 19300 36737
rect 19340 36660 19392 36712
rect 2228 36567 2280 36576
rect 2228 36533 2237 36567
rect 2237 36533 2271 36567
rect 2271 36533 2280 36567
rect 2228 36524 2280 36533
rect 5816 36524 5868 36576
rect 8668 36524 8720 36576
rect 11060 36524 11112 36576
rect 12072 36524 12124 36576
rect 20536 36660 20588 36712
rect 23940 36796 23992 36848
rect 22560 36771 22612 36780
rect 22560 36737 22569 36771
rect 22569 36737 22603 36771
rect 22603 36737 22612 36771
rect 22560 36728 22612 36737
rect 22744 36703 22796 36712
rect 22744 36669 22753 36703
rect 22753 36669 22787 36703
rect 22787 36669 22796 36703
rect 22744 36660 22796 36669
rect 23664 36703 23716 36712
rect 23664 36669 23673 36703
rect 23673 36669 23707 36703
rect 23707 36669 23716 36703
rect 23664 36660 23716 36669
rect 25964 36771 26016 36780
rect 25964 36737 25973 36771
rect 25973 36737 26007 36771
rect 26007 36737 26016 36771
rect 25964 36728 26016 36737
rect 27068 36728 27120 36780
rect 28172 36771 28224 36780
rect 28172 36737 28181 36771
rect 28181 36737 28215 36771
rect 28215 36737 28224 36771
rect 28172 36728 28224 36737
rect 29000 36796 29052 36848
rect 30196 36728 30248 36780
rect 25228 36660 25280 36712
rect 33140 36864 33192 36916
rect 16396 36524 16448 36576
rect 21180 36567 21232 36576
rect 21180 36533 21189 36567
rect 21189 36533 21223 36567
rect 21223 36533 21232 36567
rect 21180 36524 21232 36533
rect 22192 36567 22244 36576
rect 22192 36533 22201 36567
rect 22201 36533 22235 36567
rect 22235 36533 22244 36567
rect 22192 36524 22244 36533
rect 23112 36567 23164 36576
rect 23112 36533 23121 36567
rect 23121 36533 23155 36567
rect 23155 36533 23164 36567
rect 23112 36524 23164 36533
rect 24860 36524 24912 36576
rect 26976 36567 27028 36576
rect 26976 36533 26985 36567
rect 26985 36533 27019 36567
rect 27019 36533 27028 36567
rect 26976 36524 27028 36533
rect 27436 36524 27488 36576
rect 27528 36567 27580 36576
rect 27528 36533 27537 36567
rect 27537 36533 27571 36567
rect 27571 36533 27580 36567
rect 27528 36524 27580 36533
rect 27620 36524 27672 36576
rect 31116 36524 31168 36576
rect 32680 36703 32732 36712
rect 32680 36669 32689 36703
rect 32689 36669 32723 36703
rect 32723 36669 32732 36703
rect 32680 36660 32732 36669
rect 33232 36703 33284 36712
rect 33232 36669 33241 36703
rect 33241 36669 33275 36703
rect 33275 36669 33284 36703
rect 33232 36660 33284 36669
rect 33416 36728 33468 36780
rect 33876 36907 33928 36916
rect 33876 36873 33885 36907
rect 33885 36873 33919 36907
rect 33919 36873 33928 36907
rect 33876 36864 33928 36873
rect 34060 36907 34112 36916
rect 34060 36873 34069 36907
rect 34069 36873 34103 36907
rect 34103 36873 34112 36907
rect 34060 36864 34112 36873
rect 35348 36864 35400 36916
rect 35808 36796 35860 36848
rect 41604 36864 41656 36916
rect 41788 36864 41840 36916
rect 42248 36864 42300 36916
rect 33876 36728 33928 36780
rect 33968 36771 34020 36780
rect 33968 36737 33977 36771
rect 33977 36737 34011 36771
rect 34011 36737 34020 36771
rect 33968 36728 34020 36737
rect 34244 36771 34296 36780
rect 34244 36737 34253 36771
rect 34253 36737 34287 36771
rect 34287 36737 34296 36771
rect 34244 36728 34296 36737
rect 32956 36592 33008 36644
rect 33324 36592 33376 36644
rect 33232 36524 33284 36576
rect 38016 36771 38068 36780
rect 38016 36737 38025 36771
rect 38025 36737 38059 36771
rect 38059 36737 38068 36771
rect 38016 36728 38068 36737
rect 38660 36728 38712 36780
rect 38844 36660 38896 36712
rect 39948 36592 40000 36644
rect 40132 36592 40184 36644
rect 35992 36524 36044 36576
rect 37740 36567 37792 36576
rect 37740 36533 37749 36567
rect 37749 36533 37783 36567
rect 37783 36533 37792 36567
rect 37740 36524 37792 36533
rect 42248 36771 42300 36780
rect 42248 36737 42257 36771
rect 42257 36737 42291 36771
rect 42291 36737 42300 36771
rect 42248 36728 42300 36737
rect 44272 36864 44324 36916
rect 42984 36796 43036 36848
rect 43076 36524 43128 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4620 36320 4672 36372
rect 8208 36320 8260 36372
rect 13268 36320 13320 36372
rect 21180 36320 21232 36372
rect 21732 36363 21784 36372
rect 21732 36329 21741 36363
rect 21741 36329 21775 36363
rect 21775 36329 21784 36363
rect 21732 36320 21784 36329
rect 22192 36320 22244 36372
rect 23664 36320 23716 36372
rect 24400 36363 24452 36372
rect 24400 36329 24409 36363
rect 24409 36329 24443 36363
rect 24443 36329 24452 36363
rect 24400 36320 24452 36329
rect 28172 36320 28224 36372
rect 31668 36320 31720 36372
rect 8668 36295 8720 36304
rect 8668 36261 8677 36295
rect 8677 36261 8711 36295
rect 8711 36261 8720 36295
rect 8668 36252 8720 36261
rect 8852 36252 8904 36304
rect 9864 36252 9916 36304
rect 10692 36252 10744 36304
rect 6736 36184 6788 36236
rect 9404 36184 9456 36236
rect 6092 36159 6144 36168
rect 6092 36125 6101 36159
rect 6101 36125 6135 36159
rect 6135 36125 6144 36159
rect 6092 36116 6144 36125
rect 4068 36091 4120 36100
rect 4068 36057 4077 36091
rect 4077 36057 4111 36091
rect 4111 36057 4120 36091
rect 4068 36048 4120 36057
rect 5816 36048 5868 36100
rect 5724 35980 5776 36032
rect 7196 36091 7248 36100
rect 7196 36057 7205 36091
rect 7205 36057 7239 36091
rect 7239 36057 7248 36091
rect 7196 36048 7248 36057
rect 7380 35980 7432 36032
rect 8484 36116 8536 36168
rect 14004 36184 14056 36236
rect 16948 36184 17000 36236
rect 22100 36252 22152 36304
rect 17500 36184 17552 36236
rect 20720 36184 20772 36236
rect 24860 36252 24912 36304
rect 12164 36048 12216 36100
rect 16488 36116 16540 36168
rect 23112 36184 23164 36236
rect 23572 36184 23624 36236
rect 25412 36184 25464 36236
rect 26976 36184 27028 36236
rect 23756 36159 23808 36168
rect 23756 36125 23765 36159
rect 23765 36125 23799 36159
rect 23799 36125 23808 36159
rect 23756 36116 23808 36125
rect 23940 36159 23992 36168
rect 23940 36125 23949 36159
rect 23949 36125 23983 36159
rect 23983 36125 23992 36159
rect 23940 36116 23992 36125
rect 24032 36159 24084 36168
rect 24032 36125 24041 36159
rect 24041 36125 24075 36159
rect 24075 36125 24084 36159
rect 24032 36116 24084 36125
rect 24860 36116 24912 36168
rect 24952 36159 25004 36168
rect 24952 36125 24960 36159
rect 24960 36125 24994 36159
rect 24994 36125 25004 36159
rect 24952 36116 25004 36125
rect 12440 35980 12492 36032
rect 13452 35980 13504 36032
rect 15200 36091 15252 36100
rect 15200 36057 15209 36091
rect 15209 36057 15243 36091
rect 15243 36057 15252 36091
rect 15200 36048 15252 36057
rect 20628 36048 20680 36100
rect 22468 36048 22520 36100
rect 14096 36023 14148 36032
rect 14096 35989 14105 36023
rect 14105 35989 14139 36023
rect 14139 35989 14148 36023
rect 14096 35980 14148 35989
rect 16764 36023 16816 36032
rect 16764 35989 16773 36023
rect 16773 35989 16807 36023
rect 16807 35989 16816 36023
rect 16764 35980 16816 35989
rect 20536 35980 20588 36032
rect 23848 36048 23900 36100
rect 24768 36091 24820 36100
rect 24768 36057 24777 36091
rect 24777 36057 24811 36091
rect 24811 36057 24820 36091
rect 24768 36048 24820 36057
rect 25228 36116 25280 36168
rect 25964 36116 26016 36168
rect 29000 36116 29052 36168
rect 31116 36184 31168 36236
rect 31392 36227 31444 36236
rect 31392 36193 31401 36227
rect 31401 36193 31435 36227
rect 31435 36193 31444 36227
rect 31392 36184 31444 36193
rect 26792 36048 26844 36100
rect 29368 36048 29420 36100
rect 28080 36023 28132 36032
rect 28080 35989 28089 36023
rect 28089 35989 28123 36023
rect 28123 35989 28132 36023
rect 28080 35980 28132 35989
rect 28540 35980 28592 36032
rect 29644 36023 29696 36032
rect 29644 35989 29653 36023
rect 29653 35989 29687 36023
rect 29687 35989 29696 36023
rect 29644 35980 29696 35989
rect 30564 36116 30616 36168
rect 31576 36116 31628 36168
rect 32404 36363 32456 36372
rect 32404 36329 32413 36363
rect 32413 36329 32447 36363
rect 32447 36329 32456 36363
rect 32404 36320 32456 36329
rect 32680 36320 32732 36372
rect 33140 36320 33192 36372
rect 33968 36320 34020 36372
rect 34244 36320 34296 36372
rect 38844 36363 38896 36372
rect 38844 36329 38853 36363
rect 38853 36329 38887 36363
rect 38887 36329 38896 36363
rect 38844 36320 38896 36329
rect 41420 36320 41472 36372
rect 42616 36320 42668 36372
rect 43168 36320 43220 36372
rect 33324 36252 33376 36304
rect 33876 36184 33928 36236
rect 37740 36184 37792 36236
rect 40132 36227 40184 36236
rect 40132 36193 40141 36227
rect 40141 36193 40175 36227
rect 40175 36193 40184 36227
rect 40132 36184 40184 36193
rect 30012 36091 30064 36100
rect 30012 36057 30021 36091
rect 30021 36057 30055 36091
rect 30055 36057 30064 36091
rect 30012 36048 30064 36057
rect 30104 36091 30156 36100
rect 30104 36057 30139 36091
rect 30139 36057 30156 36091
rect 30104 36048 30156 36057
rect 30656 35980 30708 36032
rect 31116 36023 31168 36032
rect 31116 35989 31125 36023
rect 31125 35989 31159 36023
rect 31159 35989 31168 36023
rect 33324 36159 33376 36168
rect 33324 36125 33333 36159
rect 33333 36125 33367 36159
rect 33367 36125 33376 36159
rect 33324 36116 33376 36125
rect 33508 36116 33560 36168
rect 36912 36116 36964 36168
rect 37096 36159 37148 36168
rect 37096 36125 37105 36159
rect 37105 36125 37139 36159
rect 37139 36125 37148 36159
rect 37096 36116 37148 36125
rect 39580 36116 39632 36168
rect 39948 36159 40000 36168
rect 39948 36125 39957 36159
rect 39957 36125 39991 36159
rect 39991 36125 40000 36159
rect 39948 36116 40000 36125
rect 42708 36159 42760 36168
rect 42708 36125 42717 36159
rect 42717 36125 42751 36159
rect 42751 36125 42760 36159
rect 42708 36116 42760 36125
rect 43076 36116 43128 36168
rect 33600 36091 33652 36100
rect 33600 36057 33609 36091
rect 33609 36057 33643 36091
rect 33643 36057 33652 36091
rect 33600 36048 33652 36057
rect 31116 35980 31168 35989
rect 32128 36023 32180 36032
rect 32128 35989 32137 36023
rect 32137 35989 32171 36023
rect 32171 35989 32180 36023
rect 32128 35980 32180 35989
rect 32496 35980 32548 36032
rect 33140 35980 33192 36032
rect 34152 36048 34204 36100
rect 38844 35980 38896 36032
rect 39764 35980 39816 36032
rect 42248 35980 42300 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4068 35776 4120 35828
rect 6092 35776 6144 35828
rect 7196 35776 7248 35828
rect 12440 35776 12492 35828
rect 13360 35776 13412 35828
rect 14096 35776 14148 35828
rect 15200 35776 15252 35828
rect 16764 35776 16816 35828
rect 16856 35776 16908 35828
rect 20536 35776 20588 35828
rect 2228 35640 2280 35692
rect 5540 35708 5592 35760
rect 15936 35708 15988 35760
rect 6920 35640 6972 35692
rect 7564 35640 7616 35692
rect 7656 35683 7708 35692
rect 7656 35649 7665 35683
rect 7665 35649 7699 35683
rect 7699 35649 7708 35683
rect 7656 35640 7708 35649
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 5632 35479 5684 35488
rect 5632 35445 5641 35479
rect 5641 35445 5675 35479
rect 5675 35445 5684 35479
rect 5632 35436 5684 35445
rect 12808 35436 12860 35488
rect 16764 35640 16816 35692
rect 20260 35708 20312 35760
rect 18604 35615 18656 35624
rect 18604 35581 18613 35615
rect 18613 35581 18647 35615
rect 18647 35581 18656 35615
rect 18604 35572 18656 35581
rect 19248 35572 19300 35624
rect 22560 35776 22612 35828
rect 24952 35776 25004 35828
rect 27068 35776 27120 35828
rect 28080 35776 28132 35828
rect 18052 35436 18104 35488
rect 18972 35436 19024 35488
rect 19248 35436 19300 35488
rect 20444 35436 20496 35488
rect 20628 35436 20680 35488
rect 25964 35708 26016 35760
rect 26424 35708 26476 35760
rect 23572 35683 23624 35692
rect 23572 35649 23581 35683
rect 23581 35649 23615 35683
rect 23615 35649 23624 35683
rect 23572 35640 23624 35649
rect 22100 35572 22152 35624
rect 26056 35615 26108 35624
rect 26056 35581 26065 35615
rect 26065 35581 26099 35615
rect 26099 35581 26108 35615
rect 26056 35572 26108 35581
rect 27896 35708 27948 35760
rect 29644 35776 29696 35828
rect 30564 35776 30616 35828
rect 30656 35819 30708 35828
rect 30656 35785 30665 35819
rect 30665 35785 30699 35819
rect 30699 35785 30708 35819
rect 30656 35776 30708 35785
rect 29368 35708 29420 35760
rect 31760 35776 31812 35828
rect 32128 35776 32180 35828
rect 28172 35640 28224 35692
rect 28540 35640 28592 35692
rect 31116 35708 31168 35760
rect 31208 35708 31260 35760
rect 31668 35708 31720 35760
rect 27896 35615 27948 35624
rect 27896 35581 27905 35615
rect 27905 35581 27939 35615
rect 27939 35581 27948 35615
rect 27896 35572 27948 35581
rect 28632 35615 28684 35624
rect 28632 35581 28641 35615
rect 28641 35581 28675 35615
rect 28675 35581 28684 35615
rect 28632 35572 28684 35581
rect 31392 35640 31444 35692
rect 32588 35751 32640 35760
rect 32588 35717 32597 35751
rect 32597 35717 32631 35751
rect 32631 35717 32640 35751
rect 32588 35708 32640 35717
rect 32312 35683 32364 35692
rect 32312 35649 32336 35683
rect 32336 35649 32364 35683
rect 32312 35640 32364 35649
rect 33232 35751 33284 35760
rect 33232 35717 33241 35751
rect 33241 35717 33275 35751
rect 33275 35717 33284 35751
rect 33232 35708 33284 35717
rect 33324 35708 33376 35760
rect 36912 35708 36964 35760
rect 39764 35776 39816 35828
rect 26792 35436 26844 35488
rect 27528 35436 27580 35488
rect 27620 35479 27672 35488
rect 27620 35445 27629 35479
rect 27629 35445 27663 35479
rect 27663 35445 27672 35479
rect 27620 35436 27672 35445
rect 31392 35504 31444 35556
rect 33508 35683 33560 35692
rect 33508 35649 33517 35683
rect 33517 35649 33551 35683
rect 33551 35649 33560 35683
rect 33508 35640 33560 35649
rect 33600 35572 33652 35624
rect 36084 35615 36136 35624
rect 36084 35581 36093 35615
rect 36093 35581 36127 35615
rect 36127 35581 36136 35615
rect 36084 35572 36136 35581
rect 36360 35615 36412 35624
rect 36360 35581 36369 35615
rect 36369 35581 36403 35615
rect 36403 35581 36412 35615
rect 36360 35572 36412 35581
rect 37096 35572 37148 35624
rect 39396 35615 39448 35624
rect 39396 35581 39405 35615
rect 39405 35581 39439 35615
rect 39439 35581 39448 35615
rect 39396 35572 39448 35581
rect 38844 35504 38896 35556
rect 40960 35572 41012 35624
rect 31852 35436 31904 35488
rect 31944 35479 31996 35488
rect 31944 35445 31953 35479
rect 31953 35445 31987 35479
rect 31987 35445 31996 35479
rect 31944 35436 31996 35445
rect 33140 35436 33192 35488
rect 34428 35436 34480 35488
rect 39396 35436 39448 35488
rect 39856 35436 39908 35488
rect 40132 35436 40184 35488
rect 42616 35436 42668 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5080 35028 5132 35080
rect 5540 35232 5592 35284
rect 6092 35232 6144 35284
rect 7656 35275 7708 35284
rect 7656 35241 7665 35275
rect 7665 35241 7699 35275
rect 7699 35241 7708 35275
rect 7656 35232 7708 35241
rect 5448 35164 5500 35216
rect 5540 35028 5592 35080
rect 7472 35207 7524 35216
rect 7472 35173 7481 35207
rect 7481 35173 7515 35207
rect 7515 35173 7524 35207
rect 14280 35232 14332 35284
rect 15568 35232 15620 35284
rect 16212 35232 16264 35284
rect 7472 35164 7524 35173
rect 8484 35164 8536 35216
rect 6736 35096 6788 35148
rect 8300 35096 8352 35148
rect 7380 35028 7432 35080
rect 6736 34892 6788 34944
rect 7564 34960 7616 35012
rect 8852 35028 8904 35080
rect 8944 35071 8996 35080
rect 8944 35037 8953 35071
rect 8953 35037 8987 35071
rect 8987 35037 8996 35071
rect 8944 35028 8996 35037
rect 12256 35096 12308 35148
rect 18604 35232 18656 35284
rect 23756 35232 23808 35284
rect 25964 35232 26016 35284
rect 31944 35232 31996 35284
rect 8668 34892 8720 34944
rect 9404 35028 9456 35080
rect 11060 35028 11112 35080
rect 12624 35028 12676 35080
rect 16856 35096 16908 35148
rect 16948 35096 17000 35148
rect 20260 35096 20312 35148
rect 26424 35139 26476 35148
rect 18420 35028 18472 35080
rect 18880 35071 18932 35080
rect 18880 35037 18889 35071
rect 18889 35037 18923 35071
rect 18923 35037 18932 35071
rect 18880 35028 18932 35037
rect 20628 35028 20680 35080
rect 17316 35003 17368 35012
rect 17316 34969 17325 35003
rect 17325 34969 17359 35003
rect 17359 34969 17368 35003
rect 17316 34960 17368 34969
rect 12256 34892 12308 34944
rect 14832 34892 14884 34944
rect 15752 34935 15804 34944
rect 15752 34901 15761 34935
rect 15761 34901 15795 34935
rect 15795 34901 15804 34935
rect 15752 34892 15804 34901
rect 16212 34892 16264 34944
rect 22744 34960 22796 35012
rect 25044 35071 25096 35080
rect 25044 35037 25053 35071
rect 25053 35037 25087 35071
rect 25087 35037 25096 35071
rect 25044 35028 25096 35037
rect 25688 35028 25740 35080
rect 26424 35105 26433 35139
rect 26433 35105 26467 35139
rect 26467 35105 26476 35139
rect 26424 35096 26476 35105
rect 31760 35071 31812 35080
rect 31760 35037 31769 35071
rect 31769 35037 31803 35071
rect 31803 35037 31812 35071
rect 31760 35028 31812 35037
rect 34428 35096 34480 35148
rect 36360 35232 36412 35284
rect 39580 35232 39632 35284
rect 39948 35232 40000 35284
rect 40960 35232 41012 35284
rect 41144 35275 41196 35284
rect 41144 35241 41153 35275
rect 41153 35241 41187 35275
rect 41187 35241 41196 35275
rect 41144 35232 41196 35241
rect 39856 35207 39908 35216
rect 39856 35173 39865 35207
rect 39865 35173 39899 35207
rect 39899 35173 39908 35207
rect 39856 35164 39908 35173
rect 40132 35164 40184 35216
rect 38752 35139 38804 35148
rect 38752 35105 38761 35139
rect 38761 35105 38795 35139
rect 38795 35105 38804 35139
rect 38752 35096 38804 35105
rect 32036 35028 32088 35080
rect 35808 35028 35860 35080
rect 39120 35071 39172 35080
rect 39120 35037 39129 35071
rect 39129 35037 39163 35071
rect 39163 35037 39172 35071
rect 39120 35028 39172 35037
rect 32404 34960 32456 35012
rect 19340 34892 19392 34944
rect 22560 34892 22612 34944
rect 24032 34892 24084 34944
rect 24492 34935 24544 34944
rect 24492 34901 24501 34935
rect 24501 34901 24535 34935
rect 24535 34901 24544 34935
rect 24492 34892 24544 34901
rect 27620 34892 27672 34944
rect 35348 34892 35400 34944
rect 36176 35003 36228 35012
rect 36176 34969 36185 35003
rect 36185 34969 36219 35003
rect 36219 34969 36228 35003
rect 36176 34960 36228 34969
rect 36912 34960 36964 35012
rect 39764 35028 39816 35080
rect 42708 35139 42760 35148
rect 42708 35105 42717 35139
rect 42717 35105 42751 35139
rect 42751 35105 42760 35139
rect 42708 35096 42760 35105
rect 40868 35071 40920 35080
rect 40868 35037 40877 35071
rect 40877 35037 40911 35071
rect 40911 35037 40920 35071
rect 40868 35028 40920 35037
rect 42248 35028 42300 35080
rect 43444 35028 43496 35080
rect 36544 34892 36596 34944
rect 37648 34935 37700 34944
rect 37648 34901 37657 34935
rect 37657 34901 37691 34935
rect 37691 34901 37700 34935
rect 37648 34892 37700 34901
rect 39488 34935 39540 34944
rect 39488 34901 39497 34935
rect 39497 34901 39531 34935
rect 39531 34901 39540 34935
rect 39488 34892 39540 34901
rect 42064 34960 42116 35012
rect 42156 34892 42208 34944
rect 43260 34935 43312 34944
rect 43260 34901 43269 34935
rect 43269 34901 43303 34935
rect 43303 34901 43312 34935
rect 43260 34892 43312 34901
rect 43720 34892 43772 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 5632 34731 5684 34740
rect 5632 34697 5641 34731
rect 5641 34697 5675 34731
rect 5675 34697 5684 34731
rect 5632 34688 5684 34697
rect 6000 34688 6052 34740
rect 6092 34688 6144 34740
rect 6644 34688 6696 34740
rect 6736 34731 6788 34740
rect 6736 34697 6745 34731
rect 6745 34697 6779 34731
rect 6779 34697 6788 34731
rect 6736 34688 6788 34697
rect 7472 34688 7524 34740
rect 8300 34731 8352 34740
rect 8300 34697 8309 34731
rect 8309 34697 8343 34731
rect 8343 34697 8352 34731
rect 8300 34688 8352 34697
rect 8668 34688 8720 34740
rect 9404 34688 9456 34740
rect 13452 34688 13504 34740
rect 6184 34620 6236 34672
rect 6368 34595 6420 34604
rect 6368 34561 6377 34595
rect 6377 34561 6411 34595
rect 6411 34561 6420 34595
rect 6368 34552 6420 34561
rect 6460 34552 6512 34604
rect 6644 34595 6696 34604
rect 6644 34561 6653 34595
rect 6653 34561 6687 34595
rect 6687 34561 6696 34595
rect 6644 34552 6696 34561
rect 8484 34552 8536 34604
rect 8852 34552 8904 34604
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 11060 34620 11112 34672
rect 11520 34595 11572 34604
rect 11520 34561 11529 34595
rect 11529 34561 11563 34595
rect 11563 34561 11572 34595
rect 11520 34552 11572 34561
rect 12624 34620 12676 34672
rect 12532 34595 12584 34604
rect 12532 34561 12541 34595
rect 12541 34561 12575 34595
rect 12575 34561 12584 34595
rect 12532 34552 12584 34561
rect 12716 34595 12768 34604
rect 12716 34561 12725 34595
rect 12725 34561 12759 34595
rect 12759 34561 12768 34595
rect 12716 34552 12768 34561
rect 12808 34552 12860 34604
rect 13084 34552 13136 34604
rect 15660 34688 15712 34740
rect 16212 34731 16264 34740
rect 16212 34697 16221 34731
rect 16221 34697 16255 34731
rect 16255 34697 16264 34731
rect 16212 34688 16264 34697
rect 16856 34688 16908 34740
rect 17316 34688 17368 34740
rect 16488 34620 16540 34672
rect 16580 34620 16632 34672
rect 17132 34552 17184 34604
rect 17224 34595 17276 34604
rect 17224 34561 17233 34595
rect 17233 34561 17267 34595
rect 17267 34561 17276 34595
rect 17224 34552 17276 34561
rect 18788 34688 18840 34740
rect 18880 34731 18932 34740
rect 18880 34697 18889 34731
rect 18889 34697 18923 34731
rect 18923 34697 18932 34731
rect 18880 34688 18932 34697
rect 19248 34688 19300 34740
rect 5080 34484 5132 34536
rect 5448 34484 5500 34536
rect 8668 34527 8720 34536
rect 8668 34493 8677 34527
rect 8677 34493 8711 34527
rect 8711 34493 8720 34527
rect 8668 34484 8720 34493
rect 13360 34484 13412 34536
rect 14740 34527 14792 34536
rect 14740 34493 14749 34527
rect 14749 34493 14783 34527
rect 14783 34493 14792 34527
rect 14740 34484 14792 34493
rect 18052 34484 18104 34536
rect 19248 34595 19300 34604
rect 19248 34561 19257 34595
rect 19257 34561 19291 34595
rect 19291 34561 19300 34595
rect 19248 34552 19300 34561
rect 8852 34459 8904 34468
rect 8852 34425 8861 34459
rect 8861 34425 8895 34459
rect 8895 34425 8904 34459
rect 8852 34416 8904 34425
rect 19064 34416 19116 34468
rect 22008 34484 22060 34536
rect 22560 34416 22612 34468
rect 26056 34688 26108 34740
rect 27896 34688 27948 34740
rect 30196 34688 30248 34740
rect 33508 34688 33560 34740
rect 24492 34663 24544 34672
rect 24492 34629 24501 34663
rect 24501 34629 24535 34663
rect 24535 34629 24544 34663
rect 24492 34620 24544 34629
rect 25228 34620 25280 34672
rect 28448 34620 28500 34672
rect 23572 34552 23624 34604
rect 23664 34552 23716 34604
rect 24032 34595 24084 34604
rect 24032 34561 24041 34595
rect 24041 34561 24075 34595
rect 24075 34561 24084 34595
rect 24032 34552 24084 34561
rect 27252 34595 27304 34604
rect 27252 34561 27261 34595
rect 27261 34561 27295 34595
rect 27295 34561 27304 34595
rect 27252 34552 27304 34561
rect 27528 34595 27580 34604
rect 27528 34561 27537 34595
rect 27537 34561 27571 34595
rect 27571 34561 27580 34595
rect 27528 34552 27580 34561
rect 26792 34484 26844 34536
rect 34612 34620 34664 34672
rect 35348 34663 35400 34672
rect 35348 34629 35357 34663
rect 35357 34629 35391 34663
rect 35391 34629 35400 34663
rect 35348 34620 35400 34629
rect 36084 34688 36136 34740
rect 36176 34620 36228 34672
rect 37648 34688 37700 34740
rect 37924 34688 37976 34740
rect 39120 34688 39172 34740
rect 36544 34620 36596 34672
rect 42064 34688 42116 34740
rect 42248 34731 42300 34740
rect 42248 34697 42257 34731
rect 42257 34697 42291 34731
rect 42291 34697 42300 34731
rect 42248 34688 42300 34697
rect 30748 34595 30800 34604
rect 30748 34561 30757 34595
rect 30757 34561 30791 34595
rect 30791 34561 30800 34595
rect 30748 34552 30800 34561
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 32312 34484 32364 34536
rect 35440 34595 35492 34604
rect 35440 34561 35449 34595
rect 35449 34561 35483 34595
rect 35483 34561 35492 34595
rect 35440 34552 35492 34561
rect 35348 34484 35400 34536
rect 35808 34484 35860 34536
rect 36268 34484 36320 34536
rect 36544 34484 36596 34536
rect 31024 34416 31076 34468
rect 9036 34348 9088 34400
rect 9312 34391 9364 34400
rect 9312 34357 9342 34391
rect 9342 34357 9364 34391
rect 9312 34348 9364 34357
rect 10784 34391 10836 34400
rect 10784 34357 10793 34391
rect 10793 34357 10827 34391
rect 10827 34357 10836 34391
rect 10784 34348 10836 34357
rect 11612 34391 11664 34400
rect 11612 34357 11621 34391
rect 11621 34357 11655 34391
rect 11655 34357 11664 34391
rect 11612 34348 11664 34357
rect 12992 34391 13044 34400
rect 12992 34357 13001 34391
rect 13001 34357 13035 34391
rect 13035 34357 13044 34391
rect 12992 34348 13044 34357
rect 23480 34391 23532 34400
rect 23480 34357 23489 34391
rect 23489 34357 23523 34391
rect 23523 34357 23532 34391
rect 23480 34348 23532 34357
rect 23572 34391 23624 34400
rect 23572 34357 23581 34391
rect 23581 34357 23615 34391
rect 23615 34357 23624 34391
rect 23572 34348 23624 34357
rect 26884 34348 26936 34400
rect 27068 34348 27120 34400
rect 36268 34348 36320 34400
rect 38016 34552 38068 34604
rect 38384 34595 38436 34604
rect 38384 34561 38393 34595
rect 38393 34561 38427 34595
rect 38427 34561 38436 34595
rect 38384 34552 38436 34561
rect 39488 34552 39540 34604
rect 41420 34552 41472 34604
rect 42156 34552 42208 34604
rect 42708 34688 42760 34740
rect 42616 34620 42668 34672
rect 43720 34620 43772 34672
rect 44272 34595 44324 34604
rect 44272 34561 44281 34595
rect 44281 34561 44315 34595
rect 44315 34561 44324 34595
rect 44272 34552 44324 34561
rect 37648 34391 37700 34400
rect 37648 34357 37657 34391
rect 37657 34357 37691 34391
rect 37691 34357 37700 34391
rect 37648 34348 37700 34357
rect 38476 34348 38528 34400
rect 39396 34348 39448 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5540 34144 5592 34196
rect 9312 34144 9364 34196
rect 12716 34144 12768 34196
rect 12900 34144 12952 34196
rect 6092 34076 6144 34128
rect 12624 34076 12676 34128
rect 14740 34187 14792 34196
rect 14740 34153 14749 34187
rect 14749 34153 14783 34187
rect 14783 34153 14792 34187
rect 14740 34144 14792 34153
rect 15660 34144 15712 34196
rect 17960 34144 18012 34196
rect 21548 34144 21600 34196
rect 25044 34187 25096 34196
rect 25044 34153 25053 34187
rect 25053 34153 25087 34187
rect 25087 34153 25096 34187
rect 25044 34144 25096 34153
rect 28448 34187 28500 34196
rect 28448 34153 28457 34187
rect 28457 34153 28491 34187
rect 28491 34153 28500 34187
rect 28448 34144 28500 34153
rect 30748 34144 30800 34196
rect 30932 34144 30984 34196
rect 31116 34187 31168 34196
rect 31116 34153 31125 34187
rect 31125 34153 31159 34187
rect 31159 34153 31168 34187
rect 31116 34144 31168 34153
rect 31392 34144 31444 34196
rect 32864 34187 32916 34196
rect 32864 34153 32873 34187
rect 32873 34153 32907 34187
rect 32907 34153 32916 34187
rect 32864 34144 32916 34153
rect 33324 34144 33376 34196
rect 33784 34144 33836 34196
rect 34060 34187 34112 34196
rect 34060 34153 34069 34187
rect 34069 34153 34103 34187
rect 34103 34153 34112 34187
rect 34060 34144 34112 34153
rect 35348 34144 35400 34196
rect 39488 34144 39540 34196
rect 43444 34144 43496 34196
rect 6184 33940 6236 33992
rect 10784 34008 10836 34060
rect 11336 34008 11388 34060
rect 6368 33940 6420 33992
rect 8852 33940 8904 33992
rect 9036 33940 9088 33992
rect 12348 34008 12400 34060
rect 5540 33804 5592 33856
rect 8944 33804 8996 33856
rect 11612 33983 11664 33992
rect 11612 33949 11621 33983
rect 11621 33949 11655 33983
rect 11655 33949 11664 33983
rect 11612 33940 11664 33949
rect 11796 33940 11848 33992
rect 12072 33983 12124 33992
rect 12072 33949 12081 33983
rect 12081 33949 12115 33983
rect 12115 33949 12124 33983
rect 12072 33940 12124 33949
rect 12256 33940 12308 33992
rect 12532 33983 12584 33992
rect 12532 33949 12541 33983
rect 12541 33949 12575 33983
rect 12575 33949 12584 33983
rect 12532 33940 12584 33949
rect 11980 33915 12032 33924
rect 11980 33881 11989 33915
rect 11989 33881 12023 33915
rect 12023 33881 12032 33915
rect 11980 33872 12032 33881
rect 19340 34076 19392 34128
rect 20812 34076 20864 34128
rect 22284 34076 22336 34128
rect 30564 34076 30616 34128
rect 31024 34076 31076 34128
rect 12992 34008 13044 34060
rect 13176 33983 13228 33992
rect 13176 33949 13185 33983
rect 13185 33949 13219 33983
rect 13219 33949 13228 33983
rect 13176 33940 13228 33949
rect 13452 33983 13504 33992
rect 13452 33949 13461 33983
rect 13461 33949 13495 33983
rect 13495 33949 13504 33983
rect 13452 33940 13504 33949
rect 12808 33872 12860 33924
rect 13084 33872 13136 33924
rect 11796 33804 11848 33856
rect 12164 33804 12216 33856
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 12440 33804 12492 33856
rect 14188 33940 14240 33992
rect 14464 33940 14516 33992
rect 14924 33983 14976 33992
rect 14924 33949 14933 33983
rect 14933 33949 14967 33983
rect 14967 33949 14976 33983
rect 14924 33940 14976 33949
rect 15844 33940 15896 33992
rect 20904 34008 20956 34060
rect 22560 34051 22612 34060
rect 22560 34017 22569 34051
rect 22569 34017 22603 34051
rect 22603 34017 22612 34051
rect 22560 34008 22612 34017
rect 23480 34008 23532 34060
rect 23572 34008 23624 34060
rect 24676 34008 24728 34060
rect 24768 34008 24820 34060
rect 27068 34008 27120 34060
rect 21456 33940 21508 33992
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 24860 33983 24912 33992
rect 24860 33949 24874 33983
rect 24874 33949 24908 33983
rect 24908 33949 24912 33983
rect 24860 33940 24912 33949
rect 26056 33940 26108 33992
rect 26608 33940 26660 33992
rect 17592 33872 17644 33924
rect 19156 33872 19208 33924
rect 23020 33872 23072 33924
rect 13820 33847 13872 33856
rect 13820 33813 13829 33847
rect 13829 33813 13863 33847
rect 13863 33813 13872 33847
rect 13820 33804 13872 33813
rect 20352 33847 20404 33856
rect 20352 33813 20361 33847
rect 20361 33813 20395 33847
rect 20395 33813 20404 33847
rect 20352 33804 20404 33813
rect 22744 33847 22796 33856
rect 22744 33813 22753 33847
rect 22753 33813 22787 33847
rect 22787 33813 22796 33847
rect 22744 33804 22796 33813
rect 23572 33872 23624 33924
rect 26424 33872 26476 33924
rect 27436 33872 27488 33924
rect 23388 33847 23440 33856
rect 23388 33813 23397 33847
rect 23397 33813 23431 33847
rect 23431 33813 23440 33847
rect 23388 33804 23440 33813
rect 24584 33804 24636 33856
rect 29828 33804 29880 33856
rect 33508 34008 33560 34060
rect 37280 34076 37332 34128
rect 31392 33983 31444 33992
rect 31392 33949 31401 33983
rect 31401 33949 31435 33983
rect 31435 33949 31444 33983
rect 31392 33940 31444 33949
rect 32312 33983 32364 33992
rect 32312 33949 32321 33983
rect 32321 33949 32355 33983
rect 32355 33949 32364 33983
rect 32312 33940 32364 33949
rect 32496 33983 32548 33992
rect 32496 33949 32505 33983
rect 32505 33949 32539 33983
rect 32539 33949 32548 33983
rect 32496 33940 32548 33949
rect 32588 33983 32640 33992
rect 32588 33949 32597 33983
rect 32597 33949 32631 33983
rect 32631 33949 32640 33983
rect 32588 33940 32640 33949
rect 33692 33983 33744 33992
rect 33692 33949 33701 33983
rect 33701 33949 33735 33983
rect 33735 33949 33744 33983
rect 33692 33940 33744 33949
rect 32772 33915 32824 33924
rect 32772 33881 32781 33915
rect 32781 33881 32815 33915
rect 32815 33881 32824 33915
rect 32772 33872 32824 33881
rect 34796 34051 34848 34060
rect 34796 34017 34805 34051
rect 34805 34017 34839 34051
rect 34839 34017 34848 34051
rect 34796 34008 34848 34017
rect 38476 34008 38528 34060
rect 39856 33940 39908 33992
rect 40868 34008 40920 34060
rect 41420 34051 41472 34060
rect 41420 34017 41429 34051
rect 41429 34017 41463 34051
rect 41463 34017 41472 34051
rect 41420 34008 41472 34017
rect 31208 33804 31260 33856
rect 32036 33847 32088 33856
rect 32036 33813 32045 33847
rect 32045 33813 32079 33847
rect 32079 33813 32088 33847
rect 32036 33804 32088 33813
rect 32128 33847 32180 33856
rect 32128 33813 32137 33847
rect 32137 33813 32171 33847
rect 32171 33813 32180 33847
rect 32128 33804 32180 33813
rect 33048 33804 33100 33856
rect 33232 33804 33284 33856
rect 34428 33847 34480 33856
rect 34428 33813 34437 33847
rect 34437 33813 34471 33847
rect 34471 33813 34480 33847
rect 34428 33804 34480 33813
rect 36912 33847 36964 33856
rect 36912 33813 36921 33847
rect 36921 33813 36955 33847
rect 36955 33813 36964 33847
rect 36912 33804 36964 33813
rect 38752 33804 38804 33856
rect 39764 33804 39816 33856
rect 40408 33847 40460 33856
rect 40408 33813 40417 33847
rect 40417 33813 40451 33847
rect 40451 33813 40460 33847
rect 40408 33804 40460 33813
rect 40592 33847 40644 33856
rect 40592 33813 40601 33847
rect 40601 33813 40635 33847
rect 40635 33813 40644 33847
rect 42064 33983 42116 33992
rect 42064 33949 42073 33983
rect 42073 33949 42107 33983
rect 42107 33949 42116 33983
rect 42064 33940 42116 33949
rect 42156 33940 42208 33992
rect 43260 33940 43312 33992
rect 44640 34008 44692 34060
rect 40592 33804 40644 33813
rect 43904 33804 43956 33856
rect 44088 33847 44140 33856
rect 44088 33813 44097 33847
rect 44097 33813 44131 33847
rect 44131 33813 44140 33847
rect 44088 33804 44140 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 6368 33643 6420 33652
rect 6368 33609 6377 33643
rect 6377 33609 6411 33643
rect 6411 33609 6420 33643
rect 6368 33600 6420 33609
rect 8392 33600 8444 33652
rect 11980 33600 12032 33652
rect 12716 33600 12768 33652
rect 5172 33464 5224 33516
rect 13820 33600 13872 33652
rect 14924 33600 14976 33652
rect 15752 33600 15804 33652
rect 20260 33643 20312 33652
rect 20260 33609 20269 33643
rect 20269 33609 20303 33643
rect 20303 33609 20312 33643
rect 20260 33600 20312 33609
rect 20720 33600 20772 33652
rect 21088 33600 21140 33652
rect 22008 33643 22060 33652
rect 22008 33609 22017 33643
rect 22017 33609 22051 33643
rect 22051 33609 22060 33643
rect 22008 33600 22060 33609
rect 3884 33439 3936 33448
rect 3884 33405 3893 33439
rect 3893 33405 3927 33439
rect 3927 33405 3936 33439
rect 3884 33396 3936 33405
rect 4620 33396 4672 33448
rect 11612 33464 11664 33516
rect 11888 33507 11940 33516
rect 11888 33473 11897 33507
rect 11897 33473 11931 33507
rect 11931 33473 11940 33507
rect 11888 33464 11940 33473
rect 11980 33507 12032 33516
rect 11980 33473 11989 33507
rect 11989 33473 12023 33507
rect 12023 33473 12032 33507
rect 11980 33464 12032 33473
rect 25044 33600 25096 33652
rect 23388 33532 23440 33584
rect 23572 33532 23624 33584
rect 26240 33600 26292 33652
rect 26424 33600 26476 33652
rect 12256 33464 12308 33516
rect 12624 33464 12676 33516
rect 12992 33464 13044 33516
rect 8024 33396 8076 33448
rect 9772 33328 9824 33380
rect 12164 33328 12216 33380
rect 12440 33328 12492 33380
rect 5816 33303 5868 33312
rect 5816 33269 5825 33303
rect 5825 33269 5859 33303
rect 5859 33269 5868 33303
rect 5816 33260 5868 33269
rect 12072 33260 12124 33312
rect 13268 33328 13320 33380
rect 15844 33464 15896 33516
rect 16028 33328 16080 33380
rect 12900 33303 12952 33312
rect 12900 33269 12909 33303
rect 12909 33269 12943 33303
rect 12943 33269 12952 33303
rect 12900 33260 12952 33269
rect 13176 33260 13228 33312
rect 13820 33260 13872 33312
rect 15936 33260 15988 33312
rect 18420 33507 18472 33516
rect 18420 33473 18429 33507
rect 18429 33473 18463 33507
rect 18463 33473 18472 33507
rect 18420 33464 18472 33473
rect 17132 33439 17184 33448
rect 17132 33405 17141 33439
rect 17141 33405 17175 33439
rect 17175 33405 17184 33439
rect 17132 33396 17184 33405
rect 17316 33396 17368 33448
rect 17224 33260 17276 33312
rect 18512 33439 18564 33448
rect 18512 33405 18521 33439
rect 18521 33405 18555 33439
rect 18555 33405 18564 33439
rect 18512 33396 18564 33405
rect 19340 33507 19392 33516
rect 19340 33473 19349 33507
rect 19349 33473 19383 33507
rect 19383 33473 19392 33507
rect 19340 33464 19392 33473
rect 19432 33464 19484 33516
rect 20168 33464 20220 33516
rect 19524 33260 19576 33312
rect 20628 33396 20680 33448
rect 20628 33303 20680 33312
rect 20628 33269 20637 33303
rect 20637 33269 20671 33303
rect 20671 33269 20680 33303
rect 20628 33260 20680 33269
rect 21272 33464 21324 33516
rect 21456 33507 21508 33516
rect 21456 33473 21465 33507
rect 21465 33473 21499 33507
rect 21499 33473 21508 33507
rect 21456 33464 21508 33473
rect 21548 33464 21600 33516
rect 26516 33532 26568 33584
rect 27896 33600 27948 33652
rect 28540 33600 28592 33652
rect 31392 33600 31444 33652
rect 32036 33600 32088 33652
rect 32312 33643 32364 33652
rect 32312 33609 32339 33643
rect 32339 33609 32364 33643
rect 32312 33600 32364 33609
rect 33416 33600 33468 33652
rect 27528 33532 27580 33584
rect 29828 33532 29880 33584
rect 32128 33532 32180 33584
rect 32496 33575 32548 33584
rect 32496 33541 32505 33575
rect 32505 33541 32539 33575
rect 32539 33541 32548 33575
rect 32496 33532 32548 33541
rect 33692 33600 33744 33652
rect 26884 33464 26936 33516
rect 29000 33464 29052 33516
rect 20904 33396 20956 33448
rect 20996 33439 21048 33448
rect 20996 33405 21005 33439
rect 21005 33405 21039 33439
rect 21039 33405 21048 33439
rect 20996 33396 21048 33405
rect 24768 33328 24820 33380
rect 21180 33260 21232 33312
rect 23848 33303 23900 33312
rect 23848 33269 23857 33303
rect 23857 33269 23891 33303
rect 23891 33269 23900 33303
rect 23848 33260 23900 33269
rect 26608 33396 26660 33448
rect 28632 33396 28684 33448
rect 26424 33328 26476 33380
rect 31576 33396 31628 33448
rect 32772 33507 32824 33516
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 33048 33507 33100 33516
rect 33048 33473 33057 33507
rect 33057 33473 33091 33507
rect 33091 33473 33100 33507
rect 33048 33464 33100 33473
rect 33232 33507 33284 33516
rect 33232 33473 33241 33507
rect 33241 33473 33275 33507
rect 33275 33473 33284 33507
rect 33232 33464 33284 33473
rect 33324 33507 33376 33516
rect 33324 33473 33333 33507
rect 33333 33473 33367 33507
rect 33367 33473 33376 33507
rect 33324 33464 33376 33473
rect 33784 33507 33836 33516
rect 33784 33473 33798 33507
rect 33798 33473 33832 33507
rect 33832 33473 33836 33507
rect 34428 33600 34480 33652
rect 34520 33600 34572 33652
rect 33784 33464 33836 33473
rect 36544 33600 36596 33652
rect 36912 33600 36964 33652
rect 37280 33643 37332 33652
rect 37280 33609 37289 33643
rect 37289 33609 37323 33643
rect 37323 33609 37332 33643
rect 37280 33600 37332 33609
rect 39764 33600 39816 33652
rect 40868 33600 40920 33652
rect 42064 33600 42116 33652
rect 35348 33464 35400 33516
rect 35440 33464 35492 33516
rect 38292 33532 38344 33584
rect 36820 33464 36872 33516
rect 33876 33328 33928 33380
rect 34704 33328 34756 33380
rect 32588 33260 32640 33312
rect 33048 33260 33100 33312
rect 38384 33260 38436 33312
rect 40132 33396 40184 33448
rect 39764 33260 39816 33312
rect 43444 33532 43496 33584
rect 43904 33575 43956 33584
rect 43904 33541 43913 33575
rect 43913 33541 43947 33575
rect 43947 33541 43956 33575
rect 43904 33532 43956 33541
rect 42524 33260 42576 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 33099 4672 33108
rect 4620 33065 4629 33099
rect 4629 33065 4663 33099
rect 4663 33065 4672 33099
rect 4620 33056 4672 33065
rect 5816 33056 5868 33108
rect 8300 33056 8352 33108
rect 9128 33056 9180 33108
rect 12072 33056 12124 33108
rect 12624 33056 12676 33108
rect 13820 33031 13872 33040
rect 13820 32997 13829 33031
rect 13829 32997 13863 33031
rect 13863 32997 13872 33031
rect 13820 32988 13872 32997
rect 6920 32963 6972 32972
rect 6920 32929 6929 32963
rect 6929 32929 6963 32963
rect 6963 32929 6972 32963
rect 6920 32920 6972 32929
rect 12440 32920 12492 32972
rect 3884 32852 3936 32904
rect 5540 32852 5592 32904
rect 5724 32852 5776 32904
rect 6828 32784 6880 32836
rect 12900 32852 12952 32904
rect 13360 32852 13412 32904
rect 14188 32852 14240 32904
rect 14556 33056 14608 33108
rect 17224 33056 17276 33108
rect 17592 33056 17644 33108
rect 18512 33056 18564 33108
rect 19432 33099 19484 33108
rect 19432 33065 19441 33099
rect 19441 33065 19475 33099
rect 19475 33065 19484 33099
rect 19432 33056 19484 33065
rect 20168 33056 20220 33108
rect 14464 32920 14516 32972
rect 15660 32963 15712 32972
rect 15660 32929 15669 32963
rect 15669 32929 15703 32963
rect 15703 32929 15712 32963
rect 15660 32920 15712 32929
rect 20996 32988 21048 33040
rect 21272 33031 21324 33040
rect 21272 32997 21281 33031
rect 21281 32997 21315 33031
rect 21315 32997 21324 33031
rect 21272 32988 21324 32997
rect 7196 32827 7248 32836
rect 7196 32793 7205 32827
rect 7205 32793 7239 32827
rect 7239 32793 7248 32827
rect 7196 32784 7248 32793
rect 8484 32784 8536 32836
rect 9312 32784 9364 32836
rect 15936 32827 15988 32836
rect 15936 32793 15945 32827
rect 15945 32793 15979 32827
rect 15979 32793 15988 32827
rect 15936 32784 15988 32793
rect 17224 32784 17276 32836
rect 20352 32920 20404 32972
rect 17868 32852 17920 32904
rect 18880 32852 18932 32904
rect 18420 32784 18472 32836
rect 11704 32716 11756 32768
rect 20076 32852 20128 32904
rect 20812 32852 20864 32904
rect 21640 32852 21692 32904
rect 21364 32784 21416 32836
rect 22284 33056 22336 33108
rect 22744 33056 22796 33108
rect 23848 33056 23900 33108
rect 24676 33056 24728 33108
rect 26516 33099 26568 33108
rect 26516 33065 26525 33099
rect 26525 33065 26559 33099
rect 26559 33065 26568 33099
rect 26516 33056 26568 33065
rect 28632 33099 28684 33108
rect 28632 33065 28641 33099
rect 28641 33065 28675 33099
rect 28675 33065 28684 33099
rect 28632 33056 28684 33065
rect 34704 33056 34756 33108
rect 34796 33056 34848 33108
rect 23572 32895 23624 32904
rect 23572 32861 23581 32895
rect 23581 32861 23615 32895
rect 23615 32861 23624 32895
rect 23572 32852 23624 32861
rect 23664 32852 23716 32904
rect 26332 32988 26384 33040
rect 33876 32988 33928 33040
rect 35348 33056 35400 33108
rect 38292 33056 38344 33108
rect 40132 33099 40184 33108
rect 40132 33065 40141 33099
rect 40141 33065 40175 33099
rect 40175 33065 40184 33099
rect 40132 33056 40184 33065
rect 27252 32920 27304 32972
rect 20260 32716 20312 32768
rect 21180 32716 21232 32768
rect 24860 32895 24912 32904
rect 24860 32861 24874 32895
rect 24874 32861 24908 32895
rect 24908 32861 24912 32895
rect 24860 32852 24912 32861
rect 26424 32852 26476 32904
rect 24676 32827 24728 32836
rect 24676 32793 24685 32827
rect 24685 32793 24719 32827
rect 24719 32793 24728 32827
rect 24676 32784 24728 32793
rect 25688 32784 25740 32836
rect 27160 32895 27212 32904
rect 27160 32861 27169 32895
rect 27169 32861 27203 32895
rect 27203 32861 27212 32895
rect 27160 32852 27212 32861
rect 31392 32895 31444 32904
rect 31392 32861 31401 32895
rect 31401 32861 31435 32895
rect 31435 32861 31444 32895
rect 31392 32852 31444 32861
rect 31208 32784 31260 32836
rect 33508 32852 33560 32904
rect 34520 32920 34572 32972
rect 34060 32852 34112 32904
rect 40408 32988 40460 33040
rect 44088 32988 44140 33040
rect 43352 32963 43404 32972
rect 43352 32929 43361 32963
rect 43361 32929 43395 32963
rect 43395 32929 43404 32963
rect 43352 32920 43404 32929
rect 43536 32920 43588 32972
rect 35256 32895 35308 32904
rect 35256 32861 35265 32895
rect 35265 32861 35299 32895
rect 35299 32861 35308 32895
rect 35256 32852 35308 32861
rect 37648 32895 37700 32904
rect 37648 32861 37657 32895
rect 37657 32861 37691 32895
rect 37691 32861 37700 32895
rect 37648 32852 37700 32861
rect 38568 32852 38620 32904
rect 40592 32852 40644 32904
rect 39396 32784 39448 32836
rect 40040 32827 40092 32836
rect 40040 32793 40049 32827
rect 40049 32793 40083 32827
rect 40083 32793 40092 32827
rect 40040 32784 40092 32793
rect 24952 32716 25004 32768
rect 30932 32759 30984 32768
rect 30932 32725 30941 32759
rect 30941 32725 30975 32759
rect 30975 32725 30984 32759
rect 30932 32716 30984 32725
rect 31392 32759 31444 32768
rect 31392 32725 31401 32759
rect 31401 32725 31435 32759
rect 31435 32725 31444 32759
rect 31392 32716 31444 32725
rect 33416 32716 33468 32768
rect 34520 32716 34572 32768
rect 43812 32759 43864 32768
rect 43812 32725 43821 32759
rect 43821 32725 43855 32759
rect 43855 32725 43864 32759
rect 43812 32716 43864 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 7196 32512 7248 32564
rect 8024 32512 8076 32564
rect 7012 32444 7064 32496
rect 7288 32444 7340 32496
rect 16580 32512 16632 32564
rect 6184 32419 6236 32428
rect 6184 32385 6193 32419
rect 6193 32385 6227 32419
rect 6227 32385 6236 32419
rect 6184 32376 6236 32385
rect 8024 32419 8076 32428
rect 8024 32385 8033 32419
rect 8033 32385 8067 32419
rect 8067 32385 8076 32419
rect 8024 32376 8076 32385
rect 7656 32308 7708 32360
rect 9128 32376 9180 32428
rect 11612 32376 11664 32428
rect 11704 32376 11756 32428
rect 17960 32444 18012 32496
rect 5172 32240 5224 32292
rect 8392 32240 8444 32292
rect 9772 32308 9824 32360
rect 14648 32308 14700 32360
rect 15660 32376 15712 32428
rect 16304 32419 16356 32428
rect 16304 32385 16313 32419
rect 16313 32385 16347 32419
rect 16347 32385 16356 32419
rect 16304 32376 16356 32385
rect 22284 32512 22336 32564
rect 26608 32512 26660 32564
rect 27896 32555 27948 32564
rect 27896 32521 27905 32555
rect 27905 32521 27939 32555
rect 27939 32521 27948 32555
rect 27896 32512 27948 32521
rect 33324 32512 33376 32564
rect 35256 32512 35308 32564
rect 43812 32512 43864 32564
rect 26424 32444 26476 32496
rect 26240 32376 26292 32428
rect 23664 32308 23716 32360
rect 25136 32351 25188 32360
rect 25136 32317 25145 32351
rect 25145 32317 25179 32351
rect 25179 32317 25188 32351
rect 25136 32308 25188 32317
rect 5816 32172 5868 32224
rect 8484 32172 8536 32224
rect 10968 32215 11020 32224
rect 10968 32181 10977 32215
rect 10977 32181 11011 32215
rect 11011 32181 11020 32215
rect 10968 32172 11020 32181
rect 11336 32172 11388 32224
rect 15844 32172 15896 32224
rect 18696 32240 18748 32292
rect 24400 32240 24452 32292
rect 31208 32444 31260 32496
rect 31392 32444 31444 32496
rect 33600 32444 33652 32496
rect 34520 32487 34572 32496
rect 30932 32419 30984 32428
rect 30932 32385 30941 32419
rect 30941 32385 30975 32419
rect 30975 32385 30984 32419
rect 30932 32376 30984 32385
rect 29736 32308 29788 32360
rect 30656 32308 30708 32360
rect 31300 32308 31352 32360
rect 32128 32308 32180 32360
rect 34520 32453 34529 32487
rect 34529 32453 34563 32487
rect 34563 32453 34572 32487
rect 34520 32444 34572 32453
rect 34704 32376 34756 32428
rect 42432 32376 42484 32428
rect 36176 32308 36228 32360
rect 26884 32240 26936 32292
rect 17592 32172 17644 32224
rect 18052 32172 18104 32224
rect 18512 32215 18564 32224
rect 18512 32181 18521 32215
rect 18521 32181 18555 32215
rect 18555 32181 18564 32215
rect 18512 32172 18564 32181
rect 20812 32172 20864 32224
rect 21180 32172 21232 32224
rect 22192 32215 22244 32224
rect 22192 32181 22201 32215
rect 22201 32181 22235 32215
rect 22235 32181 22244 32215
rect 22192 32172 22244 32181
rect 30564 32172 30616 32224
rect 31024 32215 31076 32224
rect 31024 32181 31033 32215
rect 31033 32181 31067 32215
rect 31067 32181 31076 32215
rect 31024 32172 31076 32181
rect 31208 32240 31260 32292
rect 31576 32240 31628 32292
rect 33784 32240 33836 32292
rect 35348 32172 35400 32224
rect 38016 32172 38068 32224
rect 42248 32215 42300 32224
rect 42248 32181 42257 32215
rect 42257 32181 42291 32215
rect 42291 32181 42300 32215
rect 42248 32172 42300 32181
rect 43352 32215 43404 32224
rect 43352 32181 43361 32215
rect 43361 32181 43395 32215
rect 43395 32181 43404 32215
rect 43352 32172 43404 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7196 32011 7248 32020
rect 7196 31977 7205 32011
rect 7205 31977 7239 32011
rect 7239 31977 7248 32011
rect 7196 31968 7248 31977
rect 7748 31968 7800 32020
rect 10968 31968 11020 32020
rect 11244 31968 11296 32020
rect 11336 31968 11388 32020
rect 3884 31832 3936 31884
rect 5816 31832 5868 31884
rect 6920 31832 6972 31884
rect 8024 31943 8076 31952
rect 8024 31909 8033 31943
rect 8033 31909 8067 31943
rect 8067 31909 8076 31943
rect 8024 31900 8076 31909
rect 5172 31696 5224 31748
rect 7104 31696 7156 31748
rect 7748 31696 7800 31748
rect 8576 31764 8628 31816
rect 8300 31739 8352 31748
rect 8300 31705 8309 31739
rect 8309 31705 8343 31739
rect 8343 31705 8352 31739
rect 8300 31696 8352 31705
rect 8392 31696 8444 31748
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 9312 31696 9364 31748
rect 9588 31739 9640 31748
rect 9588 31705 9597 31739
rect 9597 31705 9631 31739
rect 9631 31705 9640 31739
rect 9588 31696 9640 31705
rect 8576 31628 8628 31680
rect 9036 31671 9088 31680
rect 9036 31637 9045 31671
rect 9045 31637 9079 31671
rect 9079 31637 9088 31671
rect 9036 31628 9088 31637
rect 11244 31807 11296 31816
rect 11244 31773 11253 31807
rect 11253 31773 11287 31807
rect 11287 31773 11296 31807
rect 11244 31764 11296 31773
rect 16304 31968 16356 32020
rect 20260 31968 20312 32020
rect 24860 31968 24912 32020
rect 25136 31968 25188 32020
rect 27160 31968 27212 32020
rect 30564 31968 30616 32020
rect 30656 31968 30708 32020
rect 32128 31968 32180 32020
rect 34060 32011 34112 32020
rect 34060 31977 34069 32011
rect 34069 31977 34103 32011
rect 34103 31977 34112 32011
rect 34060 31968 34112 31977
rect 37464 31968 37516 32020
rect 39488 31968 39540 32020
rect 12532 31900 12584 31952
rect 15752 31900 15804 31952
rect 16396 31900 16448 31952
rect 19432 31900 19484 31952
rect 20812 31900 20864 31952
rect 12164 31764 12216 31816
rect 11980 31739 12032 31748
rect 11980 31705 11989 31739
rect 11989 31705 12023 31739
rect 12023 31705 12032 31739
rect 12440 31764 12492 31816
rect 15200 31832 15252 31884
rect 11980 31696 12032 31705
rect 11704 31628 11756 31680
rect 14372 31628 14424 31680
rect 15292 31764 15344 31816
rect 17316 31875 17368 31884
rect 17316 31841 17325 31875
rect 17325 31841 17359 31875
rect 17359 31841 17368 31875
rect 17316 31832 17368 31841
rect 20720 31832 20772 31884
rect 15476 31807 15528 31816
rect 15476 31773 15485 31807
rect 15485 31773 15519 31807
rect 15519 31773 15528 31807
rect 15476 31764 15528 31773
rect 15568 31696 15620 31748
rect 15108 31628 15160 31680
rect 18512 31764 18564 31816
rect 20444 31764 20496 31816
rect 19340 31696 19392 31748
rect 20168 31696 20220 31748
rect 24952 31832 25004 31884
rect 24032 31764 24084 31816
rect 24860 31807 24912 31816
rect 24860 31773 24867 31807
rect 24867 31773 24912 31807
rect 24860 31764 24912 31773
rect 29736 31783 29746 31816
rect 29746 31783 29780 31816
rect 29780 31783 29788 31816
rect 29736 31764 29788 31783
rect 31760 31900 31812 31952
rect 41052 31943 41104 31952
rect 29920 31807 29972 31816
rect 29920 31773 29929 31807
rect 29929 31773 29963 31807
rect 29963 31773 29972 31807
rect 29920 31764 29972 31773
rect 30104 31764 30156 31816
rect 30472 31764 30524 31816
rect 21548 31696 21600 31748
rect 24584 31696 24636 31748
rect 26424 31696 26476 31748
rect 19984 31671 20036 31680
rect 19984 31637 19993 31671
rect 19993 31637 20027 31671
rect 20027 31637 20036 31671
rect 19984 31628 20036 31637
rect 20076 31628 20128 31680
rect 20260 31671 20312 31680
rect 20260 31637 20269 31671
rect 20269 31637 20303 31671
rect 20303 31637 20312 31671
rect 20260 31628 20312 31637
rect 20444 31671 20496 31680
rect 20444 31637 20453 31671
rect 20453 31637 20487 31671
rect 20487 31637 20496 31671
rect 20444 31628 20496 31637
rect 20536 31671 20588 31680
rect 20536 31637 20545 31671
rect 20545 31637 20579 31671
rect 20579 31637 20588 31671
rect 20536 31628 20588 31637
rect 20996 31628 21048 31680
rect 24492 31628 24544 31680
rect 27068 31628 27120 31680
rect 29552 31671 29604 31680
rect 29552 31637 29561 31671
rect 29561 31637 29595 31671
rect 29595 31637 29604 31671
rect 29552 31628 29604 31637
rect 30748 31696 30800 31748
rect 31024 31764 31076 31816
rect 31116 31764 31168 31816
rect 31300 31764 31352 31816
rect 31576 31807 31628 31816
rect 31576 31773 31585 31807
rect 31585 31773 31619 31807
rect 31619 31773 31628 31807
rect 31576 31764 31628 31773
rect 31944 31875 31996 31884
rect 31944 31841 31953 31875
rect 31953 31841 31987 31875
rect 31987 31841 31996 31875
rect 31944 31832 31996 31841
rect 38016 31832 38068 31884
rect 38384 31832 38436 31884
rect 31760 31696 31812 31748
rect 36544 31764 36596 31816
rect 33232 31696 33284 31748
rect 34336 31696 34388 31748
rect 34428 31739 34480 31748
rect 34428 31705 34437 31739
rect 34437 31705 34471 31739
rect 34471 31705 34480 31739
rect 34428 31696 34480 31705
rect 36820 31807 36872 31816
rect 36820 31773 36853 31807
rect 36853 31773 36872 31807
rect 41052 31909 41061 31943
rect 41061 31909 41095 31943
rect 41095 31909 41104 31943
rect 41052 31900 41104 31909
rect 38568 31832 38620 31884
rect 39672 31832 39724 31884
rect 39764 31832 39816 31884
rect 40040 31832 40092 31884
rect 36820 31764 36872 31773
rect 37464 31696 37516 31748
rect 36820 31628 36872 31680
rect 38108 31628 38160 31680
rect 40776 31807 40828 31816
rect 40776 31773 40785 31807
rect 40785 31773 40819 31807
rect 40819 31773 40828 31807
rect 40776 31764 40828 31773
rect 42892 31968 42944 32020
rect 42524 31875 42576 31884
rect 42524 31841 42533 31875
rect 42533 31841 42567 31875
rect 42567 31841 42576 31875
rect 42524 31832 42576 31841
rect 43352 31832 43404 31884
rect 44272 31875 44324 31884
rect 44272 31841 44281 31875
rect 44281 31841 44315 31875
rect 44315 31841 44324 31875
rect 44272 31832 44324 31841
rect 42156 31807 42208 31816
rect 42156 31773 42165 31807
rect 42165 31773 42199 31807
rect 42199 31773 42208 31807
rect 42156 31764 42208 31773
rect 39672 31696 39724 31748
rect 40684 31696 40736 31748
rect 43444 31696 43496 31748
rect 39212 31628 39264 31680
rect 39764 31628 39816 31680
rect 41144 31628 41196 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 6276 31424 6328 31476
rect 8484 31467 8536 31476
rect 8484 31433 8493 31467
rect 8493 31433 8527 31467
rect 8527 31433 8536 31467
rect 8484 31424 8536 31433
rect 9036 31424 9088 31476
rect 9588 31424 9640 31476
rect 11980 31467 12032 31476
rect 11980 31433 11989 31467
rect 11989 31433 12023 31467
rect 12023 31433 12032 31467
rect 11980 31424 12032 31433
rect 5540 31288 5592 31340
rect 7380 31356 7432 31408
rect 8116 31399 8168 31408
rect 8116 31365 8125 31399
rect 8125 31365 8159 31399
rect 8159 31365 8168 31399
rect 8116 31356 8168 31365
rect 7104 31288 7156 31340
rect 8300 31152 8352 31204
rect 8576 31288 8628 31340
rect 8668 31288 8720 31340
rect 9128 31331 9180 31340
rect 9128 31297 9137 31331
rect 9137 31297 9171 31331
rect 9171 31297 9180 31331
rect 9128 31288 9180 31297
rect 11796 31288 11848 31340
rect 12624 31288 12676 31340
rect 14004 31424 14056 31476
rect 14464 31424 14516 31476
rect 19340 31424 19392 31476
rect 19616 31424 19668 31476
rect 21272 31424 21324 31476
rect 24860 31424 24912 31476
rect 25044 31424 25096 31476
rect 32864 31424 32916 31476
rect 14556 31399 14608 31408
rect 14556 31365 14565 31399
rect 14565 31365 14599 31399
rect 14599 31365 14608 31399
rect 14556 31356 14608 31365
rect 14648 31399 14700 31408
rect 14648 31365 14657 31399
rect 14657 31365 14691 31399
rect 14691 31365 14700 31399
rect 14648 31356 14700 31365
rect 13176 31220 13228 31272
rect 13728 31263 13780 31272
rect 13728 31229 13737 31263
rect 13737 31229 13771 31263
rect 13771 31229 13780 31263
rect 13728 31220 13780 31229
rect 14188 31331 14240 31340
rect 14188 31297 14197 31331
rect 14197 31297 14231 31331
rect 14231 31297 14240 31331
rect 14188 31288 14240 31297
rect 14280 31288 14332 31340
rect 14832 31331 14884 31340
rect 14832 31297 14840 31331
rect 14840 31297 14874 31331
rect 14874 31297 14884 31331
rect 14832 31288 14884 31297
rect 14924 31331 14976 31340
rect 14924 31297 14933 31331
rect 14933 31297 14967 31331
rect 14967 31297 14976 31331
rect 14924 31288 14976 31297
rect 15568 31356 15620 31408
rect 15292 31331 15344 31340
rect 15292 31297 15301 31331
rect 15301 31297 15335 31331
rect 15335 31297 15344 31331
rect 15292 31288 15344 31297
rect 15752 31331 15804 31340
rect 15752 31297 15761 31331
rect 15761 31297 15795 31331
rect 15795 31297 15804 31331
rect 15752 31288 15804 31297
rect 15844 31288 15896 31340
rect 6000 31127 6052 31136
rect 6000 31093 6009 31127
rect 6009 31093 6043 31127
rect 6043 31093 6052 31127
rect 6000 31084 6052 31093
rect 6920 31084 6972 31136
rect 7748 31084 7800 31136
rect 15660 31263 15712 31272
rect 15660 31229 15669 31263
rect 15669 31229 15703 31263
rect 15703 31229 15712 31263
rect 15660 31220 15712 31229
rect 16028 31263 16080 31272
rect 16028 31229 16037 31263
rect 16037 31229 16071 31263
rect 16071 31229 16080 31263
rect 16028 31220 16080 31229
rect 15476 31152 15528 31204
rect 16488 31288 16540 31340
rect 19248 31288 19300 31340
rect 13820 31127 13872 31136
rect 13820 31093 13829 31127
rect 13829 31093 13863 31127
rect 13863 31093 13872 31127
rect 13820 31084 13872 31093
rect 14280 31127 14332 31136
rect 14280 31093 14289 31127
rect 14289 31093 14323 31127
rect 14323 31093 14332 31127
rect 14280 31084 14332 31093
rect 14556 31084 14608 31136
rect 15016 31127 15068 31136
rect 15016 31093 15025 31127
rect 15025 31093 15059 31127
rect 15059 31093 15068 31127
rect 15016 31084 15068 31093
rect 15384 31084 15436 31136
rect 19432 31152 19484 31204
rect 18420 31084 18472 31136
rect 19340 31084 19392 31136
rect 20628 31356 20680 31408
rect 20812 31399 20864 31408
rect 20812 31365 20821 31399
rect 20821 31365 20855 31399
rect 20855 31365 20864 31399
rect 20812 31356 20864 31365
rect 21548 31356 21600 31408
rect 23572 31356 23624 31408
rect 26424 31399 26476 31408
rect 26424 31365 26433 31399
rect 26433 31365 26467 31399
rect 26467 31365 26476 31399
rect 26424 31356 26476 31365
rect 21088 31331 21140 31340
rect 21088 31297 21097 31331
rect 21097 31297 21131 31331
rect 21131 31297 21140 31331
rect 21088 31288 21140 31297
rect 21364 31331 21416 31340
rect 21364 31297 21373 31331
rect 21373 31297 21407 31331
rect 21407 31297 21416 31331
rect 21364 31288 21416 31297
rect 19800 31152 19852 31204
rect 20812 31220 20864 31272
rect 21548 31263 21600 31272
rect 21548 31229 21557 31263
rect 21557 31229 21591 31263
rect 21591 31229 21600 31263
rect 21548 31220 21600 31229
rect 22560 31263 22612 31272
rect 22560 31229 22569 31263
rect 22569 31229 22603 31263
rect 22603 31229 22612 31263
rect 22560 31220 22612 31229
rect 22836 31263 22888 31272
rect 22836 31229 22845 31263
rect 22845 31229 22879 31263
rect 22879 31229 22888 31263
rect 22836 31220 22888 31229
rect 25872 31263 25924 31272
rect 25872 31229 25881 31263
rect 25881 31229 25915 31263
rect 25915 31229 25924 31263
rect 25872 31220 25924 31229
rect 27528 31356 27580 31408
rect 28632 31356 28684 31408
rect 30012 31356 30064 31408
rect 26792 31288 26844 31340
rect 28264 31331 28316 31340
rect 28264 31297 28273 31331
rect 28273 31297 28307 31331
rect 28307 31297 28316 31331
rect 28264 31288 28316 31297
rect 30380 31331 30432 31340
rect 30380 31297 30389 31331
rect 30389 31297 30423 31331
rect 30423 31297 30432 31331
rect 30380 31288 30432 31297
rect 30472 31331 30524 31340
rect 30472 31297 30481 31331
rect 30481 31297 30515 31331
rect 30515 31297 30524 31331
rect 30472 31288 30524 31297
rect 31116 31356 31168 31408
rect 31576 31356 31628 31408
rect 31392 31288 31444 31340
rect 35348 31424 35400 31476
rect 35808 31424 35860 31476
rect 27436 31220 27488 31272
rect 20076 31152 20128 31204
rect 20904 31084 20956 31136
rect 23848 31084 23900 31136
rect 26056 31127 26108 31136
rect 26056 31093 26065 31127
rect 26065 31093 26099 31127
rect 26099 31093 26108 31127
rect 26056 31084 26108 31093
rect 29552 31220 29604 31272
rect 33232 31331 33284 31340
rect 33232 31297 33241 31331
rect 33241 31297 33275 31331
rect 33275 31297 33284 31331
rect 33232 31288 33284 31297
rect 33508 31220 33560 31272
rect 29644 31152 29696 31204
rect 31944 31152 31996 31204
rect 32680 31152 32732 31204
rect 29276 31084 29328 31136
rect 32772 31127 32824 31136
rect 32772 31093 32781 31127
rect 32781 31093 32815 31127
rect 32815 31093 32824 31127
rect 32772 31084 32824 31093
rect 32864 31084 32916 31136
rect 38752 31399 38804 31408
rect 38752 31365 38761 31399
rect 38761 31365 38795 31399
rect 38795 31365 38804 31399
rect 38752 31356 38804 31365
rect 39212 31356 39264 31408
rect 38016 31288 38068 31340
rect 38476 31331 38528 31340
rect 38476 31297 38485 31331
rect 38485 31297 38519 31331
rect 38519 31297 38528 31331
rect 38476 31288 38528 31297
rect 42156 31424 42208 31476
rect 42432 31467 42484 31476
rect 42432 31433 42441 31467
rect 42441 31433 42475 31467
rect 42475 31433 42484 31467
rect 42432 31424 42484 31433
rect 42892 31467 42944 31476
rect 42892 31433 42901 31467
rect 42901 31433 42935 31467
rect 42935 31433 42944 31467
rect 42892 31424 42944 31433
rect 40684 31356 40736 31408
rect 42800 31331 42852 31340
rect 42800 31297 42809 31331
rect 42809 31297 42843 31331
rect 42843 31297 42852 31331
rect 42800 31288 42852 31297
rect 38384 31220 38436 31272
rect 39764 31152 39816 31204
rect 37924 31084 37976 31136
rect 40040 31084 40092 31136
rect 40592 31263 40644 31272
rect 40592 31229 40601 31263
rect 40601 31229 40635 31263
rect 40635 31229 40644 31263
rect 40592 31220 40644 31229
rect 43168 31220 43220 31272
rect 40776 31084 40828 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3884 30880 3936 30932
rect 6000 30880 6052 30932
rect 8300 30880 8352 30932
rect 13820 30880 13872 30932
rect 14280 30923 14332 30932
rect 14280 30889 14304 30923
rect 14304 30889 14332 30923
rect 14280 30880 14332 30889
rect 14372 30923 14424 30932
rect 14372 30889 14381 30923
rect 14381 30889 14415 30923
rect 14415 30889 14424 30923
rect 14372 30880 14424 30889
rect 14556 30923 14608 30932
rect 14556 30889 14565 30923
rect 14565 30889 14599 30923
rect 14599 30889 14608 30923
rect 14556 30880 14608 30889
rect 15016 30880 15068 30932
rect 17316 30880 17368 30932
rect 19248 30880 19300 30932
rect 19524 30923 19576 30932
rect 19524 30889 19533 30923
rect 19533 30889 19567 30923
rect 19567 30889 19576 30923
rect 19524 30880 19576 30889
rect 19708 30880 19760 30932
rect 7196 30744 7248 30796
rect 5172 30676 5224 30728
rect 5632 30676 5684 30728
rect 6092 30719 6144 30728
rect 6092 30685 6101 30719
rect 6101 30685 6135 30719
rect 6135 30685 6144 30719
rect 6092 30676 6144 30685
rect 5816 30651 5868 30660
rect 5816 30617 5825 30651
rect 5825 30617 5859 30651
rect 5859 30617 5868 30651
rect 5816 30608 5868 30617
rect 13084 30812 13136 30864
rect 13176 30812 13228 30864
rect 7564 30719 7616 30728
rect 7564 30685 7573 30719
rect 7573 30685 7607 30719
rect 7607 30685 7616 30719
rect 7564 30676 7616 30685
rect 7380 30608 7432 30660
rect 8208 30719 8260 30728
rect 8208 30685 8217 30719
rect 8217 30685 8251 30719
rect 8251 30685 8260 30719
rect 8208 30676 8260 30685
rect 7748 30651 7800 30660
rect 7748 30617 7757 30651
rect 7757 30617 7791 30651
rect 7791 30617 7800 30651
rect 7748 30608 7800 30617
rect 10508 30719 10560 30728
rect 10508 30685 10517 30719
rect 10517 30685 10551 30719
rect 10551 30685 10560 30719
rect 10508 30676 10560 30685
rect 11704 30719 11756 30728
rect 11704 30685 11714 30719
rect 11714 30685 11748 30719
rect 11748 30685 11756 30719
rect 11704 30676 11756 30685
rect 12072 30719 12124 30728
rect 12072 30685 12086 30719
rect 12086 30685 12120 30719
rect 12120 30685 12124 30719
rect 12072 30676 12124 30685
rect 7932 30583 7984 30592
rect 7932 30549 7941 30583
rect 7941 30549 7975 30583
rect 7975 30549 7984 30583
rect 7932 30540 7984 30549
rect 11980 30540 12032 30592
rect 12440 30608 12492 30660
rect 12900 30676 12952 30728
rect 13544 30812 13596 30864
rect 15752 30812 15804 30864
rect 19616 30812 19668 30864
rect 13544 30719 13596 30728
rect 13544 30685 13553 30719
rect 13553 30685 13587 30719
rect 13587 30685 13596 30719
rect 13544 30676 13596 30685
rect 13820 30676 13872 30728
rect 12348 30583 12400 30592
rect 12348 30549 12357 30583
rect 12357 30549 12391 30583
rect 12391 30549 12400 30583
rect 12348 30540 12400 30549
rect 12992 30540 13044 30592
rect 13360 30540 13412 30592
rect 13912 30540 13964 30592
rect 14188 30744 14240 30796
rect 14280 30744 14332 30796
rect 14832 30744 14884 30796
rect 15384 30787 15436 30796
rect 15384 30753 15393 30787
rect 15393 30753 15427 30787
rect 15427 30753 15436 30787
rect 15384 30744 15436 30753
rect 17132 30744 17184 30796
rect 19892 30812 19944 30864
rect 20076 30855 20128 30864
rect 20076 30821 20085 30855
rect 20085 30821 20119 30855
rect 20119 30821 20128 30855
rect 20076 30812 20128 30821
rect 20536 30880 20588 30932
rect 21088 30880 21140 30932
rect 21180 30880 21232 30932
rect 22836 30880 22888 30932
rect 25872 30880 25924 30932
rect 26056 30880 26108 30932
rect 29000 30880 29052 30932
rect 30012 30880 30064 30932
rect 14096 30651 14148 30660
rect 14096 30617 14105 30651
rect 14105 30617 14139 30651
rect 14139 30617 14148 30651
rect 14096 30608 14148 30617
rect 14648 30608 14700 30660
rect 15660 30676 15712 30728
rect 16488 30608 16540 30660
rect 18328 30719 18380 30728
rect 18328 30685 18337 30719
rect 18337 30685 18371 30719
rect 18371 30685 18380 30719
rect 18328 30676 18380 30685
rect 18420 30676 18472 30728
rect 18788 30719 18840 30728
rect 18788 30685 18797 30719
rect 18797 30685 18831 30719
rect 18831 30685 18840 30719
rect 18788 30676 18840 30685
rect 18972 30719 19024 30728
rect 18972 30685 18981 30719
rect 18981 30685 19015 30719
rect 19015 30685 19024 30719
rect 18972 30676 19024 30685
rect 19708 30719 19760 30728
rect 19708 30685 19717 30719
rect 19717 30685 19751 30719
rect 19751 30685 19760 30719
rect 19708 30676 19760 30685
rect 20076 30676 20128 30728
rect 20260 30676 20312 30728
rect 20260 30540 20312 30592
rect 20536 30719 20588 30728
rect 20536 30685 20545 30719
rect 20545 30685 20579 30719
rect 20579 30685 20588 30719
rect 20536 30676 20588 30685
rect 20812 30719 20864 30728
rect 20812 30685 20821 30719
rect 20821 30685 20855 30719
rect 20855 30685 20864 30719
rect 20812 30676 20864 30685
rect 21180 30719 21232 30728
rect 21180 30685 21189 30719
rect 21189 30685 21223 30719
rect 21223 30685 21232 30719
rect 21180 30676 21232 30685
rect 21272 30676 21324 30728
rect 22008 30719 22060 30728
rect 22008 30685 22017 30719
rect 22017 30685 22051 30719
rect 22051 30685 22060 30719
rect 22008 30676 22060 30685
rect 23756 30744 23808 30796
rect 24124 30787 24176 30796
rect 24124 30753 24133 30787
rect 24133 30753 24167 30787
rect 24167 30753 24176 30787
rect 24124 30744 24176 30753
rect 29276 30855 29328 30864
rect 29276 30821 29285 30855
rect 29285 30821 29319 30855
rect 29319 30821 29328 30855
rect 29276 30812 29328 30821
rect 32036 30880 32088 30932
rect 34428 30880 34480 30932
rect 35992 30880 36044 30932
rect 38384 30880 38436 30932
rect 38752 30880 38804 30932
rect 40592 30923 40644 30932
rect 40592 30889 40601 30923
rect 40601 30889 40635 30923
rect 40635 30889 40644 30923
rect 40592 30880 40644 30889
rect 41052 30880 41104 30932
rect 41328 30880 41380 30932
rect 42156 30880 42208 30932
rect 28264 30744 28316 30796
rect 33692 30787 33744 30796
rect 33692 30753 33701 30787
rect 33701 30753 33735 30787
rect 33735 30753 33744 30787
rect 33692 30744 33744 30753
rect 23940 30676 23992 30728
rect 29460 30676 29512 30728
rect 30380 30719 30432 30728
rect 30380 30685 30389 30719
rect 30389 30685 30423 30719
rect 30423 30685 30432 30719
rect 30380 30676 30432 30685
rect 31300 30719 31352 30728
rect 31300 30685 31309 30719
rect 31309 30685 31343 30719
rect 31343 30685 31352 30719
rect 31300 30676 31352 30685
rect 34244 30744 34296 30796
rect 20812 30540 20864 30592
rect 20904 30540 20956 30592
rect 26700 30608 26752 30660
rect 22468 30540 22520 30592
rect 23388 30540 23440 30592
rect 26240 30540 26292 30592
rect 27804 30651 27856 30660
rect 27804 30617 27813 30651
rect 27813 30617 27847 30651
rect 27847 30617 27856 30651
rect 27804 30608 27856 30617
rect 34152 30676 34204 30728
rect 31852 30608 31904 30660
rect 32036 30608 32088 30660
rect 29092 30540 29144 30592
rect 33232 30608 33284 30660
rect 36820 30812 36872 30864
rect 34796 30787 34848 30796
rect 34796 30753 34805 30787
rect 34805 30753 34839 30787
rect 34839 30753 34848 30787
rect 34796 30744 34848 30753
rect 35348 30676 35400 30728
rect 37924 30719 37976 30728
rect 37924 30685 37933 30719
rect 37933 30685 37967 30719
rect 37967 30685 37976 30719
rect 37924 30676 37976 30685
rect 38200 30719 38252 30728
rect 38200 30685 38209 30719
rect 38209 30685 38243 30719
rect 38243 30685 38252 30719
rect 38200 30676 38252 30685
rect 38752 30676 38804 30728
rect 33140 30583 33192 30592
rect 33140 30549 33149 30583
rect 33149 30549 33183 30583
rect 33183 30549 33192 30583
rect 33140 30540 33192 30549
rect 35256 30583 35308 30592
rect 35256 30549 35265 30583
rect 35265 30549 35299 30583
rect 35299 30549 35308 30583
rect 35256 30540 35308 30549
rect 35716 30608 35768 30660
rect 36452 30540 36504 30592
rect 38016 30608 38068 30660
rect 38568 30651 38620 30660
rect 38568 30617 38577 30651
rect 38577 30617 38611 30651
rect 38611 30617 38620 30651
rect 38568 30608 38620 30617
rect 41144 30787 41196 30796
rect 41144 30753 41153 30787
rect 41153 30753 41187 30787
rect 41187 30753 41196 30787
rect 41144 30744 41196 30753
rect 42800 30744 42852 30796
rect 43352 30744 43404 30796
rect 39488 30719 39540 30728
rect 39488 30685 39497 30719
rect 39497 30685 39531 30719
rect 39531 30685 39540 30719
rect 39488 30676 39540 30685
rect 39764 30676 39816 30728
rect 38844 30583 38896 30592
rect 38844 30549 38853 30583
rect 38853 30549 38887 30583
rect 38887 30549 38896 30583
rect 38844 30540 38896 30549
rect 39120 30540 39172 30592
rect 39304 30651 39356 30660
rect 39304 30617 39313 30651
rect 39313 30617 39347 30651
rect 39347 30617 39356 30651
rect 39304 30608 39356 30617
rect 40500 30676 40552 30728
rect 40776 30676 40828 30728
rect 41972 30676 42024 30728
rect 43444 30676 43496 30728
rect 41880 30540 41932 30592
rect 43076 30540 43128 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5632 30379 5684 30388
rect 5632 30345 5641 30379
rect 5641 30345 5675 30379
rect 5675 30345 5684 30379
rect 5632 30336 5684 30345
rect 6092 30379 6144 30388
rect 6092 30345 6101 30379
rect 6101 30345 6135 30379
rect 6135 30345 6144 30379
rect 6092 30336 6144 30345
rect 7380 30379 7432 30388
rect 7380 30345 7389 30379
rect 7389 30345 7423 30379
rect 7423 30345 7432 30379
rect 7380 30336 7432 30345
rect 7564 30336 7616 30388
rect 7840 30336 7892 30388
rect 5448 30039 5500 30048
rect 5448 30005 5457 30039
rect 5457 30005 5491 30039
rect 5491 30005 5500 30039
rect 5448 29996 5500 30005
rect 12072 30336 12124 30388
rect 9312 30200 9364 30252
rect 9496 30200 9548 30252
rect 12164 30268 12216 30320
rect 12900 30336 12952 30388
rect 13636 30336 13688 30388
rect 13728 30336 13780 30388
rect 5724 30132 5776 30184
rect 6000 30132 6052 30184
rect 6920 30132 6972 30184
rect 8024 30175 8076 30184
rect 8024 30141 8033 30175
rect 8033 30141 8067 30175
rect 8067 30141 8076 30175
rect 8024 30132 8076 30141
rect 7564 30064 7616 30116
rect 12716 30200 12768 30252
rect 12256 30132 12308 30184
rect 12992 30200 13044 30252
rect 13176 30268 13228 30320
rect 18788 30336 18840 30388
rect 19432 30336 19484 30388
rect 15200 30311 15252 30320
rect 15200 30277 15209 30311
rect 15209 30277 15243 30311
rect 15243 30277 15252 30311
rect 15200 30268 15252 30277
rect 18420 30268 18472 30320
rect 5816 29996 5868 30048
rect 12624 30107 12676 30116
rect 12624 30073 12633 30107
rect 12633 30073 12667 30107
rect 12667 30073 12676 30107
rect 12624 30064 12676 30073
rect 13820 30132 13872 30184
rect 14004 30175 14056 30184
rect 14004 30141 14013 30175
rect 14013 30141 14047 30175
rect 14047 30141 14056 30175
rect 14004 30132 14056 30141
rect 15568 30132 15620 30184
rect 11612 29996 11664 30048
rect 11888 29996 11940 30048
rect 13360 30039 13412 30048
rect 13360 30005 13369 30039
rect 13369 30005 13403 30039
rect 13403 30005 13412 30039
rect 13360 29996 13412 30005
rect 18052 30200 18104 30252
rect 18328 30200 18380 30252
rect 16580 30132 16632 30184
rect 18052 30064 18104 30116
rect 17316 29996 17368 30048
rect 17960 29996 18012 30048
rect 18972 30243 19024 30252
rect 18972 30209 18973 30243
rect 18973 30209 19007 30243
rect 19007 30209 19024 30243
rect 18972 30200 19024 30209
rect 19340 30243 19392 30252
rect 19340 30209 19349 30243
rect 19349 30209 19383 30243
rect 19383 30209 19392 30243
rect 19340 30200 19392 30209
rect 19800 30200 19852 30252
rect 20168 30268 20220 30320
rect 20444 30336 20496 30388
rect 22008 30336 22060 30388
rect 23940 30379 23992 30388
rect 23940 30345 23949 30379
rect 23949 30345 23983 30379
rect 23983 30345 23992 30379
rect 23940 30336 23992 30345
rect 26700 30336 26752 30388
rect 27436 30336 27488 30388
rect 27804 30336 27856 30388
rect 26424 30268 26476 30320
rect 27528 30268 27580 30320
rect 30104 30336 30156 30388
rect 29092 30268 29144 30320
rect 20352 30243 20404 30252
rect 20352 30209 20386 30243
rect 20386 30209 20404 30243
rect 20904 30243 20956 30252
rect 20352 30200 20404 30209
rect 19432 30175 19484 30184
rect 19432 30141 19441 30175
rect 19441 30141 19475 30175
rect 19475 30141 19484 30175
rect 19432 30132 19484 30141
rect 19984 30064 20036 30116
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 23572 30200 23624 30252
rect 20628 30132 20680 30184
rect 20812 30175 20864 30184
rect 20812 30141 20821 30175
rect 20821 30141 20855 30175
rect 20855 30141 20864 30175
rect 20812 30132 20864 30141
rect 20996 30175 21048 30184
rect 20996 30141 21005 30175
rect 21005 30141 21039 30175
rect 21039 30141 21048 30175
rect 20996 30132 21048 30141
rect 18604 30039 18656 30048
rect 18604 30005 18613 30039
rect 18613 30005 18647 30039
rect 18647 30005 18656 30039
rect 18604 29996 18656 30005
rect 19432 29996 19484 30048
rect 22468 30175 22520 30184
rect 22468 30141 22477 30175
rect 22477 30141 22511 30175
rect 22511 30141 22520 30175
rect 22468 30132 22520 30141
rect 24400 30175 24452 30184
rect 24400 30141 24409 30175
rect 24409 30141 24443 30175
rect 24443 30141 24452 30175
rect 24400 30132 24452 30141
rect 24492 30132 24544 30184
rect 26424 30132 26476 30184
rect 27896 30200 27948 30252
rect 29000 30132 29052 30184
rect 29460 30311 29512 30320
rect 29460 30277 29469 30311
rect 29469 30277 29503 30311
rect 29503 30277 29512 30311
rect 29460 30268 29512 30277
rect 29184 30132 29236 30184
rect 29644 30243 29696 30252
rect 29644 30209 29653 30243
rect 29653 30209 29687 30243
rect 29687 30209 29696 30243
rect 29644 30200 29696 30209
rect 30196 30200 30248 30252
rect 23572 30064 23624 30116
rect 29736 30132 29788 30184
rect 31852 30336 31904 30388
rect 32680 30336 32732 30388
rect 32772 30336 32824 30388
rect 33140 30336 33192 30388
rect 33324 30379 33376 30388
rect 33324 30345 33326 30379
rect 33326 30345 33360 30379
rect 33360 30345 33376 30379
rect 33324 30336 33376 30345
rect 32588 30243 32640 30252
rect 32588 30209 32597 30243
rect 32597 30209 32631 30243
rect 32631 30209 32640 30243
rect 32588 30200 32640 30209
rect 34796 30336 34848 30388
rect 35256 30336 35308 30388
rect 35716 30336 35768 30388
rect 36728 30336 36780 30388
rect 38200 30336 38252 30388
rect 38476 30336 38528 30388
rect 33140 30243 33192 30252
rect 33140 30209 33149 30243
rect 33149 30209 33183 30243
rect 33183 30209 33192 30243
rect 33140 30200 33192 30209
rect 33692 30243 33744 30252
rect 33692 30209 33701 30243
rect 33701 30209 33735 30243
rect 33735 30209 33744 30243
rect 33692 30200 33744 30209
rect 34060 30243 34112 30252
rect 34060 30209 34069 30243
rect 34069 30209 34103 30243
rect 34103 30209 34112 30243
rect 34060 30200 34112 30209
rect 34244 30243 34296 30252
rect 34244 30209 34253 30243
rect 34253 30209 34287 30243
rect 34287 30209 34296 30243
rect 34244 30200 34296 30209
rect 34428 30243 34480 30252
rect 34428 30209 34437 30243
rect 34437 30209 34471 30243
rect 34471 30209 34480 30243
rect 34428 30200 34480 30209
rect 34152 30132 34204 30184
rect 35440 30243 35492 30252
rect 35440 30209 35449 30243
rect 35449 30209 35483 30243
rect 35483 30209 35492 30243
rect 35440 30200 35492 30209
rect 35992 30200 36044 30252
rect 36452 30243 36504 30252
rect 36452 30209 36461 30243
rect 36461 30209 36495 30243
rect 36495 30209 36504 30243
rect 36452 30200 36504 30209
rect 36544 30200 36596 30252
rect 37832 30243 37884 30252
rect 37832 30209 37841 30243
rect 37841 30209 37875 30243
rect 37875 30209 37884 30243
rect 37832 30200 37884 30209
rect 38844 30336 38896 30388
rect 40500 30336 40552 30388
rect 39120 30268 39172 30320
rect 36728 30175 36780 30184
rect 36728 30141 36737 30175
rect 36737 30141 36771 30175
rect 36771 30141 36780 30175
rect 36728 30132 36780 30141
rect 41880 30243 41932 30252
rect 41880 30209 41889 30243
rect 41889 30209 41923 30243
rect 41923 30209 41932 30243
rect 41880 30200 41932 30209
rect 43076 30379 43128 30388
rect 43076 30345 43085 30379
rect 43085 30345 43119 30379
rect 43119 30345 43128 30379
rect 43076 30336 43128 30345
rect 43168 30200 43220 30252
rect 39764 30132 39816 30184
rect 41144 30175 41196 30184
rect 41144 30141 41153 30175
rect 41153 30141 41187 30175
rect 41187 30141 41196 30175
rect 41144 30132 41196 30141
rect 42524 30175 42576 30184
rect 42524 30141 42533 30175
rect 42533 30141 42567 30175
rect 42567 30141 42576 30175
rect 42524 30132 42576 30141
rect 22560 29996 22612 30048
rect 23204 29996 23256 30048
rect 27620 29996 27672 30048
rect 32864 29996 32916 30048
rect 38016 30064 38068 30116
rect 33508 29996 33560 30048
rect 36912 29996 36964 30048
rect 38108 30039 38160 30048
rect 38108 30005 38117 30039
rect 38117 30005 38151 30039
rect 38151 30005 38160 30039
rect 38108 29996 38160 30005
rect 39212 29996 39264 30048
rect 40592 30039 40644 30048
rect 40592 30005 40601 30039
rect 40601 30005 40635 30039
rect 40635 30005 40644 30039
rect 40592 29996 40644 30005
rect 41052 29996 41104 30048
rect 41236 29996 41288 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3884 29792 3936 29844
rect 5448 29792 5500 29844
rect 7932 29792 7984 29844
rect 8024 29792 8076 29844
rect 12532 29792 12584 29844
rect 13360 29792 13412 29844
rect 13820 29792 13872 29844
rect 6000 29656 6052 29708
rect 10416 29724 10468 29776
rect 5172 29588 5224 29640
rect 4068 29563 4120 29572
rect 4068 29529 4077 29563
rect 4077 29529 4111 29563
rect 4111 29529 4120 29563
rect 4068 29520 4120 29529
rect 5724 29520 5776 29572
rect 7380 29588 7432 29640
rect 7656 29588 7708 29640
rect 8944 29699 8996 29708
rect 8944 29665 8953 29699
rect 8953 29665 8987 29699
rect 8987 29665 8996 29699
rect 8944 29656 8996 29665
rect 6184 29495 6236 29504
rect 6184 29461 6193 29495
rect 6193 29461 6227 29495
rect 6227 29461 6236 29495
rect 6184 29452 6236 29461
rect 6552 29563 6604 29572
rect 6552 29529 6561 29563
rect 6561 29529 6595 29563
rect 6595 29529 6604 29563
rect 6552 29520 6604 29529
rect 8208 29588 8260 29640
rect 11060 29588 11112 29640
rect 11520 29631 11572 29640
rect 11520 29597 11529 29631
rect 11529 29597 11563 29631
rect 11563 29597 11572 29631
rect 11520 29588 11572 29597
rect 11612 29631 11664 29640
rect 11612 29597 11622 29631
rect 11622 29597 11656 29631
rect 11656 29597 11664 29631
rect 11612 29588 11664 29597
rect 11796 29631 11848 29640
rect 11796 29597 11805 29631
rect 11805 29597 11839 29631
rect 11839 29597 11848 29631
rect 11796 29588 11848 29597
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 12624 29631 12676 29640
rect 12624 29597 12633 29631
rect 12633 29597 12667 29631
rect 12667 29597 12676 29631
rect 12624 29588 12676 29597
rect 18604 29792 18656 29844
rect 20812 29792 20864 29844
rect 21180 29792 21232 29844
rect 24400 29792 24452 29844
rect 26240 29792 26292 29844
rect 27620 29835 27672 29844
rect 27620 29801 27629 29835
rect 27629 29801 27663 29835
rect 27663 29801 27672 29835
rect 27620 29792 27672 29801
rect 34060 29792 34112 29844
rect 35440 29792 35492 29844
rect 35900 29792 35952 29844
rect 38568 29792 38620 29844
rect 41144 29792 41196 29844
rect 42524 29792 42576 29844
rect 15384 29656 15436 29708
rect 16580 29656 16632 29708
rect 17224 29656 17276 29708
rect 18236 29656 18288 29708
rect 19064 29656 19116 29708
rect 20260 29656 20312 29708
rect 20996 29656 21048 29708
rect 24124 29656 24176 29708
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 16028 29563 16080 29572
rect 16028 29529 16037 29563
rect 16037 29529 16071 29563
rect 16071 29529 16080 29563
rect 16028 29520 16080 29529
rect 17316 29520 17368 29572
rect 8852 29452 8904 29504
rect 11244 29452 11296 29504
rect 12992 29452 13044 29504
rect 14280 29452 14332 29504
rect 17500 29495 17552 29504
rect 17500 29461 17509 29495
rect 17509 29461 17543 29495
rect 17543 29461 17552 29495
rect 17500 29452 17552 29461
rect 17868 29495 17920 29504
rect 17868 29461 17877 29495
rect 17877 29461 17911 29495
rect 17911 29461 17920 29495
rect 17868 29452 17920 29461
rect 18328 29495 18380 29504
rect 18328 29461 18337 29495
rect 18337 29461 18371 29495
rect 18371 29461 18380 29495
rect 18328 29452 18380 29461
rect 20352 29452 20404 29504
rect 24492 29588 24544 29640
rect 27436 29631 27488 29640
rect 27436 29597 27445 29631
rect 27445 29597 27479 29631
rect 27479 29597 27488 29631
rect 27436 29588 27488 29597
rect 33968 29631 34020 29640
rect 33968 29597 33977 29631
rect 33977 29597 34011 29631
rect 34011 29597 34020 29631
rect 33968 29588 34020 29597
rect 34704 29588 34756 29640
rect 41236 29656 41288 29708
rect 43076 29656 43128 29708
rect 38752 29631 38804 29640
rect 38752 29597 38761 29631
rect 38761 29597 38795 29631
rect 38795 29597 38804 29631
rect 38752 29588 38804 29597
rect 39120 29588 39172 29640
rect 33692 29563 33744 29572
rect 33692 29529 33701 29563
rect 33701 29529 33735 29563
rect 33735 29529 33744 29563
rect 33692 29520 33744 29529
rect 38016 29520 38068 29572
rect 38476 29520 38528 29572
rect 26332 29452 26384 29504
rect 27620 29452 27672 29504
rect 33416 29452 33468 29504
rect 34428 29452 34480 29504
rect 38844 29520 38896 29572
rect 39856 29631 39908 29640
rect 39856 29597 39865 29631
rect 39865 29597 39899 29631
rect 39899 29597 39908 29631
rect 39856 29588 39908 29597
rect 40776 29588 40828 29640
rect 41052 29520 41104 29572
rect 38936 29452 38988 29504
rect 40500 29495 40552 29504
rect 40500 29461 40509 29495
rect 40509 29461 40543 29495
rect 40543 29461 40552 29495
rect 40500 29452 40552 29461
rect 40684 29452 40736 29504
rect 42984 29520 43036 29572
rect 42708 29495 42760 29504
rect 42708 29461 42717 29495
rect 42717 29461 42751 29495
rect 42751 29461 42760 29495
rect 42708 29452 42760 29461
rect 43076 29495 43128 29504
rect 43076 29461 43085 29495
rect 43085 29461 43119 29495
rect 43119 29461 43128 29495
rect 43076 29452 43128 29461
rect 43168 29452 43220 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4068 29248 4120 29300
rect 7748 29248 7800 29300
rect 8668 29248 8720 29300
rect 5448 29180 5500 29232
rect 5540 29223 5592 29232
rect 5540 29189 5549 29223
rect 5549 29189 5583 29223
rect 5583 29189 5592 29223
rect 5540 29180 5592 29189
rect 7196 29180 7248 29232
rect 9496 29248 9548 29300
rect 11060 29291 11112 29300
rect 11060 29257 11069 29291
rect 11069 29257 11103 29291
rect 11103 29257 11112 29291
rect 11060 29248 11112 29257
rect 15108 29248 15160 29300
rect 16028 29248 16080 29300
rect 16948 29248 17000 29300
rect 17500 29248 17552 29300
rect 17868 29248 17920 29300
rect 18052 29291 18104 29300
rect 18052 29257 18061 29291
rect 18061 29257 18095 29291
rect 18095 29257 18104 29291
rect 18052 29248 18104 29257
rect 18328 29248 18380 29300
rect 13084 29180 13136 29232
rect 13452 29180 13504 29232
rect 13728 29180 13780 29232
rect 9220 29112 9272 29164
rect 9312 29087 9364 29096
rect 9312 29053 9321 29087
rect 9321 29053 9355 29087
rect 9355 29053 9364 29087
rect 9312 29044 9364 29053
rect 17132 29155 17184 29164
rect 17132 29121 17141 29155
rect 17141 29121 17175 29155
rect 17175 29121 17184 29155
rect 17132 29112 17184 29121
rect 20536 29248 20588 29300
rect 20904 29248 20956 29300
rect 20260 29223 20312 29232
rect 20260 29189 20269 29223
rect 20269 29189 20303 29223
rect 20303 29189 20312 29223
rect 20260 29180 20312 29189
rect 18696 29112 18748 29164
rect 19340 29112 19392 29164
rect 19984 29112 20036 29164
rect 20444 29180 20496 29232
rect 16948 28976 17000 29028
rect 20812 29112 20864 29164
rect 20996 29112 21048 29164
rect 22192 29180 22244 29232
rect 23020 29223 23072 29232
rect 23020 29189 23029 29223
rect 23029 29189 23063 29223
rect 23063 29189 23072 29223
rect 23020 29180 23072 29189
rect 29000 29248 29052 29300
rect 33968 29248 34020 29300
rect 37832 29248 37884 29300
rect 26332 29112 26384 29164
rect 27436 29112 27488 29164
rect 27896 29155 27948 29164
rect 27896 29121 27905 29155
rect 27905 29121 27939 29155
rect 27939 29121 27948 29155
rect 27896 29112 27948 29121
rect 29092 29112 29144 29164
rect 27528 29044 27580 29096
rect 6184 28908 6236 28960
rect 17500 28908 17552 28960
rect 24676 28908 24728 28960
rect 26792 28908 26844 28960
rect 27620 28908 27672 28960
rect 31208 29112 31260 29164
rect 31576 29112 31628 29164
rect 33416 29155 33468 29164
rect 33416 29121 33425 29155
rect 33425 29121 33459 29155
rect 33459 29121 33468 29155
rect 33416 29112 33468 29121
rect 34612 29180 34664 29232
rect 34704 29180 34756 29232
rect 33692 29112 33744 29164
rect 38936 29180 38988 29232
rect 40592 29248 40644 29300
rect 42708 29248 42760 29300
rect 36544 29087 36596 29096
rect 36544 29053 36553 29087
rect 36553 29053 36587 29087
rect 36587 29053 36596 29087
rect 36544 29044 36596 29053
rect 37832 29087 37884 29096
rect 37832 29053 37841 29087
rect 37841 29053 37875 29087
rect 37875 29053 37884 29087
rect 37832 29044 37884 29053
rect 31024 28976 31076 29028
rect 32128 28976 32180 29028
rect 33968 28976 34020 29028
rect 34520 28976 34572 29028
rect 38200 28976 38252 29028
rect 38660 29155 38712 29164
rect 38660 29121 38669 29155
rect 38669 29121 38703 29155
rect 38703 29121 38712 29155
rect 38660 29112 38712 29121
rect 39304 29112 39356 29164
rect 42800 29180 42852 29232
rect 40868 29044 40920 29096
rect 42892 29044 42944 29096
rect 39212 28976 39264 29028
rect 31944 28908 31996 28960
rect 35992 28951 36044 28960
rect 35992 28917 36001 28951
rect 36001 28917 36035 28951
rect 36035 28917 36044 28951
rect 35992 28908 36044 28917
rect 38844 28908 38896 28960
rect 38936 28951 38988 28960
rect 38936 28917 38945 28951
rect 38945 28917 38979 28951
rect 38979 28917 38988 28951
rect 38936 28908 38988 28917
rect 39948 28908 40000 28960
rect 42432 28908 42484 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 7104 28747 7156 28756
rect 7104 28713 7113 28747
rect 7113 28713 7147 28747
rect 7147 28713 7156 28747
rect 7104 28704 7156 28713
rect 9220 28704 9272 28756
rect 10416 28704 10468 28756
rect 11520 28747 11572 28756
rect 11520 28713 11529 28747
rect 11529 28713 11563 28747
rect 11563 28713 11572 28747
rect 11520 28704 11572 28713
rect 14924 28704 14976 28756
rect 16948 28704 17000 28756
rect 19984 28704 20036 28756
rect 21180 28704 21232 28756
rect 29092 28747 29144 28756
rect 29092 28713 29101 28747
rect 29101 28713 29135 28747
rect 29135 28713 29144 28747
rect 29092 28704 29144 28713
rect 5540 28568 5592 28620
rect 6552 28568 6604 28620
rect 7196 28568 7248 28620
rect 7472 28568 7524 28620
rect 9036 28568 9088 28620
rect 20352 28636 20404 28688
rect 14924 28568 14976 28620
rect 6092 28364 6144 28416
rect 7196 28432 7248 28484
rect 7472 28364 7524 28416
rect 7748 28364 7800 28416
rect 11612 28500 11664 28552
rect 11980 28543 12032 28552
rect 11980 28509 11989 28543
rect 11989 28509 12023 28543
rect 12023 28509 12032 28543
rect 11980 28500 12032 28509
rect 12808 28543 12860 28552
rect 12808 28509 12817 28543
rect 12817 28509 12851 28543
rect 12851 28509 12860 28543
rect 12808 28500 12860 28509
rect 18052 28568 18104 28620
rect 20076 28568 20128 28620
rect 16396 28543 16448 28552
rect 16396 28509 16405 28543
rect 16405 28509 16439 28543
rect 16439 28509 16448 28543
rect 16396 28500 16448 28509
rect 16672 28500 16724 28552
rect 18512 28543 18564 28552
rect 18512 28509 18521 28543
rect 18521 28509 18555 28543
rect 18555 28509 18564 28543
rect 18512 28500 18564 28509
rect 20168 28500 20220 28552
rect 20996 28568 21048 28620
rect 22744 28611 22796 28620
rect 22744 28577 22753 28611
rect 22753 28577 22787 28611
rect 22787 28577 22796 28611
rect 22744 28568 22796 28577
rect 23848 28568 23900 28620
rect 20812 28500 20864 28552
rect 8760 28364 8812 28416
rect 9588 28364 9640 28416
rect 12072 28407 12124 28416
rect 12072 28373 12081 28407
rect 12081 28373 12115 28407
rect 12115 28373 12124 28407
rect 12072 28364 12124 28373
rect 12256 28407 12308 28416
rect 12256 28373 12265 28407
rect 12265 28373 12299 28407
rect 12299 28373 12308 28407
rect 12256 28364 12308 28373
rect 19340 28432 19392 28484
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 21732 28432 21784 28484
rect 24032 28500 24084 28552
rect 32588 28704 32640 28756
rect 33968 28747 34020 28756
rect 33968 28713 33977 28747
rect 33977 28713 34011 28747
rect 34011 28713 34020 28747
rect 33968 28704 34020 28713
rect 36912 28704 36964 28756
rect 37924 28704 37976 28756
rect 42892 28704 42944 28756
rect 31576 28636 31628 28688
rect 26240 28500 26292 28552
rect 27436 28543 27488 28552
rect 27436 28509 27445 28543
rect 27445 28509 27479 28543
rect 27479 28509 27488 28543
rect 27436 28500 27488 28509
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 17960 28407 18012 28416
rect 17960 28373 17969 28407
rect 17969 28373 18003 28407
rect 18003 28373 18012 28407
rect 17960 28364 18012 28373
rect 19984 28364 20036 28416
rect 21548 28364 21600 28416
rect 22100 28364 22152 28416
rect 22560 28407 22612 28416
rect 22560 28373 22569 28407
rect 22569 28373 22603 28407
rect 22603 28373 22612 28407
rect 22560 28364 22612 28373
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 31208 28611 31260 28620
rect 31208 28577 31217 28611
rect 31217 28577 31251 28611
rect 31251 28577 31260 28611
rect 31208 28568 31260 28577
rect 32128 28679 32180 28688
rect 32128 28645 32137 28679
rect 32137 28645 32171 28679
rect 32171 28645 32180 28679
rect 32128 28636 32180 28645
rect 32956 28611 33008 28620
rect 32956 28577 32965 28611
rect 32965 28577 32999 28611
rect 32999 28577 33008 28611
rect 32956 28568 33008 28577
rect 30564 28500 30616 28552
rect 31024 28543 31076 28552
rect 31024 28509 31033 28543
rect 31033 28509 31067 28543
rect 31067 28509 31076 28543
rect 31024 28500 31076 28509
rect 29184 28432 29236 28484
rect 23756 28407 23808 28416
rect 23756 28373 23765 28407
rect 23765 28373 23799 28407
rect 23799 28373 23808 28407
rect 23756 28364 23808 28373
rect 27620 28364 27672 28416
rect 27896 28364 27948 28416
rect 29736 28407 29788 28416
rect 29736 28373 29745 28407
rect 29745 28373 29779 28407
rect 29779 28373 29788 28407
rect 29736 28364 29788 28373
rect 30196 28432 30248 28484
rect 31392 28432 31444 28484
rect 30472 28364 30524 28416
rect 31760 28432 31812 28484
rect 32312 28543 32364 28552
rect 32312 28509 32321 28543
rect 32321 28509 32355 28543
rect 32355 28509 32364 28543
rect 32312 28500 32364 28509
rect 35992 28568 36044 28620
rect 40776 28568 40828 28620
rect 41972 28568 42024 28620
rect 33508 28432 33560 28484
rect 35348 28500 35400 28552
rect 37832 28500 37884 28552
rect 38568 28500 38620 28552
rect 39948 28500 40000 28552
rect 43076 28568 43128 28620
rect 35992 28432 36044 28484
rect 40684 28475 40736 28484
rect 40684 28441 40693 28475
rect 40693 28441 40727 28475
rect 40727 28441 40736 28475
rect 40684 28432 40736 28441
rect 41144 28432 41196 28484
rect 42432 28432 42484 28484
rect 42984 28432 43036 28484
rect 32036 28364 32088 28416
rect 32680 28407 32732 28416
rect 32680 28373 32689 28407
rect 32689 28373 32723 28407
rect 32723 28373 32732 28407
rect 32680 28364 32732 28373
rect 34336 28364 34388 28416
rect 38200 28364 38252 28416
rect 38844 28364 38896 28416
rect 42340 28364 42392 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5540 28067 5592 28076
rect 5540 28033 5549 28067
rect 5549 28033 5583 28067
rect 5583 28033 5592 28067
rect 5540 28024 5592 28033
rect 7104 28092 7156 28144
rect 5816 28067 5868 28076
rect 5816 28033 5837 28067
rect 5837 28033 5868 28067
rect 5816 28024 5868 28033
rect 6092 28067 6144 28076
rect 6092 28033 6101 28067
rect 6101 28033 6135 28067
rect 6135 28033 6144 28067
rect 6092 28024 6144 28033
rect 7840 28135 7892 28144
rect 7840 28101 7849 28135
rect 7849 28101 7883 28135
rect 7883 28101 7892 28135
rect 7840 28092 7892 28101
rect 6368 27888 6420 27940
rect 7196 27956 7248 28008
rect 7472 28024 7524 28076
rect 9036 28160 9088 28212
rect 9588 28203 9640 28212
rect 9588 28169 9597 28203
rect 9597 28169 9631 28203
rect 9631 28169 9640 28203
rect 9588 28160 9640 28169
rect 8760 28024 8812 28076
rect 9404 28135 9456 28144
rect 9404 28101 9413 28135
rect 9413 28101 9447 28135
rect 9447 28101 9456 28135
rect 9404 28092 9456 28101
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 9680 28067 9732 28076
rect 9680 28033 9689 28067
rect 9689 28033 9723 28067
rect 9723 28033 9732 28067
rect 9680 28024 9732 28033
rect 10324 28024 10376 28076
rect 12256 28160 12308 28212
rect 12440 28203 12492 28212
rect 12440 28169 12449 28203
rect 12449 28169 12483 28203
rect 12483 28169 12492 28203
rect 12440 28160 12492 28169
rect 11612 28092 11664 28144
rect 12072 28092 12124 28144
rect 16396 28160 16448 28212
rect 15660 28092 15712 28144
rect 7840 27888 7892 27940
rect 8392 27888 8444 27940
rect 12624 28067 12676 28076
rect 12624 28033 12628 28067
rect 12628 28033 12662 28067
rect 12662 28033 12676 28067
rect 12624 28024 12676 28033
rect 12532 27956 12584 28008
rect 12992 28067 13044 28076
rect 12992 28033 13000 28067
rect 13000 28033 13034 28067
rect 13034 28033 13044 28067
rect 12992 28024 13044 28033
rect 13084 28067 13136 28076
rect 13084 28033 13093 28067
rect 13093 28033 13127 28067
rect 13127 28033 13136 28067
rect 13084 28024 13136 28033
rect 13912 28024 13964 28076
rect 16948 28160 17000 28212
rect 17132 28160 17184 28212
rect 17960 28160 18012 28212
rect 20076 28160 20128 28212
rect 20812 28160 20864 28212
rect 23020 28160 23072 28212
rect 23112 28160 23164 28212
rect 23664 28160 23716 28212
rect 23756 28160 23808 28212
rect 25320 28160 25372 28212
rect 26240 28160 26292 28212
rect 13820 27956 13872 28008
rect 16672 27956 16724 28008
rect 17040 28024 17092 28076
rect 17500 28024 17552 28076
rect 29736 28160 29788 28212
rect 29920 28160 29972 28212
rect 29368 28092 29420 28144
rect 30472 28203 30524 28212
rect 30472 28169 30481 28203
rect 30481 28169 30515 28203
rect 30515 28169 30524 28203
rect 30472 28160 30524 28169
rect 31668 28160 31720 28212
rect 32312 28160 32364 28212
rect 32956 28160 33008 28212
rect 36544 28160 36596 28212
rect 30840 28135 30892 28144
rect 30840 28101 30864 28135
rect 30864 28101 30892 28135
rect 20076 28024 20128 28076
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 19156 27999 19208 28008
rect 19156 27965 19165 27999
rect 19165 27965 19199 27999
rect 19199 27965 19208 27999
rect 19156 27956 19208 27965
rect 19708 27956 19760 28008
rect 19984 27999 20036 28008
rect 19984 27965 19993 27999
rect 19993 27965 20027 27999
rect 20027 27965 20036 27999
rect 19984 27956 20036 27965
rect 20628 28067 20680 28076
rect 20628 28033 20637 28067
rect 20637 28033 20671 28067
rect 20671 28033 20680 28067
rect 20628 28024 20680 28033
rect 21548 28024 21600 28076
rect 21732 27956 21784 28008
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 27344 28067 27396 28076
rect 27344 28033 27353 28067
rect 27353 28033 27387 28067
rect 27387 28033 27396 28067
rect 27344 28024 27396 28033
rect 28080 28067 28132 28076
rect 28080 28033 28089 28067
rect 28089 28033 28123 28067
rect 28123 28033 28132 28067
rect 28080 28024 28132 28033
rect 22560 27956 22612 28008
rect 24676 27999 24728 28008
rect 5356 27863 5408 27872
rect 5356 27829 5365 27863
rect 5365 27829 5399 27863
rect 5399 27829 5408 27863
rect 5356 27820 5408 27829
rect 5908 27820 5960 27872
rect 7380 27820 7432 27872
rect 8208 27820 8260 27872
rect 8484 27863 8536 27872
rect 8484 27829 8493 27863
rect 8493 27829 8527 27863
rect 8527 27829 8536 27863
rect 8484 27820 8536 27829
rect 11152 27863 11204 27872
rect 11152 27829 11161 27863
rect 11161 27829 11195 27863
rect 11195 27829 11204 27863
rect 11152 27820 11204 27829
rect 12992 27820 13044 27872
rect 15844 27863 15896 27872
rect 15844 27829 15853 27863
rect 15853 27829 15887 27863
rect 15887 27829 15896 27863
rect 15844 27820 15896 27829
rect 17132 27863 17184 27872
rect 17132 27829 17141 27863
rect 17141 27829 17175 27863
rect 17175 27829 17184 27863
rect 17132 27820 17184 27829
rect 17224 27820 17276 27872
rect 23296 27820 23348 27872
rect 24676 27965 24685 27999
rect 24685 27965 24719 27999
rect 24719 27965 24728 27999
rect 24676 27956 24728 27965
rect 24952 27999 25004 28008
rect 24952 27965 24961 27999
rect 24961 27965 24995 27999
rect 24995 27965 25004 27999
rect 24952 27956 25004 27965
rect 28540 27956 28592 28008
rect 30564 27956 30616 28008
rect 30840 28092 30892 28101
rect 31208 28092 31260 28144
rect 31116 28067 31168 28076
rect 31116 28033 31125 28067
rect 31125 28033 31159 28067
rect 31159 28033 31168 28067
rect 31116 28024 31168 28033
rect 31944 28067 31996 28076
rect 31944 28033 31953 28067
rect 31953 28033 31987 28067
rect 31987 28033 31996 28067
rect 31944 28024 31996 28033
rect 32036 28024 32088 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 33876 28092 33928 28144
rect 33600 27999 33652 28008
rect 33600 27965 33609 27999
rect 33609 27965 33643 27999
rect 33643 27965 33652 27999
rect 33600 27956 33652 27965
rect 34336 27956 34388 28008
rect 35900 28067 35952 28076
rect 35900 28033 35909 28067
rect 35909 28033 35943 28067
rect 35943 28033 35952 28067
rect 35900 28024 35952 28033
rect 35716 27956 35768 28008
rect 36176 28024 36228 28076
rect 38200 28160 38252 28212
rect 40684 28160 40736 28212
rect 37280 28092 37332 28144
rect 38016 28092 38068 28144
rect 40500 28092 40552 28144
rect 36912 27999 36964 28008
rect 36912 27965 36921 27999
rect 36921 27965 36955 27999
rect 36955 27965 36964 27999
rect 36912 27956 36964 27965
rect 35992 27888 36044 27940
rect 37188 27888 37240 27940
rect 24584 27863 24636 27872
rect 24584 27829 24593 27863
rect 24593 27829 24627 27863
rect 24627 27829 24636 27863
rect 24584 27820 24636 27829
rect 27896 27863 27948 27872
rect 27896 27829 27905 27863
rect 27905 27829 27939 27863
rect 27939 27829 27948 27863
rect 27896 27820 27948 27829
rect 28724 27820 28776 27872
rect 30840 27820 30892 27872
rect 31116 27820 31168 27872
rect 31760 27820 31812 27872
rect 34704 27820 34756 27872
rect 37556 27999 37608 28008
rect 37556 27965 37565 27999
rect 37565 27965 37599 27999
rect 37599 27965 37608 27999
rect 37556 27956 37608 27965
rect 38016 27956 38068 28008
rect 39304 28024 39356 28076
rect 42524 28067 42576 28076
rect 42524 28033 42533 28067
rect 42533 28033 42567 28067
rect 42567 28033 42576 28067
rect 42524 28024 42576 28033
rect 38568 27888 38620 27940
rect 40224 27956 40276 28008
rect 40868 27999 40920 28008
rect 40868 27965 40877 27999
rect 40877 27965 40911 27999
rect 40911 27965 40920 27999
rect 40868 27956 40920 27965
rect 41696 27999 41748 28008
rect 41696 27965 41705 27999
rect 41705 27965 41739 27999
rect 41739 27965 41748 27999
rect 41696 27956 41748 27965
rect 38108 27820 38160 27872
rect 39212 27820 39264 27872
rect 40040 27820 40092 27872
rect 44272 27820 44324 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5356 27616 5408 27668
rect 6368 27616 6420 27668
rect 8392 27659 8444 27668
rect 8392 27625 8401 27659
rect 8401 27625 8435 27659
rect 8435 27625 8444 27659
rect 8392 27616 8444 27625
rect 11152 27616 11204 27668
rect 12808 27616 12860 27668
rect 13084 27616 13136 27668
rect 13912 27616 13964 27668
rect 15660 27616 15712 27668
rect 17040 27616 17092 27668
rect 17224 27616 17276 27668
rect 6920 27480 6972 27532
rect 12624 27480 12676 27532
rect 940 27412 992 27464
rect 6644 27455 6696 27464
rect 6644 27421 6653 27455
rect 6653 27421 6687 27455
rect 6687 27421 6696 27455
rect 6644 27412 6696 27421
rect 9312 27412 9364 27464
rect 9680 27412 9732 27464
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 15108 27523 15160 27532
rect 15108 27489 15117 27523
rect 15117 27489 15151 27523
rect 15151 27489 15160 27523
rect 15108 27480 15160 27489
rect 7380 27344 7432 27396
rect 8208 27344 8260 27396
rect 9588 27344 9640 27396
rect 12440 27344 12492 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 7104 27276 7156 27328
rect 14648 27412 14700 27464
rect 15844 27412 15896 27464
rect 15936 27412 15988 27464
rect 16948 27548 17000 27600
rect 19156 27548 19208 27600
rect 19708 27659 19760 27668
rect 19708 27625 19717 27659
rect 19717 27625 19751 27659
rect 19751 27625 19760 27659
rect 19708 27616 19760 27625
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 16672 27412 16724 27464
rect 18052 27480 18104 27532
rect 14924 27319 14976 27328
rect 14924 27285 14933 27319
rect 14933 27285 14967 27319
rect 14967 27285 14976 27319
rect 14924 27276 14976 27285
rect 16580 27276 16632 27328
rect 18052 27344 18104 27396
rect 19156 27344 19208 27396
rect 20076 27616 20128 27668
rect 22560 27616 22612 27668
rect 24400 27616 24452 27668
rect 24584 27616 24636 27668
rect 33600 27616 33652 27668
rect 35716 27616 35768 27668
rect 37648 27616 37700 27668
rect 39580 27616 39632 27668
rect 23112 27548 23164 27600
rect 21640 27455 21692 27464
rect 21640 27421 21649 27455
rect 21649 27421 21683 27455
rect 21683 27421 21692 27455
rect 21640 27412 21692 27421
rect 23480 27480 23532 27532
rect 24676 27480 24728 27532
rect 36176 27548 36228 27600
rect 37740 27548 37792 27600
rect 38384 27548 38436 27600
rect 39856 27548 39908 27600
rect 41696 27548 41748 27600
rect 26332 27480 26384 27532
rect 34336 27480 34388 27532
rect 35808 27480 35860 27532
rect 24400 27455 24452 27464
rect 24400 27421 24409 27455
rect 24409 27421 24443 27455
rect 24443 27421 24452 27455
rect 24400 27412 24452 27421
rect 24952 27412 25004 27464
rect 28356 27455 28408 27464
rect 28356 27421 28365 27455
rect 28365 27421 28399 27455
rect 28399 27421 28408 27455
rect 28356 27412 28408 27421
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 32680 27412 32732 27464
rect 33232 27412 33284 27464
rect 33784 27412 33836 27464
rect 37464 27480 37516 27532
rect 21916 27387 21968 27396
rect 21916 27353 21925 27387
rect 21925 27353 21959 27387
rect 21959 27353 21968 27387
rect 21916 27344 21968 27353
rect 23756 27319 23808 27328
rect 23756 27285 23765 27319
rect 23765 27285 23799 27319
rect 23799 27285 23808 27319
rect 23756 27276 23808 27285
rect 25320 27344 25372 27396
rect 29368 27344 29420 27396
rect 30012 27344 30064 27396
rect 32588 27344 32640 27396
rect 29460 27276 29512 27328
rect 31944 27319 31996 27328
rect 31944 27285 31953 27319
rect 31953 27285 31987 27319
rect 31987 27285 31996 27319
rect 31944 27276 31996 27285
rect 32404 27276 32456 27328
rect 32864 27276 32916 27328
rect 33876 27276 33928 27328
rect 35164 27387 35216 27396
rect 35164 27353 35173 27387
rect 35173 27353 35207 27387
rect 35207 27353 35216 27387
rect 35164 27344 35216 27353
rect 35348 27276 35400 27328
rect 35992 27276 36044 27328
rect 38660 27412 38712 27464
rect 38844 27412 38896 27464
rect 39120 27455 39172 27464
rect 39120 27421 39129 27455
rect 39129 27421 39163 27455
rect 39163 27421 39172 27455
rect 39120 27412 39172 27421
rect 37740 27344 37792 27396
rect 38476 27344 38528 27396
rect 39212 27344 39264 27396
rect 40776 27412 40828 27464
rect 41052 27480 41104 27532
rect 36728 27276 36780 27328
rect 38108 27276 38160 27328
rect 39856 27319 39908 27328
rect 39856 27285 39865 27319
rect 39865 27285 39899 27319
rect 39899 27285 39908 27319
rect 39856 27276 39908 27285
rect 41328 27344 41380 27396
rect 42800 27480 42852 27532
rect 43168 27412 43220 27464
rect 43812 27455 43864 27464
rect 43812 27421 43821 27455
rect 43821 27421 43855 27455
rect 43855 27421 43864 27455
rect 43812 27412 43864 27421
rect 41236 27276 41288 27328
rect 42800 27319 42852 27328
rect 42800 27285 42809 27319
rect 42809 27285 42843 27319
rect 42843 27285 42852 27319
rect 42800 27276 42852 27285
rect 42892 27276 42944 27328
rect 43996 27319 44048 27328
rect 43996 27285 44005 27319
rect 44005 27285 44039 27319
rect 44039 27285 44048 27319
rect 43996 27276 44048 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 10324 27115 10376 27124
rect 10324 27081 10333 27115
rect 10333 27081 10367 27115
rect 10367 27081 10376 27115
rect 10324 27072 10376 27081
rect 14924 27072 14976 27124
rect 16764 27072 16816 27124
rect 8484 27004 8536 27056
rect 6644 26868 6696 26920
rect 8576 26911 8628 26920
rect 8576 26877 8585 26911
rect 8585 26877 8619 26911
rect 8619 26877 8628 26911
rect 8576 26868 8628 26877
rect 9588 26868 9640 26920
rect 12440 27004 12492 27056
rect 17132 27072 17184 27124
rect 18512 27072 18564 27124
rect 21916 27072 21968 27124
rect 22100 27072 22152 27124
rect 24400 27072 24452 27124
rect 26240 27072 26292 27124
rect 29644 27072 29696 27124
rect 18052 26936 18104 26988
rect 19432 26936 19484 26988
rect 20628 26936 20680 26988
rect 30196 27004 30248 27056
rect 11428 26868 11480 26920
rect 13728 26868 13780 26920
rect 16580 26868 16632 26920
rect 15660 26800 15712 26852
rect 18328 26868 18380 26920
rect 20260 26868 20312 26920
rect 23480 26868 23532 26920
rect 24308 26911 24360 26920
rect 24308 26877 24317 26911
rect 24317 26877 24351 26911
rect 24351 26877 24360 26911
rect 24308 26868 24360 26877
rect 25320 26868 25372 26920
rect 28356 26868 28408 26920
rect 28724 26911 28776 26920
rect 28724 26877 28733 26911
rect 28733 26877 28767 26911
rect 28767 26877 28776 26911
rect 28724 26868 28776 26877
rect 29092 26979 29144 26988
rect 29092 26945 29101 26979
rect 29101 26945 29135 26979
rect 29135 26945 29144 26979
rect 29092 26936 29144 26945
rect 29184 26979 29236 26988
rect 29184 26945 29193 26979
rect 29193 26945 29227 26979
rect 29227 26945 29236 26979
rect 29184 26936 29236 26945
rect 29460 26979 29512 26988
rect 29460 26945 29469 26979
rect 29469 26945 29503 26979
rect 29503 26945 29512 26979
rect 29460 26936 29512 26945
rect 29552 26979 29604 26988
rect 29552 26945 29561 26979
rect 29561 26945 29595 26979
rect 29595 26945 29604 26979
rect 29552 26936 29604 26945
rect 29736 26979 29788 26988
rect 29736 26945 29745 26979
rect 29745 26945 29779 26979
rect 29779 26945 29788 26979
rect 29736 26936 29788 26945
rect 32036 27072 32088 27124
rect 32312 27115 32364 27124
rect 32312 27081 32321 27115
rect 32321 27081 32355 27115
rect 32355 27081 32364 27115
rect 32312 27072 32364 27081
rect 34520 27072 34572 27124
rect 35164 27072 35216 27124
rect 32864 26936 32916 26988
rect 34244 26936 34296 26988
rect 34428 26868 34480 26920
rect 17960 26800 18012 26852
rect 18420 26800 18472 26852
rect 25412 26800 25464 26852
rect 31300 26800 31352 26852
rect 31944 26800 31996 26852
rect 34060 26800 34112 26852
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 37464 27072 37516 27124
rect 37556 27072 37608 27124
rect 36728 26979 36780 26988
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 37740 27004 37792 27056
rect 38200 27047 38252 27056
rect 38200 27013 38209 27047
rect 38209 27013 38243 27047
rect 38243 27013 38252 27047
rect 38200 27004 38252 27013
rect 38660 27072 38712 27124
rect 42524 27072 42576 27124
rect 37372 26936 37424 26988
rect 37464 26979 37516 26988
rect 37464 26945 37473 26979
rect 37473 26945 37507 26979
rect 37507 26945 37516 26979
rect 37464 26936 37516 26945
rect 37648 26936 37700 26988
rect 37832 26979 37884 26988
rect 37832 26945 37841 26979
rect 37841 26945 37875 26979
rect 37875 26945 37884 26979
rect 37832 26936 37884 26945
rect 37924 26936 37976 26988
rect 39120 27004 39172 27056
rect 39856 27004 39908 27056
rect 39948 27004 40000 27056
rect 43260 27004 43312 27056
rect 14648 26732 14700 26784
rect 21272 26732 21324 26784
rect 29276 26732 29328 26784
rect 35900 26800 35952 26852
rect 40684 26911 40736 26920
rect 40684 26877 40693 26911
rect 40693 26877 40727 26911
rect 40727 26877 40736 26911
rect 40684 26868 40736 26877
rect 41236 26979 41288 26988
rect 41236 26945 41245 26979
rect 41245 26945 41279 26979
rect 41279 26945 41288 26979
rect 41236 26936 41288 26945
rect 44272 26979 44324 26988
rect 44272 26945 44281 26979
rect 44281 26945 44315 26979
rect 44315 26945 44324 26979
rect 44272 26936 44324 26945
rect 40960 26911 41012 26920
rect 40960 26877 40969 26911
rect 40969 26877 41003 26911
rect 41003 26877 41012 26911
rect 40960 26868 41012 26877
rect 41328 26868 41380 26920
rect 42800 26868 42852 26920
rect 43996 26911 44048 26920
rect 43996 26877 44005 26911
rect 44005 26877 44039 26911
rect 44039 26877 44048 26911
rect 43996 26868 44048 26877
rect 36176 26732 36228 26784
rect 36452 26775 36504 26784
rect 36452 26741 36461 26775
rect 36461 26741 36495 26775
rect 36495 26741 36504 26775
rect 36452 26732 36504 26741
rect 40132 26775 40184 26784
rect 40132 26741 40141 26775
rect 40141 26741 40175 26775
rect 40175 26741 40184 26775
rect 40132 26732 40184 26741
rect 42892 26800 42944 26852
rect 40960 26732 41012 26784
rect 42156 26775 42208 26784
rect 42156 26741 42165 26775
rect 42165 26741 42199 26775
rect 42199 26741 42208 26775
rect 42156 26732 42208 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1584 26528 1636 26580
rect 8576 26528 8628 26580
rect 9680 26571 9732 26580
rect 9680 26537 9689 26571
rect 9689 26537 9723 26571
rect 9723 26537 9732 26571
rect 9680 26528 9732 26537
rect 9404 26460 9456 26512
rect 5724 26392 5776 26444
rect 6276 26392 6328 26444
rect 9036 26367 9088 26376
rect 9036 26333 9045 26367
rect 9045 26333 9079 26367
rect 9079 26333 9088 26367
rect 9036 26324 9088 26333
rect 9496 26324 9548 26376
rect 13268 26528 13320 26580
rect 12532 26460 12584 26512
rect 12624 26392 12676 26444
rect 15108 26460 15160 26512
rect 17408 26460 17460 26512
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 16396 26392 16448 26444
rect 9772 26256 9824 26308
rect 10600 26256 10652 26308
rect 13912 26324 13964 26376
rect 19432 26571 19484 26580
rect 19432 26537 19441 26571
rect 19441 26537 19475 26571
rect 19475 26537 19484 26571
rect 19432 26528 19484 26537
rect 28356 26528 28408 26580
rect 31116 26528 31168 26580
rect 36452 26528 36504 26580
rect 37832 26528 37884 26580
rect 42156 26528 42208 26580
rect 43812 26528 43864 26580
rect 21640 26392 21692 26444
rect 21272 26324 21324 26376
rect 12072 26231 12124 26240
rect 12072 26197 12081 26231
rect 12081 26197 12115 26231
rect 12115 26197 12124 26231
rect 12072 26188 12124 26197
rect 13820 26188 13872 26240
rect 16580 26256 16632 26308
rect 16948 26256 17000 26308
rect 23112 26460 23164 26512
rect 23480 26435 23532 26444
rect 23480 26401 23489 26435
rect 23489 26401 23523 26435
rect 23523 26401 23532 26435
rect 23480 26392 23532 26401
rect 23572 26324 23624 26376
rect 28264 26367 28316 26376
rect 28264 26333 28273 26367
rect 28273 26333 28307 26367
rect 28307 26333 28316 26367
rect 28264 26324 28316 26333
rect 29092 26460 29144 26512
rect 29460 26460 29512 26512
rect 29736 26460 29788 26512
rect 32128 26460 32180 26512
rect 29552 26392 29604 26444
rect 14096 26231 14148 26240
rect 14096 26197 14105 26231
rect 14105 26197 14139 26231
rect 14139 26197 14148 26231
rect 14096 26188 14148 26197
rect 14556 26231 14608 26240
rect 14556 26197 14565 26231
rect 14565 26197 14599 26231
rect 14599 26197 14608 26231
rect 14556 26188 14608 26197
rect 25412 26256 25464 26308
rect 29000 26324 29052 26376
rect 30472 26435 30524 26444
rect 30472 26401 30481 26435
rect 30481 26401 30515 26435
rect 30515 26401 30524 26435
rect 30472 26392 30524 26401
rect 33876 26435 33928 26444
rect 33876 26401 33885 26435
rect 33885 26401 33919 26435
rect 33919 26401 33928 26435
rect 33876 26392 33928 26401
rect 29184 26256 29236 26308
rect 21640 26188 21692 26240
rect 23296 26188 23348 26240
rect 23572 26231 23624 26240
rect 23572 26197 23581 26231
rect 23581 26197 23615 26231
rect 23615 26197 23624 26231
rect 23572 26188 23624 26197
rect 24032 26231 24084 26240
rect 24032 26197 24041 26231
rect 24041 26197 24075 26231
rect 24075 26197 24084 26231
rect 24032 26188 24084 26197
rect 28448 26231 28500 26240
rect 28448 26197 28457 26231
rect 28457 26197 28491 26231
rect 28491 26197 28500 26231
rect 28448 26188 28500 26197
rect 29276 26188 29328 26240
rect 32036 26231 32088 26240
rect 32036 26197 32045 26231
rect 32045 26197 32079 26231
rect 32079 26197 32088 26231
rect 32036 26188 32088 26197
rect 33968 26367 34020 26376
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 40132 26435 40184 26444
rect 40132 26401 40141 26435
rect 40141 26401 40175 26435
rect 40175 26401 40184 26435
rect 40132 26392 40184 26401
rect 42340 26392 42392 26444
rect 44272 26392 44324 26444
rect 32588 26256 32640 26308
rect 33600 26299 33652 26308
rect 33600 26265 33609 26299
rect 33609 26265 33643 26299
rect 33643 26265 33652 26299
rect 33600 26256 33652 26265
rect 34060 26256 34112 26308
rect 32772 26188 32824 26240
rect 34244 26188 34296 26240
rect 35440 26324 35492 26376
rect 37096 26367 37148 26376
rect 37096 26333 37105 26367
rect 37105 26333 37139 26367
rect 37139 26333 37148 26367
rect 37096 26324 37148 26333
rect 38016 26324 38068 26376
rect 37648 26256 37700 26308
rect 38108 26256 38160 26308
rect 41144 26324 41196 26376
rect 40040 26256 40092 26308
rect 34704 26231 34756 26240
rect 34704 26197 34713 26231
rect 34713 26197 34747 26231
rect 34747 26197 34756 26231
rect 34704 26188 34756 26197
rect 35900 26188 35952 26240
rect 41604 26231 41656 26240
rect 41604 26197 41613 26231
rect 41613 26197 41647 26231
rect 41647 26197 41656 26231
rect 41604 26188 41656 26197
rect 43260 26256 43312 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5724 25984 5776 26036
rect 7840 25984 7892 26036
rect 9588 25916 9640 25968
rect 9772 25984 9824 26036
rect 12072 25984 12124 26036
rect 9036 25891 9088 25900
rect 9036 25857 9045 25891
rect 9045 25857 9079 25891
rect 9079 25857 9088 25891
rect 9036 25848 9088 25857
rect 10600 25848 10652 25900
rect 12440 25916 12492 25968
rect 13912 25984 13964 26036
rect 14556 25984 14608 26036
rect 15844 26027 15896 26036
rect 15844 25993 15853 26027
rect 15853 25993 15887 26027
rect 15887 25993 15896 26027
rect 15844 25984 15896 25993
rect 5816 25780 5868 25832
rect 6644 25780 6696 25832
rect 7932 25780 7984 25832
rect 9496 25780 9548 25832
rect 6184 25644 6236 25696
rect 9128 25687 9180 25696
rect 9128 25653 9137 25687
rect 9137 25653 9171 25687
rect 9171 25653 9180 25687
rect 9128 25644 9180 25653
rect 11060 25780 11112 25832
rect 12348 25780 12400 25832
rect 15660 25916 15712 25968
rect 16764 25916 16816 25968
rect 13728 25891 13780 25900
rect 13728 25857 13737 25891
rect 13737 25857 13771 25891
rect 13771 25857 13780 25891
rect 13728 25848 13780 25857
rect 16580 25848 16632 25900
rect 18052 25916 18104 25968
rect 13820 25780 13872 25832
rect 14372 25823 14424 25832
rect 14372 25789 14381 25823
rect 14381 25789 14415 25823
rect 14415 25789 14424 25823
rect 14372 25780 14424 25789
rect 22100 25848 22152 25900
rect 19616 25823 19668 25832
rect 19616 25789 19625 25823
rect 19625 25789 19659 25823
rect 19659 25789 19668 25823
rect 19616 25780 19668 25789
rect 17408 25712 17460 25764
rect 23572 25984 23624 26036
rect 23848 25984 23900 26036
rect 28264 25984 28316 26036
rect 25320 25916 25372 25968
rect 25412 25959 25464 25968
rect 25412 25925 25421 25959
rect 25421 25925 25455 25959
rect 25455 25925 25464 25959
rect 25412 25916 25464 25925
rect 29000 25916 29052 25968
rect 22468 25891 22520 25900
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 22468 25848 22520 25857
rect 23296 25848 23348 25900
rect 26148 25891 26200 25900
rect 26148 25857 26157 25891
rect 26157 25857 26191 25891
rect 26191 25857 26200 25891
rect 26148 25848 26200 25857
rect 23204 25823 23256 25832
rect 23204 25789 23213 25823
rect 23213 25789 23247 25823
rect 23247 25789 23256 25823
rect 23204 25780 23256 25789
rect 23664 25823 23716 25832
rect 23664 25789 23673 25823
rect 23673 25789 23707 25823
rect 23707 25789 23716 25823
rect 23664 25780 23716 25789
rect 25872 25823 25924 25832
rect 25872 25789 25881 25823
rect 25881 25789 25915 25823
rect 25915 25789 25924 25823
rect 25872 25780 25924 25789
rect 28448 25848 28500 25900
rect 29460 25984 29512 26036
rect 30472 25984 30524 26036
rect 31944 25984 31996 26036
rect 29276 25959 29328 25968
rect 29276 25925 29285 25959
rect 29285 25925 29319 25959
rect 29319 25925 29328 25959
rect 29276 25916 29328 25925
rect 29552 25959 29604 25968
rect 29552 25925 29561 25959
rect 29561 25925 29595 25959
rect 29595 25925 29604 25959
rect 29552 25916 29604 25925
rect 29736 25891 29788 25900
rect 29736 25857 29745 25891
rect 29745 25857 29779 25891
rect 29779 25857 29788 25891
rect 29736 25848 29788 25857
rect 32036 25916 32088 25968
rect 31576 25848 31628 25900
rect 32128 25891 32180 25900
rect 32128 25857 32137 25891
rect 32137 25857 32171 25891
rect 32171 25857 32180 25891
rect 32128 25848 32180 25857
rect 29184 25780 29236 25832
rect 32404 25780 32456 25832
rect 32312 25712 32364 25764
rect 33600 25984 33652 26036
rect 32864 25959 32916 25968
rect 32864 25925 32873 25959
rect 32873 25925 32907 25959
rect 32907 25925 32916 25959
rect 32864 25916 32916 25925
rect 34704 25984 34756 26036
rect 35440 25984 35492 26036
rect 35992 25984 36044 26036
rect 37096 26027 37148 26036
rect 37096 25993 37105 26027
rect 37105 25993 37139 26027
rect 37139 25993 37148 26027
rect 37096 25984 37148 25993
rect 42892 25984 42944 26036
rect 32772 25891 32824 25900
rect 32772 25857 32781 25891
rect 32781 25857 32815 25891
rect 32815 25857 32824 25891
rect 32772 25848 32824 25857
rect 34796 25848 34848 25900
rect 35900 25916 35952 25968
rect 40132 25916 40184 25968
rect 41144 25916 41196 25968
rect 35348 25891 35400 25900
rect 35348 25857 35357 25891
rect 35357 25857 35391 25891
rect 35391 25857 35400 25891
rect 35348 25848 35400 25857
rect 37372 25848 37424 25900
rect 41604 25848 41656 25900
rect 43076 25848 43128 25900
rect 32680 25780 32732 25832
rect 35716 25780 35768 25832
rect 38108 25823 38160 25832
rect 38108 25789 38117 25823
rect 38117 25789 38151 25823
rect 38151 25789 38160 25823
rect 38108 25780 38160 25789
rect 38384 25823 38436 25832
rect 38384 25789 38393 25823
rect 38393 25789 38427 25823
rect 38427 25789 38436 25823
rect 38384 25780 38436 25789
rect 42892 25780 42944 25832
rect 43168 25780 43220 25832
rect 33232 25712 33284 25764
rect 10692 25644 10744 25696
rect 13912 25687 13964 25696
rect 13912 25653 13921 25687
rect 13921 25653 13955 25687
rect 13955 25653 13964 25687
rect 13912 25644 13964 25653
rect 21088 25687 21140 25696
rect 21088 25653 21097 25687
rect 21097 25653 21131 25687
rect 21131 25653 21140 25687
rect 21088 25644 21140 25653
rect 22008 25687 22060 25696
rect 22008 25653 22017 25687
rect 22017 25653 22051 25687
rect 22051 25653 22060 25687
rect 22008 25644 22060 25653
rect 23480 25644 23532 25696
rect 26056 25644 26108 25696
rect 26332 25687 26384 25696
rect 26332 25653 26341 25687
rect 26341 25653 26375 25687
rect 26375 25653 26384 25687
rect 26332 25644 26384 25653
rect 26700 25644 26752 25696
rect 29000 25644 29052 25696
rect 29644 25644 29696 25696
rect 29736 25644 29788 25696
rect 37280 25687 37332 25696
rect 37280 25653 37289 25687
rect 37289 25653 37323 25687
rect 37323 25653 37332 25687
rect 37280 25644 37332 25653
rect 40592 25687 40644 25696
rect 40592 25653 40601 25687
rect 40601 25653 40635 25687
rect 40635 25653 40644 25687
rect 40592 25644 40644 25653
rect 41052 25644 41104 25696
rect 43444 25687 43496 25696
rect 43444 25653 43453 25687
rect 43453 25653 43487 25687
rect 43487 25653 43496 25687
rect 43444 25644 43496 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7932 25483 7984 25492
rect 7932 25449 7941 25483
rect 7941 25449 7975 25483
rect 7975 25449 7984 25483
rect 7932 25440 7984 25449
rect 9128 25440 9180 25492
rect 9588 25440 9640 25492
rect 10692 25483 10744 25492
rect 10692 25449 10713 25483
rect 10713 25449 10744 25483
rect 10692 25440 10744 25449
rect 13912 25440 13964 25492
rect 14372 25440 14424 25492
rect 18880 25483 18932 25492
rect 18880 25449 18889 25483
rect 18889 25449 18923 25483
rect 18923 25449 18932 25483
rect 18880 25440 18932 25449
rect 19616 25440 19668 25492
rect 21088 25440 21140 25492
rect 5816 25347 5868 25356
rect 5816 25313 5825 25347
rect 5825 25313 5859 25347
rect 5859 25313 5868 25347
rect 5816 25304 5868 25313
rect 6184 25304 6236 25356
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 9496 25304 9548 25356
rect 8300 25100 8352 25152
rect 9680 25304 9732 25356
rect 11060 25347 11112 25356
rect 11060 25313 11069 25347
rect 11069 25313 11103 25347
rect 11103 25313 11112 25347
rect 11060 25304 11112 25313
rect 11704 25304 11756 25356
rect 17776 25347 17828 25356
rect 17776 25313 17785 25347
rect 17785 25313 17819 25347
rect 17819 25313 17828 25347
rect 17776 25304 17828 25313
rect 12440 25236 12492 25288
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 14740 25236 14792 25288
rect 18420 25236 18472 25288
rect 11336 25211 11388 25220
rect 11336 25177 11345 25211
rect 11345 25177 11379 25211
rect 11379 25177 11388 25211
rect 11336 25168 11388 25177
rect 17132 25143 17184 25152
rect 17132 25109 17141 25143
rect 17141 25109 17175 25143
rect 17175 25109 17184 25143
rect 17132 25100 17184 25109
rect 19248 25100 19300 25152
rect 19432 25143 19484 25152
rect 19432 25109 19441 25143
rect 19441 25109 19475 25143
rect 19475 25109 19484 25143
rect 19432 25100 19484 25109
rect 20260 25236 20312 25288
rect 22468 25440 22520 25492
rect 23204 25440 23256 25492
rect 23664 25440 23716 25492
rect 21640 25304 21692 25356
rect 22008 25347 22060 25356
rect 22008 25313 22017 25347
rect 22017 25313 22051 25347
rect 22051 25313 22060 25347
rect 22008 25304 22060 25313
rect 23480 25168 23532 25220
rect 26240 25372 26292 25424
rect 26332 25372 26384 25424
rect 26700 25483 26752 25492
rect 26700 25449 26709 25483
rect 26709 25449 26743 25483
rect 26743 25449 26752 25483
rect 26700 25440 26752 25449
rect 25688 25347 25740 25356
rect 25688 25313 25697 25347
rect 25697 25313 25731 25347
rect 25731 25313 25740 25347
rect 25688 25304 25740 25313
rect 29000 25372 29052 25424
rect 24032 25236 24084 25288
rect 24216 25236 24268 25288
rect 25136 25236 25188 25288
rect 26240 25236 26292 25288
rect 23664 25100 23716 25152
rect 25872 25100 25924 25152
rect 27712 25236 27764 25288
rect 29184 25483 29236 25492
rect 29184 25449 29193 25483
rect 29193 25449 29227 25483
rect 29227 25449 29236 25483
rect 29184 25440 29236 25449
rect 29552 25440 29604 25492
rect 37280 25440 37332 25492
rect 38384 25440 38436 25492
rect 40132 25440 40184 25492
rect 40684 25440 40736 25492
rect 40960 25483 41012 25492
rect 40960 25449 40969 25483
rect 40969 25449 41003 25483
rect 41003 25449 41012 25483
rect 40960 25440 41012 25449
rect 35716 25304 35768 25356
rect 38108 25304 38160 25356
rect 43444 25304 43496 25356
rect 44272 25304 44324 25356
rect 32128 25236 32180 25288
rect 35992 25236 36044 25288
rect 39580 25279 39632 25288
rect 39580 25245 39589 25279
rect 39589 25245 39623 25279
rect 39623 25245 39632 25279
rect 39580 25236 39632 25245
rect 40224 25236 40276 25288
rect 40592 25236 40644 25288
rect 40776 25279 40828 25288
rect 40776 25245 40785 25279
rect 40785 25245 40819 25279
rect 40819 25245 40828 25279
rect 40776 25236 40828 25245
rect 41052 25279 41104 25288
rect 41052 25245 41061 25279
rect 41061 25245 41095 25279
rect 41095 25245 41104 25279
rect 41052 25236 41104 25245
rect 41236 25236 41288 25288
rect 43260 25168 43312 25220
rect 27160 25100 27212 25152
rect 31944 25143 31996 25152
rect 31944 25109 31953 25143
rect 31953 25109 31987 25143
rect 31987 25109 31996 25143
rect 31944 25100 31996 25109
rect 38016 25100 38068 25152
rect 43076 25100 43128 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 11704 24896 11756 24948
rect 15568 24939 15620 24948
rect 15568 24905 15577 24939
rect 15577 24905 15611 24939
rect 15611 24905 15620 24939
rect 15568 24896 15620 24905
rect 18420 24939 18472 24948
rect 18420 24905 18429 24939
rect 18429 24905 18463 24939
rect 18463 24905 18472 24939
rect 18420 24896 18472 24905
rect 25688 24939 25740 24948
rect 25688 24905 25697 24939
rect 25697 24905 25731 24939
rect 25731 24905 25740 24939
rect 25688 24896 25740 24905
rect 26148 24896 26200 24948
rect 15660 24828 15712 24880
rect 21640 24828 21692 24880
rect 11336 24692 11388 24744
rect 12992 24692 13044 24744
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 16580 24760 16632 24812
rect 18972 24760 19024 24812
rect 14096 24735 14148 24744
rect 14096 24701 14105 24735
rect 14105 24701 14139 24735
rect 14139 24701 14148 24735
rect 14096 24692 14148 24701
rect 16212 24735 16264 24744
rect 16212 24701 16221 24735
rect 16221 24701 16255 24735
rect 16255 24701 16264 24735
rect 16212 24692 16264 24701
rect 13820 24624 13872 24676
rect 15752 24599 15804 24608
rect 15752 24565 15761 24599
rect 15761 24565 15795 24599
rect 15795 24565 15804 24599
rect 15752 24556 15804 24565
rect 15844 24556 15896 24608
rect 16948 24735 17000 24744
rect 16948 24701 16957 24735
rect 16957 24701 16991 24735
rect 16991 24701 17000 24735
rect 16948 24692 17000 24701
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 23480 24828 23532 24880
rect 27068 24828 27120 24880
rect 27712 24939 27764 24948
rect 27712 24905 27721 24939
rect 27721 24905 27755 24939
rect 27755 24905 27764 24939
rect 27712 24896 27764 24905
rect 32128 24939 32180 24948
rect 32128 24905 32137 24939
rect 32137 24905 32171 24939
rect 32171 24905 32180 24939
rect 32128 24896 32180 24905
rect 40592 24896 40644 24948
rect 44640 24896 44692 24948
rect 26148 24803 26200 24812
rect 26148 24769 26157 24803
rect 26157 24769 26191 24803
rect 26191 24769 26200 24803
rect 26148 24760 26200 24769
rect 26240 24760 26292 24812
rect 27804 24803 27856 24812
rect 27160 24735 27212 24744
rect 27160 24701 27169 24735
rect 27169 24701 27203 24735
rect 27203 24701 27212 24735
rect 27160 24692 27212 24701
rect 23756 24624 23808 24676
rect 25872 24624 25924 24676
rect 26056 24667 26108 24676
rect 26056 24633 26065 24667
rect 26065 24633 26099 24667
rect 26099 24633 26108 24667
rect 26056 24624 26108 24633
rect 27804 24769 27813 24803
rect 27813 24769 27847 24803
rect 27847 24769 27856 24803
rect 27804 24760 27856 24769
rect 31392 24803 31444 24812
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 31576 24803 31628 24812
rect 31576 24769 31585 24803
rect 31585 24769 31619 24803
rect 31619 24769 31628 24803
rect 31576 24760 31628 24769
rect 31944 24828 31996 24880
rect 32588 24828 32640 24880
rect 32036 24760 32088 24812
rect 32312 24760 32364 24812
rect 35716 24760 35768 24812
rect 40132 24828 40184 24880
rect 37004 24760 37056 24812
rect 17684 24556 17736 24608
rect 19156 24556 19208 24608
rect 19248 24556 19300 24608
rect 22008 24556 22060 24608
rect 25136 24556 25188 24608
rect 27528 24624 27580 24676
rect 39304 24692 39356 24744
rect 27068 24599 27120 24608
rect 27068 24565 27077 24599
rect 27077 24565 27111 24599
rect 27111 24565 27120 24599
rect 27068 24556 27120 24565
rect 28540 24556 28592 24608
rect 34428 24556 34480 24608
rect 36912 24599 36964 24608
rect 36912 24565 36921 24599
rect 36921 24565 36955 24599
rect 36955 24565 36964 24599
rect 36912 24556 36964 24565
rect 39028 24599 39080 24608
rect 39028 24565 39037 24599
rect 39037 24565 39071 24599
rect 39071 24565 39080 24599
rect 39028 24556 39080 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12900 24352 12952 24404
rect 14096 24352 14148 24404
rect 15752 24352 15804 24404
rect 16948 24352 17000 24404
rect 22192 24352 22244 24404
rect 31392 24352 31444 24404
rect 13084 24284 13136 24336
rect 11060 24216 11112 24268
rect 19156 24284 19208 24336
rect 14556 24148 14608 24200
rect 16580 24216 16632 24268
rect 19984 24216 20036 24268
rect 14740 24148 14792 24200
rect 17132 24148 17184 24200
rect 22652 24259 22704 24268
rect 22652 24225 22661 24259
rect 22661 24225 22695 24259
rect 22695 24225 22704 24259
rect 22652 24216 22704 24225
rect 23572 24216 23624 24268
rect 29552 24327 29604 24336
rect 29552 24293 29561 24327
rect 29561 24293 29595 24327
rect 29595 24293 29604 24327
rect 29552 24284 29604 24293
rect 39396 24352 39448 24404
rect 42984 24352 43036 24404
rect 39028 24284 39080 24336
rect 32680 24216 32732 24268
rect 34520 24259 34572 24268
rect 34520 24225 34529 24259
rect 34529 24225 34563 24259
rect 34563 24225 34572 24259
rect 34520 24216 34572 24225
rect 11888 24123 11940 24132
rect 11888 24089 11897 24123
rect 11897 24089 11931 24123
rect 11931 24089 11940 24123
rect 11888 24080 11940 24089
rect 12440 24080 12492 24132
rect 12624 24012 12676 24064
rect 15292 24012 15344 24064
rect 17592 24123 17644 24132
rect 17592 24089 17601 24123
rect 17601 24089 17635 24123
rect 17635 24089 17644 24123
rect 17592 24080 17644 24089
rect 18052 24080 18104 24132
rect 20996 24191 21048 24200
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 22008 24148 22060 24200
rect 24584 24148 24636 24200
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 22192 24080 22244 24132
rect 29920 24148 29972 24200
rect 30012 24148 30064 24200
rect 30104 24191 30156 24200
rect 30104 24157 30113 24191
rect 30113 24157 30147 24191
rect 30147 24157 30156 24191
rect 30104 24148 30156 24157
rect 30288 24191 30340 24200
rect 30288 24157 30297 24191
rect 30297 24157 30331 24191
rect 30331 24157 30340 24191
rect 30288 24148 30340 24157
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 30840 24191 30892 24200
rect 30840 24157 30849 24191
rect 30849 24157 30883 24191
rect 30883 24157 30892 24191
rect 30840 24148 30892 24157
rect 36360 24148 36412 24200
rect 37556 24191 37608 24200
rect 37556 24157 37565 24191
rect 37565 24157 37599 24191
rect 37599 24157 37608 24191
rect 37556 24148 37608 24157
rect 40040 24216 40092 24268
rect 43536 24216 43588 24268
rect 40224 24191 40276 24200
rect 40224 24157 40233 24191
rect 40233 24157 40267 24191
rect 40267 24157 40276 24191
rect 40224 24148 40276 24157
rect 43352 24148 43404 24200
rect 33048 24123 33100 24132
rect 33048 24089 33057 24123
rect 33057 24089 33091 24123
rect 33091 24089 33100 24123
rect 33048 24080 33100 24089
rect 34796 24080 34848 24132
rect 20812 24055 20864 24064
rect 20812 24021 20821 24055
rect 20821 24021 20855 24055
rect 20855 24021 20864 24055
rect 20812 24012 20864 24021
rect 21088 24012 21140 24064
rect 22100 24012 22152 24064
rect 22284 24012 22336 24064
rect 23480 24012 23532 24064
rect 24308 24012 24360 24064
rect 29184 24012 29236 24064
rect 30104 24012 30156 24064
rect 30472 24055 30524 24064
rect 30472 24021 30481 24055
rect 30481 24021 30515 24055
rect 30515 24021 30524 24055
rect 30472 24012 30524 24021
rect 30656 24012 30708 24064
rect 34704 24055 34756 24064
rect 34704 24021 34713 24055
rect 34713 24021 34747 24055
rect 34747 24021 34756 24055
rect 34704 24012 34756 24021
rect 35808 24012 35860 24064
rect 37280 24012 37332 24064
rect 37372 24055 37424 24064
rect 37372 24021 37381 24055
rect 37381 24021 37415 24055
rect 37415 24021 37424 24055
rect 37372 24012 37424 24021
rect 39212 24012 39264 24064
rect 41144 24012 41196 24064
rect 42248 24055 42300 24064
rect 42248 24021 42257 24055
rect 42257 24021 42291 24055
rect 42291 24021 42300 24055
rect 42248 24012 42300 24021
rect 43168 24012 43220 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 11888 23808 11940 23860
rect 12900 23808 12952 23860
rect 14556 23808 14608 23860
rect 15108 23740 15160 23792
rect 17592 23808 17644 23860
rect 19248 23808 19300 23860
rect 20812 23808 20864 23860
rect 25044 23808 25096 23860
rect 29552 23808 29604 23860
rect 30472 23808 30524 23860
rect 30840 23808 30892 23860
rect 33048 23808 33100 23860
rect 20904 23740 20956 23792
rect 12992 23647 13044 23656
rect 12992 23613 13001 23647
rect 13001 23613 13035 23647
rect 13035 23613 13044 23647
rect 12992 23604 13044 23613
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 13820 23647 13872 23656
rect 13820 23613 13829 23647
rect 13829 23613 13863 23647
rect 13863 23613 13872 23647
rect 13820 23604 13872 23613
rect 19340 23604 19392 23656
rect 19432 23536 19484 23588
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 14464 23468 14516 23520
rect 15384 23511 15436 23520
rect 15384 23477 15393 23511
rect 15393 23477 15427 23511
rect 15427 23477 15436 23511
rect 15384 23468 15436 23477
rect 16212 23468 16264 23520
rect 26240 23536 26292 23588
rect 26424 23715 26476 23724
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 29736 23783 29788 23792
rect 29736 23749 29745 23783
rect 29745 23749 29779 23783
rect 29779 23749 29788 23783
rect 29736 23740 29788 23749
rect 29920 23672 29972 23724
rect 30104 23715 30156 23724
rect 30104 23681 30113 23715
rect 30113 23681 30147 23715
rect 30147 23681 30156 23715
rect 30104 23672 30156 23681
rect 30472 23715 30524 23724
rect 30472 23681 30481 23715
rect 30481 23681 30515 23715
rect 30515 23681 30524 23715
rect 30472 23672 30524 23681
rect 34704 23808 34756 23860
rect 35440 23808 35492 23860
rect 32496 23536 32548 23588
rect 34060 23715 34112 23724
rect 34060 23681 34069 23715
rect 34069 23681 34103 23715
rect 34103 23681 34112 23715
rect 34060 23672 34112 23681
rect 34152 23715 34204 23724
rect 34152 23681 34187 23715
rect 34187 23681 34204 23715
rect 34152 23672 34204 23681
rect 34612 23715 34664 23724
rect 34612 23681 34621 23715
rect 34621 23681 34655 23715
rect 34655 23681 34664 23715
rect 34612 23672 34664 23681
rect 35808 23740 35860 23792
rect 36912 23808 36964 23860
rect 39212 23808 39264 23860
rect 38660 23740 38712 23792
rect 40224 23808 40276 23860
rect 41052 23808 41104 23860
rect 42248 23808 42300 23860
rect 42800 23808 42852 23860
rect 41144 23740 41196 23792
rect 41512 23740 41564 23792
rect 37096 23647 37148 23656
rect 37096 23613 37105 23647
rect 37105 23613 37139 23647
rect 37139 23613 37148 23647
rect 37096 23604 37148 23613
rect 34704 23536 34756 23588
rect 39396 23604 39448 23656
rect 42892 23740 42944 23792
rect 42984 23672 43036 23724
rect 43352 23740 43404 23792
rect 43536 23715 43588 23724
rect 43536 23681 43545 23715
rect 43545 23681 43579 23715
rect 43579 23681 43588 23715
rect 43536 23672 43588 23681
rect 43352 23647 43404 23656
rect 43352 23613 43361 23647
rect 43361 23613 43395 23647
rect 43395 23613 43404 23647
rect 43352 23604 43404 23613
rect 21548 23468 21600 23520
rect 22284 23468 22336 23520
rect 29644 23468 29696 23520
rect 30288 23468 30340 23520
rect 35624 23468 35676 23520
rect 40132 23468 40184 23520
rect 42432 23511 42484 23520
rect 42432 23477 42441 23511
rect 42441 23477 42475 23511
rect 42475 23477 42484 23511
rect 42432 23468 42484 23477
rect 43076 23468 43128 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 13820 23264 13872 23316
rect 14372 23264 14424 23316
rect 15108 23264 15160 23316
rect 17408 23264 17460 23316
rect 17500 23264 17552 23316
rect 12992 23128 13044 23180
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 10048 22924 10100 22976
rect 10600 22967 10652 22976
rect 10600 22933 10609 22967
rect 10609 22933 10643 22967
rect 10643 22933 10652 22967
rect 10600 22924 10652 22933
rect 11796 23060 11848 23112
rect 15108 23171 15160 23180
rect 15108 23137 15117 23171
rect 15117 23137 15151 23171
rect 15151 23137 15160 23171
rect 15108 23128 15160 23137
rect 15292 23128 15344 23180
rect 15384 23060 15436 23112
rect 16396 23060 16448 23112
rect 16764 23060 16816 23112
rect 17224 23060 17276 23112
rect 14464 22992 14516 23044
rect 17500 22992 17552 23044
rect 18052 23035 18104 23044
rect 18052 23001 18061 23035
rect 18061 23001 18095 23035
rect 18095 23001 18104 23035
rect 18052 22992 18104 23001
rect 11428 22967 11480 22976
rect 11428 22933 11437 22967
rect 11437 22933 11471 22967
rect 11471 22933 11480 22967
rect 11428 22924 11480 22933
rect 14648 22924 14700 22976
rect 17040 22924 17092 22976
rect 17776 22924 17828 22976
rect 17960 22924 18012 22976
rect 20076 23128 20128 23180
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 19524 23035 19576 23044
rect 19524 23001 19533 23035
rect 19533 23001 19567 23035
rect 19567 23001 19576 23035
rect 19524 22992 19576 23001
rect 20996 23264 21048 23316
rect 21456 23264 21508 23316
rect 24216 23307 24268 23316
rect 24216 23273 24225 23307
rect 24225 23273 24259 23307
rect 24259 23273 24268 23307
rect 24216 23264 24268 23273
rect 29184 23307 29236 23316
rect 29184 23273 29193 23307
rect 29193 23273 29227 23307
rect 29227 23273 29236 23307
rect 29184 23264 29236 23273
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 21272 23128 21324 23180
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 22468 23103 22520 23112
rect 22468 23069 22477 23103
rect 22477 23069 22511 23103
rect 22511 23069 22520 23103
rect 22468 23060 22520 23069
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 30012 23264 30064 23316
rect 30288 23264 30340 23316
rect 25872 23060 25924 23112
rect 26792 23103 26844 23112
rect 26792 23069 26801 23103
rect 26801 23069 26835 23103
rect 26835 23069 26844 23103
rect 26792 23060 26844 23069
rect 28080 23103 28132 23112
rect 28080 23069 28089 23103
rect 28089 23069 28123 23103
rect 28123 23069 28132 23103
rect 28080 23060 28132 23069
rect 30472 23128 30524 23180
rect 31668 23128 31720 23180
rect 22744 23035 22796 23044
rect 22744 23001 22753 23035
rect 22753 23001 22787 23035
rect 22787 23001 22796 23035
rect 22744 22992 22796 23001
rect 24032 22992 24084 23044
rect 24124 22992 24176 23044
rect 24492 23035 24544 23044
rect 24492 23001 24501 23035
rect 24501 23001 24535 23035
rect 24535 23001 24544 23035
rect 24492 22992 24544 23001
rect 29552 23103 29604 23112
rect 29552 23069 29561 23103
rect 29561 23069 29595 23103
rect 29595 23069 29604 23103
rect 29552 23060 29604 23069
rect 29000 23035 29052 23044
rect 29000 23001 29009 23035
rect 29009 23001 29043 23035
rect 29043 23001 29052 23035
rect 29000 22992 29052 23001
rect 29828 23035 29880 23044
rect 29828 23001 29837 23035
rect 29837 23001 29871 23035
rect 29871 23001 29880 23035
rect 29828 22992 29880 23001
rect 20352 22924 20404 22976
rect 20904 22924 20956 22976
rect 21916 22924 21968 22976
rect 29092 22924 29144 22976
rect 29184 22924 29236 22976
rect 30196 22924 30248 22976
rect 37096 23264 37148 23316
rect 37372 23128 37424 23180
rect 43168 23171 43220 23180
rect 43168 23137 43177 23171
rect 43177 23137 43211 23171
rect 43211 23137 43220 23171
rect 43168 23128 43220 23137
rect 33876 23103 33928 23112
rect 33876 23069 33885 23103
rect 33885 23069 33919 23103
rect 33919 23069 33928 23103
rect 33876 23060 33928 23069
rect 34060 23103 34112 23112
rect 34060 23069 34069 23103
rect 34069 23069 34103 23103
rect 34103 23069 34112 23103
rect 34060 23060 34112 23069
rect 34520 23060 34572 23112
rect 35348 23060 35400 23112
rect 42800 23060 42852 23112
rect 43260 23060 43312 23112
rect 37280 22992 37332 23044
rect 31392 22967 31444 22976
rect 31392 22933 31401 22967
rect 31401 22933 31435 22967
rect 31435 22933 31444 22967
rect 31392 22924 31444 22933
rect 32588 22924 32640 22976
rect 32956 22924 33008 22976
rect 34244 22967 34296 22976
rect 34244 22933 34253 22967
rect 34253 22933 34287 22967
rect 34287 22933 34296 22967
rect 34244 22924 34296 22933
rect 34796 22924 34848 22976
rect 38752 22967 38804 22976
rect 38752 22933 38761 22967
rect 38761 22933 38795 22967
rect 38795 22933 38804 22967
rect 38752 22924 38804 22933
rect 42800 22924 42852 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 10048 22720 10100 22772
rect 10508 22720 10560 22772
rect 10876 22584 10928 22636
rect 11888 22627 11940 22636
rect 11888 22593 11897 22627
rect 11897 22593 11931 22627
rect 11931 22593 11940 22627
rect 11888 22584 11940 22593
rect 7748 22516 7800 22568
rect 14924 22652 14976 22704
rect 13452 22584 13504 22636
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 12992 22516 13044 22568
rect 15844 22516 15896 22568
rect 12900 22423 12952 22432
rect 12900 22389 12909 22423
rect 12909 22389 12943 22423
rect 12943 22389 12952 22423
rect 12900 22380 12952 22389
rect 17040 22652 17092 22704
rect 17408 22652 17460 22704
rect 19432 22720 19484 22772
rect 19616 22720 19668 22772
rect 20996 22720 21048 22772
rect 22744 22720 22796 22772
rect 23664 22763 23716 22772
rect 23664 22729 23673 22763
rect 23673 22729 23707 22763
rect 23707 22729 23716 22763
rect 23664 22720 23716 22729
rect 25596 22720 25648 22772
rect 26792 22720 26844 22772
rect 29000 22720 29052 22772
rect 29828 22720 29880 22772
rect 24124 22652 24176 22704
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 19708 22584 19760 22636
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 19294 22448 19346 22500
rect 19708 22448 19760 22500
rect 23388 22584 23440 22636
rect 23756 22559 23808 22568
rect 23756 22525 23765 22559
rect 23765 22525 23799 22559
rect 23799 22525 23808 22559
rect 23756 22516 23808 22525
rect 23940 22559 23992 22568
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 25688 22584 25740 22636
rect 25872 22652 25924 22704
rect 26148 22584 26200 22636
rect 28080 22625 28132 22636
rect 28080 22591 28089 22625
rect 28089 22591 28123 22625
rect 28123 22591 28132 22625
rect 28080 22584 28132 22591
rect 29276 22584 29328 22636
rect 29644 22627 29696 22636
rect 29644 22593 29653 22627
rect 29653 22593 29687 22627
rect 29687 22593 29696 22627
rect 29644 22584 29696 22593
rect 29828 22627 29880 22636
rect 29828 22593 29863 22627
rect 29863 22593 29880 22627
rect 29828 22584 29880 22593
rect 31392 22720 31444 22772
rect 31668 22720 31720 22772
rect 32588 22763 32640 22772
rect 32588 22729 32597 22763
rect 32597 22729 32631 22763
rect 32631 22729 32640 22763
rect 32588 22720 32640 22729
rect 32956 22763 33008 22772
rect 32956 22729 32965 22763
rect 32965 22729 32999 22763
rect 32999 22729 33008 22763
rect 32956 22720 33008 22729
rect 34060 22720 34112 22772
rect 34244 22720 34296 22772
rect 35348 22763 35400 22772
rect 35348 22729 35357 22763
rect 35357 22729 35391 22763
rect 35391 22729 35400 22763
rect 35348 22720 35400 22729
rect 37556 22763 37608 22772
rect 37556 22729 37565 22763
rect 37565 22729 37599 22763
rect 37599 22729 37608 22763
rect 37556 22720 37608 22729
rect 38752 22720 38804 22772
rect 30104 22516 30156 22568
rect 30380 22584 30432 22636
rect 30472 22627 30524 22636
rect 30472 22593 30481 22627
rect 30481 22593 30515 22627
rect 30515 22593 30524 22627
rect 30472 22584 30524 22593
rect 30564 22627 30616 22636
rect 30564 22593 30573 22627
rect 30573 22593 30607 22627
rect 30607 22593 30616 22627
rect 30564 22584 30616 22593
rect 30656 22627 30708 22636
rect 30656 22593 30665 22627
rect 30665 22593 30699 22627
rect 30699 22593 30708 22627
rect 30656 22584 30708 22593
rect 31760 22516 31812 22568
rect 32220 22627 32272 22636
rect 32220 22593 32229 22627
rect 32229 22593 32263 22627
rect 32263 22593 32272 22627
rect 32220 22584 32272 22593
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 25780 22448 25832 22500
rect 17592 22380 17644 22432
rect 17960 22380 18012 22432
rect 19524 22423 19576 22432
rect 19524 22389 19533 22423
rect 19533 22389 19567 22423
rect 19567 22389 19576 22423
rect 19524 22380 19576 22389
rect 20168 22380 20220 22432
rect 21824 22423 21876 22432
rect 21824 22389 21833 22423
rect 21833 22389 21867 22423
rect 21867 22389 21876 22423
rect 21824 22380 21876 22389
rect 25320 22380 25372 22432
rect 29828 22448 29880 22500
rect 30564 22448 30616 22500
rect 32404 22448 32456 22500
rect 31208 22380 31260 22432
rect 32220 22380 32272 22432
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 35808 22652 35860 22704
rect 38016 22695 38068 22704
rect 38016 22661 38025 22695
rect 38025 22661 38059 22695
rect 38059 22661 38068 22695
rect 38016 22652 38068 22661
rect 34704 22584 34756 22636
rect 37096 22627 37148 22636
rect 37096 22593 37105 22627
rect 37105 22593 37139 22627
rect 37139 22593 37148 22627
rect 37096 22584 37148 22593
rect 40132 22720 40184 22772
rect 40408 22652 40460 22704
rect 43260 22652 43312 22704
rect 36820 22559 36872 22568
rect 36820 22525 36829 22559
rect 36829 22525 36863 22559
rect 36863 22525 36872 22559
rect 36820 22516 36872 22525
rect 38108 22559 38160 22568
rect 38108 22525 38117 22559
rect 38117 22525 38151 22559
rect 38151 22525 38160 22559
rect 38108 22516 38160 22525
rect 39304 22516 39356 22568
rect 43076 22627 43128 22636
rect 43076 22593 43085 22627
rect 43085 22593 43119 22627
rect 43119 22593 43128 22627
rect 43076 22584 43128 22593
rect 43444 22584 43496 22636
rect 39856 22516 39908 22568
rect 43168 22559 43220 22568
rect 43168 22525 43177 22559
rect 43177 22525 43211 22559
rect 43211 22525 43220 22559
rect 43168 22516 43220 22525
rect 39948 22491 40000 22500
rect 39948 22457 39957 22491
rect 39957 22457 39991 22491
rect 39991 22457 40000 22491
rect 39948 22448 40000 22457
rect 40960 22448 41012 22500
rect 34520 22380 34572 22432
rect 34704 22423 34756 22432
rect 34704 22389 34713 22423
rect 34713 22389 34747 22423
rect 34747 22389 34756 22423
rect 34704 22380 34756 22389
rect 40224 22423 40276 22432
rect 40224 22389 40233 22423
rect 40233 22389 40267 22423
rect 40267 22389 40276 22423
rect 40224 22380 40276 22389
rect 41144 22380 41196 22432
rect 41696 22380 41748 22432
rect 43352 22423 43404 22432
rect 43352 22389 43361 22423
rect 43361 22389 43395 22423
rect 43395 22389 43404 22423
rect 43352 22380 43404 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 10600 22176 10652 22228
rect 11796 22176 11848 22228
rect 13452 22176 13504 22228
rect 17592 22219 17644 22228
rect 17592 22185 17601 22219
rect 17601 22185 17635 22219
rect 17635 22185 17644 22219
rect 17592 22176 17644 22185
rect 11152 22040 11204 22092
rect 12256 22040 12308 22092
rect 13544 22040 13596 22092
rect 19984 22108 20036 22160
rect 21824 22176 21876 22228
rect 25320 22219 25372 22228
rect 25320 22185 25329 22219
rect 25329 22185 25363 22219
rect 25363 22185 25372 22219
rect 25320 22176 25372 22185
rect 25964 22176 26016 22228
rect 26240 22176 26292 22228
rect 28080 22176 28132 22228
rect 28540 22176 28592 22228
rect 28908 22176 28960 22228
rect 29920 22219 29972 22228
rect 29920 22185 29929 22219
rect 29929 22185 29963 22219
rect 29963 22185 29972 22219
rect 29920 22176 29972 22185
rect 34428 22176 34480 22228
rect 25136 22108 25188 22160
rect 16672 21972 16724 22024
rect 16764 21972 16816 22024
rect 17684 21972 17736 22024
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 10876 21904 10928 21956
rect 12440 21904 12492 21956
rect 15660 21947 15712 21956
rect 15660 21913 15669 21947
rect 15669 21913 15703 21947
rect 15703 21913 15712 21947
rect 15660 21904 15712 21913
rect 17776 21904 17828 21956
rect 23020 22040 23072 22092
rect 19984 21972 20036 22024
rect 22376 21972 22428 22024
rect 23388 21972 23440 22024
rect 23848 21972 23900 22024
rect 25044 21972 25096 22024
rect 26056 22108 26108 22160
rect 28816 22108 28868 22160
rect 34612 22108 34664 22160
rect 35808 22176 35860 22228
rect 36268 22176 36320 22228
rect 40408 22219 40460 22228
rect 40408 22185 40417 22219
rect 40417 22185 40451 22219
rect 40451 22185 40460 22219
rect 40408 22176 40460 22185
rect 41236 22176 41288 22228
rect 38844 22108 38896 22160
rect 40500 22151 40552 22160
rect 40500 22117 40509 22151
rect 40509 22117 40543 22151
rect 40543 22117 40552 22151
rect 40500 22108 40552 22117
rect 29092 22040 29144 22092
rect 25688 22015 25740 22024
rect 25688 21981 25697 22015
rect 25697 21981 25731 22015
rect 25731 21981 25740 22015
rect 25688 21972 25740 21981
rect 25872 21972 25924 22024
rect 26332 22015 26384 22024
rect 26332 21981 26341 22015
rect 26341 21981 26375 22015
rect 26375 21981 26384 22015
rect 26332 21972 26384 21981
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 28954 21974 29006 22026
rect 31116 22040 31168 22092
rect 32220 22040 32272 22092
rect 34152 22040 34204 22092
rect 40132 22040 40184 22092
rect 29552 21972 29604 22024
rect 29828 22015 29880 22024
rect 29828 21981 29837 22015
rect 29837 21981 29871 22015
rect 29871 21981 29880 22015
rect 29828 21972 29880 21981
rect 30288 21972 30340 22024
rect 30748 21972 30800 22024
rect 31576 21972 31628 22024
rect 34244 21972 34296 22024
rect 34612 21972 34664 22024
rect 34704 22015 34756 22024
rect 34704 21981 34713 22015
rect 34713 21981 34747 22015
rect 34747 21981 34756 22015
rect 34704 21972 34756 21981
rect 34796 21972 34848 22024
rect 24860 21904 24912 21956
rect 27804 21904 27856 21956
rect 11060 21836 11112 21888
rect 12256 21836 12308 21888
rect 17960 21836 18012 21888
rect 19156 21836 19208 21888
rect 22192 21836 22244 21888
rect 26516 21836 26568 21888
rect 28264 21947 28316 21956
rect 28264 21913 28273 21947
rect 28273 21913 28307 21947
rect 28307 21913 28316 21947
rect 28264 21904 28316 21913
rect 28632 21904 28684 21956
rect 28816 21904 28868 21956
rect 31760 21904 31812 21956
rect 32220 21904 32272 21956
rect 32312 21904 32364 21956
rect 29184 21836 29236 21888
rect 32036 21836 32088 21888
rect 35348 21972 35400 22024
rect 35532 22015 35584 22024
rect 35532 21981 35541 22015
rect 35541 21981 35575 22015
rect 35575 21981 35584 22015
rect 35532 21972 35584 21981
rect 40224 21972 40276 22024
rect 40960 22040 41012 22092
rect 41144 22083 41196 22092
rect 41144 22049 41153 22083
rect 41153 22049 41187 22083
rect 41187 22049 41196 22083
rect 41144 22040 41196 22049
rect 41236 22083 41288 22092
rect 41236 22049 41245 22083
rect 41245 22049 41279 22083
rect 41279 22049 41288 22083
rect 41236 22040 41288 22049
rect 42892 22108 42944 22160
rect 43352 22108 43404 22160
rect 40776 22015 40828 22024
rect 40776 21981 40785 22015
rect 40785 21981 40819 22015
rect 40819 21981 40828 22015
rect 40776 21972 40828 21981
rect 36820 21836 36872 21888
rect 39488 21836 39540 21888
rect 40316 21904 40368 21956
rect 42156 22040 42208 22092
rect 41328 22015 41380 22024
rect 41328 21981 41337 22015
rect 41337 21981 41371 22015
rect 41371 21981 41380 22015
rect 41328 21972 41380 21981
rect 41512 22015 41564 22024
rect 41512 21981 41521 22015
rect 41521 21981 41555 22015
rect 41555 21981 41564 22015
rect 41512 21972 41564 21981
rect 41696 22015 41748 22024
rect 41696 21981 41705 22015
rect 41705 21981 41739 22015
rect 41739 21981 41748 22015
rect 41696 21972 41748 21981
rect 42064 21972 42116 22024
rect 42616 22015 42668 22024
rect 42616 21981 42625 22015
rect 42625 21981 42659 22015
rect 42659 21981 42668 22015
rect 42616 21972 42668 21981
rect 42800 22015 42852 22024
rect 42800 21981 42809 22015
rect 42809 21981 42843 22015
rect 42843 21981 42852 22015
rect 42800 21972 42852 21981
rect 43168 22015 43220 22024
rect 43168 21981 43177 22015
rect 43177 21981 43211 22015
rect 43211 21981 43220 22015
rect 43168 21972 43220 21981
rect 44364 22040 44416 22092
rect 43536 21972 43588 22024
rect 43628 21972 43680 22024
rect 40224 21836 40276 21888
rect 40868 21879 40920 21888
rect 40868 21845 40877 21879
rect 40877 21845 40911 21879
rect 40911 21845 40920 21879
rect 40868 21836 40920 21845
rect 41144 21836 41196 21888
rect 42340 21836 42392 21888
rect 43904 21836 43956 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 12440 21675 12492 21684
rect 12440 21641 12449 21675
rect 12449 21641 12483 21675
rect 12483 21641 12492 21675
rect 12440 21632 12492 21641
rect 15660 21632 15712 21684
rect 16672 21632 16724 21684
rect 17868 21632 17920 21684
rect 10508 21496 10560 21548
rect 12900 21496 12952 21548
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 13544 21564 13596 21616
rect 14372 21564 14424 21616
rect 19984 21632 20036 21684
rect 22008 21632 22060 21684
rect 22284 21675 22336 21684
rect 22284 21641 22293 21675
rect 22293 21641 22327 21675
rect 22327 21641 22336 21675
rect 22284 21632 22336 21641
rect 24032 21632 24084 21684
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 20352 21564 20404 21616
rect 21180 21564 21232 21616
rect 21640 21607 21692 21616
rect 21640 21573 21649 21607
rect 21649 21573 21683 21607
rect 21683 21573 21692 21607
rect 21640 21564 21692 21573
rect 15108 21428 15160 21480
rect 6920 21292 6972 21344
rect 7748 21292 7800 21344
rect 19892 21471 19944 21480
rect 19892 21437 19901 21471
rect 19901 21437 19935 21471
rect 19935 21437 19944 21471
rect 19892 21428 19944 21437
rect 22744 21496 22796 21548
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 23572 21496 23624 21548
rect 26240 21564 26292 21616
rect 28264 21632 28316 21684
rect 28632 21632 28684 21684
rect 36360 21632 36412 21684
rect 33232 21564 33284 21616
rect 33784 21607 33836 21616
rect 33784 21573 33793 21607
rect 33793 21573 33827 21607
rect 33827 21573 33836 21607
rect 33784 21564 33836 21573
rect 21272 21428 21324 21480
rect 23940 21428 23992 21480
rect 28080 21496 28132 21548
rect 28356 21496 28408 21548
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 28908 21539 28960 21548
rect 28908 21505 28917 21539
rect 28917 21505 28951 21539
rect 28951 21505 28960 21539
rect 28908 21496 28960 21505
rect 31944 21539 31996 21548
rect 31944 21505 31953 21539
rect 31953 21505 31987 21539
rect 31987 21505 31996 21539
rect 31944 21496 31996 21505
rect 33968 21496 34020 21548
rect 34520 21564 34572 21616
rect 40040 21632 40092 21684
rect 40868 21632 40920 21684
rect 41144 21632 41196 21684
rect 41512 21632 41564 21684
rect 42984 21632 43036 21684
rect 43536 21632 43588 21684
rect 38752 21539 38804 21548
rect 38752 21505 38761 21539
rect 38761 21505 38795 21539
rect 38795 21505 38804 21539
rect 38752 21496 38804 21505
rect 39488 21496 39540 21548
rect 39580 21496 39632 21548
rect 38844 21471 38896 21480
rect 38844 21437 38853 21471
rect 38853 21437 38887 21471
rect 38887 21437 38896 21471
rect 38844 21428 38896 21437
rect 34060 21403 34112 21412
rect 34060 21369 34069 21403
rect 34069 21369 34103 21403
rect 34103 21369 34112 21403
rect 39304 21428 39356 21480
rect 39948 21607 40000 21616
rect 39948 21573 39957 21607
rect 39957 21573 39991 21607
rect 39991 21573 40000 21607
rect 39948 21564 40000 21573
rect 40132 21539 40184 21548
rect 40132 21505 40141 21539
rect 40141 21505 40175 21539
rect 40175 21505 40184 21539
rect 40132 21496 40184 21505
rect 40224 21539 40276 21548
rect 40224 21505 40233 21539
rect 40233 21505 40267 21539
rect 40267 21505 40276 21539
rect 40224 21496 40276 21505
rect 40592 21539 40644 21548
rect 40592 21505 40601 21539
rect 40601 21505 40635 21539
rect 40635 21505 40644 21539
rect 40592 21496 40644 21505
rect 39948 21428 40000 21480
rect 34060 21360 34112 21369
rect 39856 21360 39908 21412
rect 42432 21496 42484 21548
rect 42524 21496 42576 21548
rect 42892 21539 42944 21548
rect 42892 21505 42901 21539
rect 42901 21505 42935 21539
rect 42935 21505 42944 21539
rect 42892 21496 42944 21505
rect 43076 21496 43128 21548
rect 43444 21496 43496 21548
rect 43628 21496 43680 21548
rect 41420 21428 41472 21480
rect 41236 21360 41288 21412
rect 41696 21428 41748 21480
rect 42064 21471 42116 21480
rect 42064 21437 42073 21471
rect 42073 21437 42107 21471
rect 42107 21437 42116 21471
rect 42064 21428 42116 21437
rect 41972 21403 42024 21412
rect 41972 21369 41981 21403
rect 41981 21369 42015 21403
rect 42015 21369 42024 21403
rect 41972 21360 42024 21369
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 25872 21292 25924 21344
rect 25964 21335 26016 21344
rect 25964 21301 25973 21335
rect 25973 21301 26007 21335
rect 26007 21301 26016 21335
rect 25964 21292 26016 21301
rect 28632 21292 28684 21344
rect 29184 21292 29236 21344
rect 29552 21292 29604 21344
rect 30840 21292 30892 21344
rect 34336 21335 34388 21344
rect 34336 21301 34345 21335
rect 34345 21301 34379 21335
rect 34379 21301 34388 21335
rect 34336 21292 34388 21301
rect 34428 21292 34480 21344
rect 39120 21335 39172 21344
rect 39120 21301 39129 21335
rect 39129 21301 39163 21335
rect 39163 21301 39172 21335
rect 39120 21292 39172 21301
rect 39396 21292 39448 21344
rect 40224 21292 40276 21344
rect 40408 21335 40460 21344
rect 40408 21301 40417 21335
rect 40417 21301 40451 21335
rect 40451 21301 40460 21335
rect 40408 21292 40460 21301
rect 41328 21292 41380 21344
rect 43168 21335 43220 21344
rect 43168 21301 43177 21335
rect 43177 21301 43211 21335
rect 43211 21301 43220 21335
rect 43168 21292 43220 21301
rect 43260 21335 43312 21344
rect 43260 21301 43269 21335
rect 43269 21301 43303 21335
rect 43303 21301 43312 21335
rect 43260 21292 43312 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13084 21088 13136 21140
rect 16028 21088 16080 21140
rect 19892 21088 19944 21140
rect 24584 21088 24636 21140
rect 25964 21088 26016 21140
rect 28724 21088 28776 21140
rect 29184 21131 29236 21140
rect 29184 21097 29193 21131
rect 29193 21097 29227 21131
rect 29227 21097 29236 21131
rect 29184 21088 29236 21097
rect 33968 21088 34020 21140
rect 34152 21088 34204 21140
rect 34336 21088 34388 21140
rect 39580 21088 39632 21140
rect 40040 21088 40092 21140
rect 41328 21131 41380 21140
rect 41328 21097 41337 21131
rect 41337 21097 41371 21131
rect 41371 21097 41380 21131
rect 41328 21088 41380 21097
rect 8300 20952 8352 21004
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 17316 20995 17368 21004
rect 17316 20961 17325 20995
rect 17325 20961 17359 20995
rect 17359 20961 17368 20995
rect 17316 20952 17368 20961
rect 13912 20884 13964 20936
rect 15108 20884 15160 20936
rect 17960 20884 18012 20936
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 22468 20995 22520 21004
rect 22468 20961 22477 20995
rect 22477 20961 22511 20995
rect 22511 20961 22520 20995
rect 22468 20952 22520 20961
rect 23112 20952 23164 21004
rect 28908 21020 28960 21072
rect 28172 20952 28224 21004
rect 30012 21020 30064 21072
rect 21640 20884 21692 20936
rect 25044 20884 25096 20936
rect 26056 20884 26108 20936
rect 24032 20816 24084 20868
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 14556 20791 14608 20800
rect 14556 20757 14565 20791
rect 14565 20757 14599 20791
rect 14599 20757 14608 20791
rect 14556 20748 14608 20757
rect 17132 20791 17184 20800
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 18328 20791 18380 20800
rect 18328 20757 18337 20791
rect 18337 20757 18371 20791
rect 18371 20757 18380 20791
rect 18328 20748 18380 20757
rect 20720 20748 20772 20800
rect 21180 20791 21232 20800
rect 21180 20757 21189 20791
rect 21189 20757 21223 20791
rect 21223 20757 21232 20791
rect 21180 20748 21232 20757
rect 25964 20748 26016 20800
rect 26976 20748 27028 20800
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 28632 20927 28684 20936
rect 28632 20893 28641 20927
rect 28641 20893 28675 20927
rect 28675 20893 28684 20927
rect 28632 20884 28684 20893
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 29828 20952 29880 21004
rect 30748 20952 30800 21004
rect 30380 20927 30432 20936
rect 30380 20893 30389 20927
rect 30389 20893 30423 20927
rect 30423 20893 30432 20927
rect 30380 20884 30432 20893
rect 31024 20884 31076 20936
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 31208 20884 31260 20936
rect 31852 20884 31904 20936
rect 29552 20859 29604 20868
rect 29552 20825 29561 20859
rect 29561 20825 29595 20859
rect 29595 20825 29604 20859
rect 29552 20816 29604 20825
rect 32220 20884 32272 20936
rect 29828 20748 29880 20800
rect 30564 20748 30616 20800
rect 32956 20791 33008 20800
rect 32956 20757 32965 20791
rect 32965 20757 32999 20791
rect 32999 20757 33008 20791
rect 32956 20748 33008 20757
rect 39028 21020 39080 21072
rect 33232 20816 33284 20868
rect 33508 20859 33560 20868
rect 33508 20825 33517 20859
rect 33517 20825 33551 20859
rect 33551 20825 33560 20859
rect 33508 20816 33560 20825
rect 34612 20884 34664 20936
rect 35624 20952 35676 21004
rect 38568 20952 38620 21004
rect 36636 20927 36688 20936
rect 36636 20893 36645 20927
rect 36645 20893 36679 20927
rect 36679 20893 36688 20927
rect 36636 20884 36688 20893
rect 33968 20816 34020 20868
rect 33692 20748 33744 20800
rect 34428 20816 34480 20868
rect 34520 20748 34572 20800
rect 34704 20791 34756 20800
rect 34704 20757 34713 20791
rect 34713 20757 34747 20791
rect 34747 20757 34756 20791
rect 34704 20748 34756 20757
rect 34796 20748 34848 20800
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 39396 20995 39448 21004
rect 39396 20961 39405 20995
rect 39405 20961 39439 20995
rect 39439 20961 39448 20995
rect 39396 20952 39448 20961
rect 40776 21020 40828 21072
rect 41420 21020 41472 21072
rect 42156 21088 42208 21140
rect 43168 21131 43220 21140
rect 43168 21097 43177 21131
rect 43177 21097 43211 21131
rect 43211 21097 43220 21131
rect 43168 21088 43220 21097
rect 43260 21088 43312 21140
rect 38292 20884 38344 20893
rect 38844 20884 38896 20936
rect 38936 20927 38988 20936
rect 38936 20893 38945 20927
rect 38945 20893 38979 20927
rect 38979 20893 38988 20927
rect 38936 20884 38988 20893
rect 39396 20748 39448 20800
rect 39948 20884 40000 20936
rect 40316 20884 40368 20936
rect 42616 21020 42668 21072
rect 42892 20952 42944 21004
rect 41236 20816 41288 20868
rect 41696 20927 41748 20936
rect 41696 20893 41705 20927
rect 41705 20893 41739 20927
rect 41739 20893 41748 20927
rect 41696 20884 41748 20893
rect 42156 20927 42208 20936
rect 42156 20893 42165 20927
rect 42165 20893 42199 20927
rect 42199 20893 42208 20927
rect 42156 20884 42208 20893
rect 42524 20927 42576 20936
rect 42524 20893 42533 20927
rect 42533 20893 42567 20927
rect 42567 20893 42576 20927
rect 42524 20884 42576 20893
rect 42616 20927 42668 20936
rect 42616 20893 42625 20927
rect 42625 20893 42659 20927
rect 42659 20893 42668 20927
rect 42616 20884 42668 20893
rect 43076 20884 43128 20936
rect 43352 20927 43404 20936
rect 43352 20893 43361 20927
rect 43361 20893 43395 20927
rect 43395 20893 43404 20927
rect 43352 20884 43404 20893
rect 43628 20927 43680 20936
rect 43628 20893 43637 20927
rect 43637 20893 43671 20927
rect 43671 20893 43680 20927
rect 43628 20884 43680 20893
rect 40224 20748 40276 20800
rect 42248 20748 42300 20800
rect 42892 20748 42944 20800
rect 42984 20748 43036 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 11980 20544 12032 20596
rect 14556 20544 14608 20596
rect 8116 20340 8168 20392
rect 14648 20476 14700 20528
rect 12348 20408 12400 20460
rect 13728 20408 13780 20460
rect 16212 20544 16264 20596
rect 19708 20587 19760 20596
rect 19708 20553 19717 20587
rect 19717 20553 19751 20587
rect 19751 20553 19760 20587
rect 19708 20544 19760 20553
rect 20628 20544 20680 20596
rect 23296 20544 23348 20596
rect 23480 20587 23532 20596
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 28540 20544 28592 20596
rect 29828 20544 29880 20596
rect 18328 20476 18380 20528
rect 20352 20476 20404 20528
rect 22560 20476 22612 20528
rect 12072 20383 12124 20392
rect 12072 20349 12081 20383
rect 12081 20349 12115 20383
rect 12115 20349 12124 20383
rect 12072 20340 12124 20349
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 14740 20340 14792 20392
rect 16028 20383 16080 20392
rect 16028 20349 16037 20383
rect 16037 20349 16071 20383
rect 16071 20349 16080 20383
rect 16028 20340 16080 20349
rect 17868 20408 17920 20460
rect 20996 20451 21048 20460
rect 20996 20417 21005 20451
rect 21005 20417 21039 20451
rect 21039 20417 21048 20451
rect 20996 20408 21048 20417
rect 28172 20408 28224 20460
rect 28356 20408 28408 20460
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29552 20451 29604 20460
rect 29552 20417 29561 20451
rect 29561 20417 29595 20451
rect 29595 20417 29604 20451
rect 29552 20408 29604 20417
rect 30104 20451 30156 20460
rect 30104 20417 30113 20451
rect 30113 20417 30147 20451
rect 30147 20417 30156 20451
rect 30104 20408 30156 20417
rect 30196 20451 30248 20460
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30196 20408 30248 20417
rect 30288 20408 30340 20460
rect 33968 20544 34020 20596
rect 34612 20544 34664 20596
rect 36636 20587 36688 20596
rect 36636 20553 36645 20587
rect 36645 20553 36679 20587
rect 36679 20553 36688 20587
rect 36636 20544 36688 20553
rect 31300 20451 31352 20460
rect 31300 20417 31309 20451
rect 31309 20417 31343 20451
rect 31343 20417 31352 20451
rect 31300 20408 31352 20417
rect 19248 20340 19300 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 23572 20340 23624 20349
rect 23940 20340 23992 20392
rect 29092 20340 29144 20392
rect 11244 20272 11296 20324
rect 10600 20204 10652 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 24860 20272 24912 20324
rect 28908 20272 28960 20324
rect 20812 20247 20864 20256
rect 20812 20213 20821 20247
rect 20821 20213 20855 20247
rect 20855 20213 20864 20247
rect 20812 20204 20864 20213
rect 26148 20204 26200 20256
rect 29828 20272 29880 20324
rect 29920 20272 29972 20324
rect 32956 20340 33008 20392
rect 33416 20272 33468 20324
rect 33692 20451 33744 20460
rect 33692 20417 33701 20451
rect 33701 20417 33735 20451
rect 33735 20417 33744 20451
rect 33692 20408 33744 20417
rect 34520 20408 34572 20460
rect 34704 20476 34756 20528
rect 36268 20408 36320 20460
rect 37648 20544 37700 20596
rect 39856 20544 39908 20596
rect 40316 20544 40368 20596
rect 42156 20544 42208 20596
rect 42524 20544 42576 20596
rect 39764 20476 39816 20528
rect 37464 20408 37516 20460
rect 38292 20408 38344 20460
rect 39028 20451 39080 20460
rect 39028 20417 39037 20451
rect 39037 20417 39071 20451
rect 39071 20417 39080 20451
rect 39028 20408 39080 20417
rect 39120 20408 39172 20460
rect 42248 20476 42300 20528
rect 43444 20476 43496 20528
rect 34060 20272 34112 20324
rect 34796 20272 34848 20324
rect 29736 20204 29788 20256
rect 33600 20204 33652 20256
rect 34336 20247 34388 20256
rect 34336 20213 34345 20247
rect 34345 20213 34379 20247
rect 34379 20213 34388 20247
rect 34336 20204 34388 20213
rect 34520 20247 34572 20256
rect 34520 20213 34529 20247
rect 34529 20213 34563 20247
rect 34563 20213 34572 20247
rect 34520 20204 34572 20213
rect 37556 20340 37608 20392
rect 36544 20272 36596 20324
rect 35900 20204 35952 20256
rect 38844 20247 38896 20256
rect 38844 20213 38853 20247
rect 38853 20213 38887 20247
rect 38887 20213 38896 20247
rect 38844 20204 38896 20213
rect 42800 20247 42852 20256
rect 42800 20213 42809 20247
rect 42809 20213 42843 20247
rect 42843 20213 42852 20247
rect 42800 20204 42852 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10600 20000 10652 20052
rect 11980 20000 12032 20052
rect 13728 20000 13780 20052
rect 14280 20000 14332 20052
rect 15476 20043 15528 20052
rect 15476 20009 15506 20043
rect 15506 20009 15528 20043
rect 15476 20000 15528 20009
rect 15844 20000 15896 20052
rect 17316 20000 17368 20052
rect 7196 19932 7248 19984
rect 8116 19932 8168 19984
rect 9496 19864 9548 19916
rect 11152 19864 11204 19916
rect 13084 19864 13136 19916
rect 15016 19864 15068 19916
rect 15200 19907 15252 19916
rect 15200 19873 15209 19907
rect 15209 19873 15243 19907
rect 15243 19873 15252 19907
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 18512 20000 18564 20052
rect 20536 20000 20588 20052
rect 22652 20000 22704 20052
rect 28356 20000 28408 20052
rect 28632 20000 28684 20052
rect 28908 20000 28960 20052
rect 15200 19864 15252 19873
rect 7012 19796 7064 19848
rect 14464 19796 14516 19848
rect 7012 19660 7064 19712
rect 10968 19728 11020 19780
rect 17316 19796 17368 19848
rect 18604 19839 18656 19848
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 19708 19796 19760 19848
rect 7840 19660 7892 19712
rect 11152 19660 11204 19712
rect 15752 19728 15804 19780
rect 16764 19728 16816 19780
rect 14556 19660 14608 19712
rect 16212 19660 16264 19712
rect 17408 19771 17460 19780
rect 17408 19737 17417 19771
rect 17417 19737 17451 19771
rect 17451 19737 17460 19771
rect 17408 19728 17460 19737
rect 18512 19728 18564 19780
rect 19248 19728 19300 19780
rect 21916 19932 21968 19984
rect 25780 19932 25832 19984
rect 22468 19864 22520 19916
rect 26332 19932 26384 19984
rect 24860 19796 24912 19848
rect 25688 19796 25740 19848
rect 26056 19907 26108 19916
rect 26056 19873 26065 19907
rect 26065 19873 26099 19907
rect 26099 19873 26108 19907
rect 26056 19864 26108 19873
rect 29368 19932 29420 19984
rect 28264 19907 28316 19916
rect 28264 19873 28273 19907
rect 28273 19873 28307 19907
rect 28307 19873 28316 19907
rect 28264 19864 28316 19873
rect 30012 20043 30064 20052
rect 30012 20009 30021 20043
rect 30021 20009 30055 20043
rect 30055 20009 30064 20043
rect 30012 20000 30064 20009
rect 30104 20000 30156 20052
rect 31024 20043 31076 20052
rect 31024 20009 31033 20043
rect 31033 20009 31067 20043
rect 31067 20009 31076 20043
rect 31024 20000 31076 20009
rect 33416 20000 33468 20052
rect 29920 19975 29972 19984
rect 29920 19941 29929 19975
rect 29929 19941 29963 19975
rect 29963 19941 29972 19975
rect 29920 19932 29972 19941
rect 25872 19796 25924 19848
rect 29000 19796 29052 19848
rect 29736 19864 29788 19916
rect 20812 19771 20864 19780
rect 20812 19737 20821 19771
rect 20821 19737 20855 19771
rect 20855 19737 20864 19771
rect 20812 19728 20864 19737
rect 22376 19728 22428 19780
rect 26148 19728 26200 19780
rect 28816 19728 28868 19780
rect 31576 19864 31628 19916
rect 32312 19907 32364 19916
rect 32312 19873 32321 19907
rect 32321 19873 32355 19907
rect 32355 19873 32364 19907
rect 32312 19864 32364 19873
rect 31760 19796 31812 19848
rect 30012 19728 30064 19780
rect 33600 19839 33652 19848
rect 33600 19805 33609 19839
rect 33609 19805 33643 19839
rect 33643 19805 33652 19839
rect 33600 19796 33652 19805
rect 36636 20000 36688 20052
rect 38292 20000 38344 20052
rect 38936 20000 38988 20052
rect 39396 19975 39448 19984
rect 39396 19941 39405 19975
rect 39405 19941 39439 19975
rect 39439 19941 39448 19975
rect 39396 19932 39448 19941
rect 36544 19864 36596 19916
rect 38568 19907 38620 19916
rect 38568 19873 38577 19907
rect 38577 19873 38611 19907
rect 38611 19873 38620 19907
rect 38568 19864 38620 19873
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 20444 19660 20496 19712
rect 20628 19660 20680 19712
rect 21180 19660 21232 19712
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 27804 19660 27856 19712
rect 29000 19660 29052 19712
rect 29184 19660 29236 19712
rect 35992 19796 36044 19848
rect 37464 19728 37516 19780
rect 40132 19839 40184 19848
rect 40132 19805 40141 19839
rect 40141 19805 40175 19839
rect 40175 19805 40184 19839
rect 40132 19796 40184 19805
rect 39764 19728 39816 19780
rect 42984 19796 43036 19848
rect 43444 19728 43496 19780
rect 33784 19660 33836 19712
rect 33876 19703 33928 19712
rect 33876 19669 33885 19703
rect 33885 19669 33919 19703
rect 33919 19669 33928 19703
rect 33876 19660 33928 19669
rect 34428 19660 34480 19712
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 39488 19703 39540 19712
rect 39488 19669 39497 19703
rect 39497 19669 39531 19703
rect 39531 19669 39540 19703
rect 39488 19660 39540 19669
rect 42524 19703 42576 19712
rect 42524 19669 42533 19703
rect 42533 19669 42567 19703
rect 42567 19669 42576 19703
rect 42524 19660 42576 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 6920 19456 6972 19508
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 14740 19456 14792 19508
rect 15200 19456 15252 19508
rect 16028 19456 16080 19508
rect 16764 19456 16816 19508
rect 7012 19388 7064 19440
rect 11612 19388 11664 19440
rect 12072 19388 12124 19440
rect 13452 19431 13504 19440
rect 13452 19397 13461 19431
rect 13461 19397 13495 19431
rect 13495 19397 13504 19431
rect 13452 19388 13504 19397
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 8484 19320 8536 19372
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 11060 19320 11112 19372
rect 14648 19320 14700 19372
rect 18420 19388 18472 19440
rect 17316 19320 17368 19372
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 20996 19456 21048 19508
rect 21180 19456 21232 19508
rect 22468 19456 22520 19508
rect 23756 19456 23808 19508
rect 26148 19456 26200 19508
rect 28264 19456 28316 19508
rect 19432 19388 19484 19440
rect 19892 19431 19944 19440
rect 19892 19397 19901 19431
rect 19901 19397 19935 19431
rect 19935 19397 19944 19431
rect 19892 19388 19944 19397
rect 22376 19388 22428 19440
rect 25780 19388 25832 19440
rect 21364 19363 21416 19372
rect 21364 19329 21373 19363
rect 21373 19329 21407 19363
rect 21407 19329 21416 19363
rect 21364 19320 21416 19329
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22468 19320 22520 19372
rect 25504 19320 25556 19372
rect 27804 19388 27856 19440
rect 26240 19320 26292 19372
rect 28816 19499 28868 19508
rect 28816 19465 28825 19499
rect 28825 19465 28859 19499
rect 28859 19465 28868 19499
rect 28816 19456 28868 19465
rect 29092 19456 29144 19508
rect 29920 19499 29972 19508
rect 29920 19465 29929 19499
rect 29929 19465 29963 19499
rect 29963 19465 29972 19499
rect 29920 19456 29972 19465
rect 7932 19295 7984 19304
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 10140 19252 10192 19304
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 21456 19184 21508 19236
rect 27712 19252 27764 19304
rect 30380 19320 30432 19372
rect 32036 19456 32088 19508
rect 33876 19456 33928 19508
rect 34520 19456 34572 19508
rect 39488 19456 39540 19508
rect 39580 19456 39632 19508
rect 42524 19456 42576 19508
rect 31576 19320 31628 19372
rect 31668 19363 31720 19372
rect 31668 19329 31677 19363
rect 31677 19329 31711 19363
rect 31711 19329 31720 19363
rect 31668 19320 31720 19329
rect 31760 19320 31812 19372
rect 32588 19320 32640 19372
rect 33784 19320 33836 19372
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 34428 19320 34480 19329
rect 42800 19456 42852 19508
rect 42708 19363 42760 19372
rect 42708 19329 42717 19363
rect 42717 19329 42751 19363
rect 42751 19329 42760 19363
rect 42708 19320 42760 19329
rect 42892 19320 42944 19372
rect 42984 19320 43036 19372
rect 43444 19320 43496 19372
rect 43628 19363 43680 19372
rect 43628 19329 43637 19363
rect 43637 19329 43671 19363
rect 43671 19329 43680 19363
rect 43628 19320 43680 19329
rect 7380 19159 7432 19168
rect 7380 19125 7389 19159
rect 7389 19125 7423 19159
rect 7423 19125 7432 19159
rect 7380 19116 7432 19125
rect 17132 19116 17184 19168
rect 17868 19116 17920 19168
rect 26148 19159 26200 19168
rect 26148 19125 26157 19159
rect 26157 19125 26191 19159
rect 26191 19125 26200 19159
rect 26148 19116 26200 19125
rect 31852 19184 31904 19236
rect 31116 19159 31168 19168
rect 31116 19125 31125 19159
rect 31125 19125 31159 19159
rect 31159 19125 31168 19159
rect 31116 19116 31168 19125
rect 33692 19159 33744 19168
rect 33692 19125 33701 19159
rect 33701 19125 33735 19159
rect 33735 19125 33744 19159
rect 33692 19116 33744 19125
rect 35808 19116 35860 19168
rect 37832 19116 37884 19168
rect 38200 19116 38252 19168
rect 42984 19159 43036 19168
rect 42984 19125 42993 19159
rect 42993 19125 43027 19159
rect 43027 19125 43036 19159
rect 42984 19116 43036 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7932 18912 7984 18964
rect 9496 18912 9548 18964
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 15016 18912 15068 18964
rect 18604 18912 18656 18964
rect 22192 18912 22244 18964
rect 23756 18955 23808 18964
rect 23756 18921 23765 18955
rect 23765 18921 23799 18955
rect 23799 18921 23808 18955
rect 23756 18912 23808 18921
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 26332 18955 26384 18964
rect 26332 18921 26341 18955
rect 26341 18921 26375 18955
rect 26375 18921 26384 18955
rect 26332 18912 26384 18921
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 8300 18776 8352 18828
rect 10784 18844 10836 18896
rect 11612 18776 11664 18828
rect 14648 18776 14700 18828
rect 940 18708 992 18760
rect 4620 18708 4672 18760
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 9220 18708 9272 18760
rect 10692 18708 10744 18760
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 4712 18572 4764 18624
rect 11888 18640 11940 18692
rect 7656 18572 7708 18624
rect 7840 18572 7892 18624
rect 11244 18572 11296 18624
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12440 18572 12492 18581
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 15752 18776 15804 18828
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 32588 18955 32640 18964
rect 32588 18921 32597 18955
rect 32597 18921 32631 18955
rect 32631 18921 32640 18955
rect 32588 18912 32640 18921
rect 33692 18912 33744 18964
rect 42340 18912 42392 18964
rect 42892 18912 42944 18964
rect 43352 18955 43404 18964
rect 43352 18921 43361 18955
rect 43361 18921 43395 18955
rect 43395 18921 43404 18955
rect 43352 18912 43404 18921
rect 32864 18844 32916 18896
rect 16028 18708 16080 18760
rect 19340 18776 19392 18828
rect 21456 18776 21508 18828
rect 23480 18776 23532 18828
rect 21916 18708 21968 18760
rect 23112 18708 23164 18760
rect 25780 18708 25832 18760
rect 25872 18708 25924 18760
rect 30840 18819 30892 18828
rect 30840 18785 30849 18819
rect 30849 18785 30883 18819
rect 30883 18785 30892 18819
rect 30840 18776 30892 18785
rect 31116 18819 31168 18828
rect 31116 18785 31125 18819
rect 31125 18785 31159 18819
rect 31159 18785 31168 18819
rect 31116 18776 31168 18785
rect 35716 18844 35768 18896
rect 38200 18844 38252 18896
rect 38936 18844 38988 18896
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 34704 18751 34756 18760
rect 34704 18717 34713 18751
rect 34713 18717 34747 18751
rect 34747 18717 34756 18751
rect 34704 18708 34756 18717
rect 35440 18708 35492 18760
rect 35808 18751 35860 18760
rect 35808 18717 35817 18751
rect 35817 18717 35851 18751
rect 35851 18717 35860 18751
rect 35808 18708 35860 18717
rect 37924 18819 37976 18828
rect 37924 18785 37933 18819
rect 37933 18785 37967 18819
rect 37967 18785 37976 18819
rect 37924 18776 37976 18785
rect 38292 18819 38344 18828
rect 38292 18785 38301 18819
rect 38301 18785 38335 18819
rect 38335 18785 38344 18819
rect 38292 18776 38344 18785
rect 40408 18776 40460 18828
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17224 18640 17276 18692
rect 17592 18683 17644 18692
rect 17592 18649 17601 18683
rect 17601 18649 17635 18683
rect 17635 18649 17644 18683
rect 17592 18640 17644 18649
rect 18880 18640 18932 18692
rect 19432 18640 19484 18692
rect 22100 18640 22152 18692
rect 29000 18640 29052 18692
rect 29368 18640 29420 18692
rect 17960 18572 18012 18624
rect 19984 18572 20036 18624
rect 21916 18615 21968 18624
rect 21916 18581 21925 18615
rect 21925 18581 21959 18615
rect 21959 18581 21968 18615
rect 21916 18572 21968 18581
rect 24676 18572 24728 18624
rect 26608 18572 26660 18624
rect 37556 18572 37608 18624
rect 37832 18683 37884 18692
rect 37832 18649 37841 18683
rect 37841 18649 37875 18683
rect 37875 18649 37884 18683
rect 37832 18640 37884 18649
rect 38752 18640 38804 18692
rect 39212 18708 39264 18760
rect 39304 18751 39356 18760
rect 39304 18717 39313 18751
rect 39313 18717 39347 18751
rect 39347 18717 39356 18751
rect 39304 18708 39356 18717
rect 40224 18640 40276 18692
rect 41236 18751 41288 18760
rect 41236 18717 41245 18751
rect 41245 18717 41279 18751
rect 41279 18717 41288 18751
rect 41236 18708 41288 18717
rect 42708 18844 42760 18896
rect 41880 18708 41932 18760
rect 41972 18751 42024 18760
rect 41972 18717 41981 18751
rect 41981 18717 42015 18751
rect 42015 18717 42024 18751
rect 41972 18708 42024 18717
rect 42984 18708 43036 18760
rect 43076 18751 43128 18760
rect 43076 18717 43085 18751
rect 43085 18717 43119 18751
rect 43119 18717 43128 18751
rect 43076 18708 43128 18717
rect 43628 18640 43680 18692
rect 38660 18615 38712 18624
rect 38660 18581 38669 18615
rect 38669 18581 38703 18615
rect 38703 18581 38712 18615
rect 38660 18572 38712 18581
rect 39672 18615 39724 18624
rect 39672 18581 39681 18615
rect 39681 18581 39715 18615
rect 39715 18581 39724 18615
rect 39672 18572 39724 18581
rect 40776 18615 40828 18624
rect 40776 18581 40785 18615
rect 40785 18581 40819 18615
rect 40819 18581 40828 18615
rect 40776 18572 40828 18581
rect 41604 18572 41656 18624
rect 43444 18572 43496 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2228 18368 2280 18420
rect 3148 18368 3200 18420
rect 4712 18300 4764 18352
rect 7380 18368 7432 18420
rect 9220 18368 9272 18420
rect 10140 18368 10192 18420
rect 10784 18368 10836 18420
rect 10876 18368 10928 18420
rect 12348 18411 12400 18420
rect 12348 18377 12357 18411
rect 12357 18377 12391 18411
rect 12391 18377 12400 18411
rect 12348 18368 12400 18377
rect 12808 18368 12860 18420
rect 17592 18368 17644 18420
rect 8484 18300 8536 18352
rect 9036 18300 9088 18352
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 14372 18300 14424 18352
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 3700 18207 3752 18216
rect 3700 18173 3709 18207
rect 3709 18173 3743 18207
rect 3743 18173 3752 18207
rect 3700 18164 3752 18173
rect 6092 18096 6144 18148
rect 7840 18164 7892 18216
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 3332 18028 3384 18080
rect 4620 18028 4672 18080
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 10784 18028 10836 18080
rect 16580 18232 16632 18284
rect 19984 18368 20036 18420
rect 20444 18300 20496 18352
rect 20812 18300 20864 18352
rect 19248 18232 19300 18284
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 23388 18368 23440 18420
rect 23756 18368 23808 18420
rect 24032 18300 24084 18352
rect 24676 18300 24728 18352
rect 26240 18368 26292 18420
rect 37924 18368 37976 18420
rect 38292 18368 38344 18420
rect 38660 18368 38712 18420
rect 38844 18368 38896 18420
rect 39580 18368 39632 18420
rect 39672 18368 39724 18420
rect 40776 18368 40828 18420
rect 41236 18368 41288 18420
rect 43628 18411 43680 18420
rect 43628 18377 43637 18411
rect 43637 18377 43671 18411
rect 43671 18377 43680 18411
rect 43628 18368 43680 18377
rect 25136 18300 25188 18352
rect 25688 18343 25740 18352
rect 25688 18309 25697 18343
rect 25697 18309 25731 18343
rect 25731 18309 25740 18343
rect 25688 18300 25740 18309
rect 19064 18164 19116 18216
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 20720 18164 20772 18216
rect 22836 18164 22888 18216
rect 23480 18164 23532 18216
rect 25596 18232 25648 18284
rect 29184 18232 29236 18284
rect 29644 18275 29696 18284
rect 29644 18241 29653 18275
rect 29653 18241 29687 18275
rect 29687 18241 29696 18275
rect 29644 18232 29696 18241
rect 30104 18275 30156 18284
rect 30104 18241 30113 18275
rect 30113 18241 30147 18275
rect 30147 18241 30156 18275
rect 30104 18232 30156 18241
rect 27068 18164 27120 18216
rect 30196 18207 30248 18216
rect 30196 18173 30205 18207
rect 30205 18173 30239 18207
rect 30239 18173 30248 18207
rect 30196 18164 30248 18173
rect 31668 18164 31720 18216
rect 35716 18164 35768 18216
rect 37464 18164 37516 18216
rect 39396 18232 39448 18284
rect 39672 18232 39724 18284
rect 42340 18300 42392 18352
rect 41604 18275 41656 18284
rect 41604 18241 41613 18275
rect 41613 18241 41647 18275
rect 41647 18241 41656 18275
rect 41604 18232 41656 18241
rect 41880 18275 41932 18284
rect 41880 18241 41889 18275
rect 41889 18241 41923 18275
rect 41923 18241 41932 18275
rect 41880 18232 41932 18241
rect 41972 18232 42024 18284
rect 43352 18275 43404 18284
rect 43352 18241 43361 18275
rect 43361 18241 43395 18275
rect 43395 18241 43404 18275
rect 43352 18232 43404 18241
rect 37188 18096 37240 18148
rect 44180 18207 44232 18216
rect 44180 18173 44189 18207
rect 44189 18173 44223 18207
rect 44223 18173 44232 18207
rect 44180 18164 44232 18173
rect 39120 18096 39172 18148
rect 39396 18096 39448 18148
rect 20628 18028 20680 18080
rect 21640 18071 21692 18080
rect 21640 18037 21649 18071
rect 21649 18037 21683 18071
rect 21683 18037 21692 18071
rect 21640 18028 21692 18037
rect 25872 18071 25924 18080
rect 25872 18037 25881 18071
rect 25881 18037 25915 18071
rect 25915 18037 25924 18071
rect 25872 18028 25924 18037
rect 26056 18028 26108 18080
rect 26240 18028 26292 18080
rect 30380 18028 30432 18080
rect 34704 18028 34756 18080
rect 35992 18028 36044 18080
rect 37280 18028 37332 18080
rect 37372 18071 37424 18080
rect 37372 18037 37381 18071
rect 37381 18037 37415 18071
rect 37415 18037 37424 18071
rect 37372 18028 37424 18037
rect 38936 18028 38988 18080
rect 39580 18028 39632 18080
rect 42800 18071 42852 18080
rect 42800 18037 42809 18071
rect 42809 18037 42843 18071
rect 42843 18037 42852 18071
rect 42800 18028 42852 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3700 17824 3752 17876
rect 9496 17824 9548 17876
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 7012 17688 7064 17740
rect 7656 17688 7708 17740
rect 11888 17867 11940 17876
rect 11888 17833 11897 17867
rect 11897 17833 11931 17867
rect 11931 17833 11940 17867
rect 11888 17824 11940 17833
rect 12992 17824 13044 17876
rect 12440 17756 12492 17808
rect 14924 17756 14976 17808
rect 17316 17756 17368 17808
rect 20720 17867 20772 17876
rect 20720 17833 20729 17867
rect 20729 17833 20763 17867
rect 20763 17833 20772 17867
rect 20720 17824 20772 17833
rect 13452 17688 13504 17740
rect 17868 17688 17920 17740
rect 2780 17620 2832 17672
rect 4712 17620 4764 17672
rect 6184 17552 6236 17604
rect 6460 17595 6512 17604
rect 6460 17561 6469 17595
rect 6469 17561 6503 17595
rect 6503 17561 6512 17595
rect 6460 17552 6512 17561
rect 6552 17552 6604 17604
rect 9036 17552 9088 17604
rect 10324 17595 10376 17604
rect 10324 17561 10333 17595
rect 10333 17561 10367 17595
rect 10367 17561 10376 17595
rect 10324 17552 10376 17561
rect 4344 17527 4396 17536
rect 4344 17493 4353 17527
rect 4353 17493 4387 17527
rect 4387 17493 4396 17527
rect 4344 17484 4396 17493
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 8668 17484 8720 17536
rect 10784 17552 10836 17604
rect 14372 17620 14424 17672
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 14648 17620 14700 17672
rect 16304 17552 16356 17604
rect 17592 17552 17644 17604
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 13452 17484 13504 17536
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 18880 17484 18932 17536
rect 21916 17824 21968 17876
rect 25872 17824 25924 17876
rect 27344 17824 27396 17876
rect 26240 17756 26292 17808
rect 21456 17620 21508 17672
rect 21640 17688 21692 17740
rect 21732 17620 21784 17672
rect 25780 17688 25832 17740
rect 27436 17756 27488 17808
rect 27620 17756 27672 17808
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 25596 17620 25648 17672
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 26332 17620 26384 17672
rect 27528 17620 27580 17672
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 30104 17824 30156 17876
rect 38752 17867 38804 17876
rect 38752 17833 38761 17867
rect 38761 17833 38795 17867
rect 38795 17833 38804 17867
rect 38752 17824 38804 17833
rect 40224 17824 40276 17876
rect 30012 17756 30064 17808
rect 30380 17756 30432 17808
rect 29184 17663 29236 17672
rect 29184 17629 29193 17663
rect 29193 17629 29227 17663
rect 29227 17629 29236 17663
rect 29184 17620 29236 17629
rect 27344 17484 27396 17536
rect 27620 17527 27672 17536
rect 27620 17493 27629 17527
rect 27629 17493 27663 17527
rect 27663 17493 27672 17527
rect 27620 17484 27672 17493
rect 27804 17527 27856 17536
rect 27804 17493 27813 17527
rect 27813 17493 27847 17527
rect 27847 17493 27856 17527
rect 27804 17484 27856 17493
rect 29552 17663 29604 17672
rect 29552 17629 29561 17663
rect 29561 17629 29595 17663
rect 29595 17629 29604 17663
rect 29552 17620 29604 17629
rect 30288 17688 30340 17740
rect 30104 17620 30156 17672
rect 33508 17756 33560 17808
rect 31576 17688 31628 17740
rect 31944 17620 31996 17672
rect 32220 17620 32272 17672
rect 32312 17620 32364 17672
rect 37280 17731 37332 17740
rect 37280 17697 37289 17731
rect 37289 17697 37323 17731
rect 37323 17697 37332 17731
rect 37280 17688 37332 17697
rect 33600 17620 33652 17672
rect 37004 17663 37056 17672
rect 31116 17552 31168 17604
rect 29644 17484 29696 17536
rect 30012 17484 30064 17536
rect 32404 17484 32456 17536
rect 35992 17484 36044 17536
rect 37004 17629 37013 17663
rect 37013 17629 37047 17663
rect 37047 17629 37056 17663
rect 37004 17620 37056 17629
rect 39396 17620 39448 17672
rect 40132 17595 40184 17604
rect 40132 17561 40141 17595
rect 40141 17561 40175 17595
rect 40175 17561 40184 17595
rect 40132 17552 40184 17561
rect 42340 17688 42392 17740
rect 42800 17824 42852 17876
rect 42800 17688 42852 17740
rect 44180 17688 44232 17740
rect 37188 17484 37240 17536
rect 39028 17527 39080 17536
rect 39028 17493 39037 17527
rect 39037 17493 39071 17527
rect 39071 17493 39080 17527
rect 39028 17484 39080 17493
rect 39948 17484 40000 17536
rect 40868 17484 40920 17536
rect 42524 17663 42576 17672
rect 42524 17629 42533 17663
rect 42533 17629 42567 17663
rect 42567 17629 42576 17663
rect 42524 17620 42576 17629
rect 42156 17484 42208 17536
rect 42432 17484 42484 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4344 17280 4396 17332
rect 5080 17280 5132 17332
rect 6460 17280 6512 17332
rect 8024 17212 8076 17264
rect 8944 17280 8996 17332
rect 10324 17280 10376 17332
rect 6920 17144 6972 17196
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 16580 17280 16632 17332
rect 17868 17280 17920 17332
rect 18880 17280 18932 17332
rect 16396 17255 16448 17264
rect 16396 17221 16405 17255
rect 16405 17221 16439 17255
rect 16439 17221 16448 17255
rect 16396 17212 16448 17221
rect 7012 17076 7064 17128
rect 8944 17076 8996 17128
rect 11980 17119 12032 17128
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 12900 17144 12952 17196
rect 13452 17144 13504 17196
rect 15476 17144 15528 17196
rect 12440 17076 12492 17128
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 14924 17076 14976 17128
rect 4712 16940 4764 16992
rect 6552 16940 6604 16992
rect 10600 16983 10652 16992
rect 10600 16949 10609 16983
rect 10609 16949 10643 16983
rect 10643 16949 10652 16983
rect 10600 16940 10652 16949
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 27804 17280 27856 17332
rect 29552 17323 29604 17332
rect 29552 17289 29561 17323
rect 29561 17289 29595 17323
rect 29595 17289 29604 17323
rect 29552 17280 29604 17289
rect 30196 17280 30248 17332
rect 20444 17255 20496 17264
rect 20444 17221 20453 17255
rect 20453 17221 20487 17255
rect 20487 17221 20496 17255
rect 20444 17212 20496 17221
rect 20812 17212 20864 17264
rect 22560 17212 22612 17264
rect 20536 17144 20588 17196
rect 20628 17144 20680 17196
rect 25688 17144 25740 17196
rect 27068 17187 27120 17196
rect 27068 17153 27077 17187
rect 27077 17153 27111 17187
rect 27111 17153 27120 17187
rect 27068 17144 27120 17153
rect 31576 17212 31628 17264
rect 29184 17144 29236 17196
rect 30472 17144 30524 17196
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 18328 17076 18380 17128
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 22192 17076 22244 17128
rect 26056 17119 26108 17128
rect 26056 17085 26065 17119
rect 26065 17085 26099 17119
rect 26099 17085 26108 17119
rect 26056 17076 26108 17085
rect 30104 17076 30156 17128
rect 30196 17076 30248 17128
rect 30564 17119 30616 17128
rect 30564 17085 30573 17119
rect 30573 17085 30607 17119
rect 30607 17085 30616 17119
rect 30564 17076 30616 17085
rect 32220 17187 32272 17196
rect 32220 17153 32229 17187
rect 32229 17153 32263 17187
rect 32263 17153 32272 17187
rect 32220 17144 32272 17153
rect 32404 17187 32456 17196
rect 32404 17153 32413 17187
rect 32413 17153 32447 17187
rect 32447 17153 32456 17187
rect 32404 17144 32456 17153
rect 34152 17280 34204 17332
rect 34428 17280 34480 17332
rect 37372 17280 37424 17332
rect 38844 17280 38896 17332
rect 39120 17280 39172 17332
rect 39212 17323 39264 17332
rect 39212 17289 39221 17323
rect 39221 17289 39255 17323
rect 39255 17289 39264 17323
rect 39212 17280 39264 17289
rect 39396 17280 39448 17332
rect 32312 17076 32364 17128
rect 33508 17187 33560 17196
rect 33508 17153 33517 17187
rect 33517 17153 33551 17187
rect 33551 17153 33560 17187
rect 33508 17144 33560 17153
rect 33600 17144 33652 17196
rect 33784 17144 33836 17196
rect 34152 17187 34204 17196
rect 34152 17153 34161 17187
rect 34161 17153 34195 17187
rect 34195 17153 34204 17187
rect 34152 17144 34204 17153
rect 34336 17144 34388 17196
rect 34704 17187 34756 17196
rect 34704 17153 34713 17187
rect 34713 17153 34747 17187
rect 34747 17153 34756 17187
rect 34704 17144 34756 17153
rect 37004 17144 37056 17196
rect 40224 17255 40276 17264
rect 40224 17221 40233 17255
rect 40233 17221 40267 17255
rect 40267 17221 40276 17255
rect 40224 17212 40276 17221
rect 37188 17076 37240 17128
rect 38752 17076 38804 17128
rect 32128 17008 32180 17060
rect 17592 16940 17644 16992
rect 18512 16940 18564 16992
rect 22652 16940 22704 16992
rect 22836 16940 22888 16992
rect 30380 16940 30432 16992
rect 31392 16940 31444 16992
rect 39764 17144 39816 17196
rect 41604 17280 41656 17332
rect 42156 17212 42208 17264
rect 43536 17280 43588 17332
rect 44180 17212 44232 17264
rect 41880 17076 41932 17128
rect 42708 17076 42760 17128
rect 33048 16983 33100 16992
rect 33048 16949 33057 16983
rect 33057 16949 33091 16983
rect 33091 16949 33100 16983
rect 33048 16940 33100 16949
rect 33692 16940 33744 16992
rect 34520 16940 34572 16992
rect 41604 16983 41656 16992
rect 41604 16949 41613 16983
rect 41613 16949 41647 16983
rect 41647 16949 41656 16983
rect 41604 16940 41656 16949
rect 42064 16983 42116 16992
rect 42064 16949 42073 16983
rect 42073 16949 42107 16983
rect 42107 16949 42116 16983
rect 42064 16940 42116 16949
rect 42156 16940 42208 16992
rect 43444 16983 43496 16992
rect 43444 16949 43453 16983
rect 43453 16949 43487 16983
rect 43487 16949 43496 16983
rect 43444 16940 43496 16949
rect 44272 16940 44324 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8944 16779 8996 16788
rect 8944 16745 8953 16779
rect 8953 16745 8987 16779
rect 8987 16745 8996 16779
rect 8944 16736 8996 16745
rect 9036 16736 9088 16788
rect 10600 16736 10652 16788
rect 12440 16736 12492 16788
rect 13084 16736 13136 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 17224 16736 17276 16788
rect 18052 16736 18104 16788
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 22192 16736 22244 16788
rect 27620 16736 27672 16788
rect 30104 16736 30156 16788
rect 33048 16736 33100 16788
rect 34152 16736 34204 16788
rect 38844 16736 38896 16788
rect 39028 16736 39080 16788
rect 40132 16736 40184 16788
rect 40868 16736 40920 16788
rect 42708 16779 42760 16788
rect 42708 16745 42717 16779
rect 42717 16745 42751 16779
rect 42751 16745 42760 16779
rect 42708 16736 42760 16745
rect 19340 16668 19392 16720
rect 9312 16532 9364 16584
rect 18328 16600 18380 16652
rect 22652 16668 22704 16720
rect 20352 16600 20404 16652
rect 21732 16600 21784 16652
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 23480 16600 23532 16652
rect 26608 16600 26660 16652
rect 27160 16600 27212 16652
rect 6828 16464 6880 16516
rect 7012 16396 7064 16448
rect 11704 16507 11756 16516
rect 11704 16473 11713 16507
rect 11713 16473 11747 16507
rect 11747 16473 11756 16507
rect 11704 16464 11756 16473
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 17592 16532 17644 16584
rect 15108 16396 15160 16448
rect 16580 16396 16632 16448
rect 20444 16532 20496 16584
rect 19984 16396 20036 16448
rect 22836 16532 22888 16584
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 23848 16396 23900 16448
rect 25688 16532 25740 16584
rect 26332 16532 26384 16584
rect 29552 16532 29604 16584
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 24676 16396 24728 16448
rect 29644 16396 29696 16448
rect 30104 16396 30156 16448
rect 32128 16600 32180 16652
rect 30472 16532 30524 16584
rect 30656 16532 30708 16584
rect 31852 16532 31904 16584
rect 32220 16532 32272 16584
rect 33508 16668 33560 16720
rect 33600 16668 33652 16720
rect 34520 16668 34572 16720
rect 30564 16396 30616 16448
rect 30840 16464 30892 16516
rect 32956 16464 33008 16516
rect 31484 16396 31536 16448
rect 34704 16532 34756 16584
rect 39948 16600 40000 16652
rect 42524 16600 42576 16652
rect 33784 16396 33836 16448
rect 33876 16396 33928 16448
rect 37464 16464 37516 16516
rect 41512 16464 41564 16516
rect 42248 16464 42300 16516
rect 35716 16439 35768 16448
rect 35716 16405 35725 16439
rect 35725 16405 35759 16439
rect 35759 16405 35768 16439
rect 35716 16396 35768 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2780 16192 2832 16244
rect 4712 16192 4764 16244
rect 6552 16124 6604 16176
rect 9588 16192 9640 16244
rect 11704 16192 11756 16244
rect 9312 16124 9364 16176
rect 9680 16124 9732 16176
rect 5724 16056 5776 16108
rect 3332 15852 3384 15904
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6000 16031 6052 16040
rect 6000 15997 6009 16031
rect 6009 15997 6043 16031
rect 6043 15997 6052 16031
rect 6000 15988 6052 15997
rect 8300 15988 8352 16040
rect 13084 16192 13136 16244
rect 16580 16192 16632 16244
rect 12440 16056 12492 16108
rect 15476 16124 15528 16176
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18328 16192 18380 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 23756 16192 23808 16244
rect 24492 16192 24544 16244
rect 26884 16192 26936 16244
rect 31852 16192 31904 16244
rect 32956 16192 33008 16244
rect 17960 16124 18012 16176
rect 25688 16124 25740 16176
rect 29276 16124 29328 16176
rect 30840 16124 30892 16176
rect 35716 16192 35768 16244
rect 42524 16192 42576 16244
rect 8668 15988 8720 16040
rect 12716 16031 12768 16040
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 12716 15988 12768 15997
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 16304 15988 16356 16040
rect 18788 16056 18840 16108
rect 21824 16056 21876 16108
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 26700 16056 26752 16108
rect 26976 16099 27028 16108
rect 26976 16065 26985 16099
rect 26985 16065 27019 16099
rect 27019 16065 27028 16099
rect 26976 16056 27028 16065
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 20076 15988 20128 16040
rect 23848 15988 23900 16040
rect 22652 15920 22704 15972
rect 22928 15920 22980 15972
rect 5632 15852 5684 15904
rect 13636 15852 13688 15904
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 22468 15852 22520 15904
rect 29092 15920 29144 15972
rect 27252 15852 27304 15904
rect 29276 15895 29328 15904
rect 29276 15861 29285 15895
rect 29285 15861 29319 15895
rect 29319 15861 29328 15895
rect 29276 15852 29328 15861
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 30288 16056 30340 16108
rect 29644 15988 29696 16040
rect 30104 15988 30156 16040
rect 30656 15988 30708 16040
rect 30840 15988 30892 16040
rect 31300 16056 31352 16108
rect 31484 16097 31536 16108
rect 31484 16063 31493 16097
rect 31493 16063 31527 16097
rect 31527 16063 31536 16097
rect 31484 16056 31536 16063
rect 31576 15988 31628 16040
rect 32220 16056 32272 16108
rect 31024 15920 31076 15972
rect 31852 15963 31904 15972
rect 31852 15929 31861 15963
rect 31861 15929 31895 15963
rect 31895 15929 31904 15963
rect 31852 15920 31904 15929
rect 33232 16099 33284 16108
rect 33232 16065 33241 16099
rect 33241 16065 33275 16099
rect 33275 16065 33284 16099
rect 33232 16056 33284 16065
rect 33324 16099 33376 16108
rect 33324 16065 33333 16099
rect 33333 16065 33367 16099
rect 33367 16065 33376 16099
rect 33324 16056 33376 16065
rect 33876 16099 33928 16108
rect 33876 16065 33885 16099
rect 33885 16065 33919 16099
rect 33919 16065 33928 16099
rect 33876 16056 33928 16065
rect 34060 16099 34112 16108
rect 34060 16065 34095 16099
rect 34095 16065 34112 16099
rect 34060 16056 34112 16065
rect 40500 16099 40552 16108
rect 40500 16065 40509 16099
rect 40509 16065 40543 16099
rect 40543 16065 40552 16099
rect 40500 16056 40552 16065
rect 43996 16099 44048 16108
rect 43996 16065 44005 16099
rect 44005 16065 44039 16099
rect 44039 16065 44048 16099
rect 43996 16056 44048 16065
rect 34612 15988 34664 16040
rect 39764 15988 39816 16040
rect 41604 15988 41656 16040
rect 42156 15988 42208 16040
rect 33508 15895 33560 15904
rect 33508 15861 33517 15895
rect 33517 15861 33551 15895
rect 33551 15861 33560 15895
rect 33508 15852 33560 15861
rect 33600 15895 33652 15904
rect 33600 15861 33609 15895
rect 33609 15861 33643 15895
rect 33643 15861 33652 15895
rect 33600 15852 33652 15861
rect 40224 15895 40276 15904
rect 40224 15861 40233 15895
rect 40233 15861 40267 15895
rect 40267 15861 40276 15895
rect 40224 15852 40276 15861
rect 44180 15895 44232 15904
rect 44180 15861 44189 15895
rect 44189 15861 44223 15895
rect 44223 15861 44232 15895
rect 44180 15852 44232 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 5356 15648 5408 15700
rect 6000 15648 6052 15700
rect 11796 15648 11848 15700
rect 13544 15648 13596 15700
rect 3332 15512 3384 15564
rect 13636 15580 13688 15632
rect 22468 15648 22520 15700
rect 7012 15512 7064 15564
rect 8300 15512 8352 15564
rect 12900 15512 12952 15564
rect 17684 15512 17736 15564
rect 18328 15512 18380 15564
rect 23112 15648 23164 15700
rect 26516 15648 26568 15700
rect 26976 15648 27028 15700
rect 29276 15648 29328 15700
rect 30104 15648 30156 15700
rect 31024 15648 31076 15700
rect 31300 15648 31352 15700
rect 6736 15444 6788 15496
rect 12348 15444 12400 15496
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 4712 15376 4764 15428
rect 10508 15419 10560 15428
rect 10508 15385 10517 15419
rect 10517 15385 10551 15419
rect 10551 15385 10560 15419
rect 10508 15376 10560 15385
rect 11060 15376 11112 15428
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 12440 15308 12492 15360
rect 15108 15444 15160 15496
rect 20352 15512 20404 15564
rect 20444 15512 20496 15564
rect 21548 15512 21600 15564
rect 23480 15512 23532 15564
rect 26608 15512 26660 15564
rect 33232 15648 33284 15700
rect 33324 15648 33376 15700
rect 33784 15648 33836 15700
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 26332 15487 26384 15496
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 26516 15444 26568 15496
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 19984 15376 20036 15428
rect 20352 15419 20404 15428
rect 20352 15385 20361 15419
rect 20361 15385 20395 15419
rect 20395 15385 20404 15419
rect 20352 15376 20404 15385
rect 20168 15308 20220 15360
rect 23204 15376 23256 15428
rect 33508 15512 33560 15564
rect 27804 15376 27856 15428
rect 24216 15308 24268 15360
rect 24676 15308 24728 15360
rect 26240 15351 26292 15360
rect 26240 15317 26249 15351
rect 26249 15317 26283 15351
rect 26283 15317 26292 15351
rect 26240 15308 26292 15317
rect 27528 15308 27580 15360
rect 29368 15444 29420 15496
rect 32772 15444 32824 15496
rect 33048 15487 33100 15496
rect 33048 15453 33057 15487
rect 33057 15453 33091 15487
rect 33091 15453 33100 15487
rect 33048 15444 33100 15453
rect 33876 15512 33928 15564
rect 33692 15487 33744 15496
rect 33692 15453 33701 15487
rect 33701 15453 33735 15487
rect 33735 15453 33744 15487
rect 33692 15444 33744 15453
rect 34612 15512 34664 15564
rect 38016 15648 38068 15700
rect 41512 15648 41564 15700
rect 42156 15648 42208 15700
rect 38016 15555 38068 15564
rect 38016 15521 38025 15555
rect 38025 15521 38059 15555
rect 38059 15521 38068 15555
rect 38016 15512 38068 15521
rect 39120 15512 39172 15564
rect 39948 15555 40000 15564
rect 39948 15521 39957 15555
rect 39957 15521 39991 15555
rect 39991 15521 40000 15555
rect 39948 15512 40000 15521
rect 40224 15555 40276 15564
rect 40224 15521 40233 15555
rect 40233 15521 40267 15555
rect 40267 15521 40276 15555
rect 40224 15512 40276 15521
rect 42524 15555 42576 15564
rect 42524 15521 42533 15555
rect 42533 15521 42567 15555
rect 42567 15521 42576 15555
rect 42524 15512 42576 15521
rect 35348 15487 35400 15496
rect 35348 15453 35357 15487
rect 35357 15453 35391 15487
rect 35391 15453 35400 15487
rect 35348 15444 35400 15453
rect 35440 15351 35492 15360
rect 35440 15317 35449 15351
rect 35449 15317 35483 15351
rect 35483 15317 35492 15351
rect 35440 15308 35492 15317
rect 37188 15376 37240 15428
rect 38108 15308 38160 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 39304 15487 39356 15496
rect 39304 15453 39313 15487
rect 39313 15453 39347 15487
rect 39347 15453 39356 15487
rect 39304 15444 39356 15453
rect 39580 15444 39632 15496
rect 41604 15444 41656 15496
rect 42064 15444 42116 15496
rect 40868 15376 40920 15428
rect 42800 15419 42852 15428
rect 42800 15385 42809 15419
rect 42809 15385 42843 15419
rect 42843 15385 42852 15419
rect 42800 15376 42852 15385
rect 43352 15376 43404 15428
rect 44272 15351 44324 15360
rect 44272 15317 44281 15351
rect 44281 15317 44315 15351
rect 44315 15317 44324 15351
rect 44272 15308 44324 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 6736 15104 6788 15156
rect 10508 15104 10560 15156
rect 12072 15104 12124 15156
rect 18328 15104 18380 15156
rect 20076 15104 20128 15156
rect 20352 15104 20404 15156
rect 3792 15036 3844 15088
rect 9036 15079 9088 15088
rect 9036 15045 9045 15079
rect 9045 15045 9079 15079
rect 9079 15045 9088 15079
rect 9036 15036 9088 15045
rect 9680 15036 9732 15088
rect 3332 14968 3384 15020
rect 4712 14968 4764 15020
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 8300 14968 8352 15020
rect 20444 15036 20496 15088
rect 21180 15104 21232 15156
rect 5632 14943 5684 14952
rect 5632 14909 5641 14943
rect 5641 14909 5675 14943
rect 5675 14909 5684 14943
rect 5632 14900 5684 14909
rect 6368 14832 6420 14884
rect 8760 14832 8812 14884
rect 14188 14832 14240 14884
rect 16488 14832 16540 14884
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 12256 14764 12308 14816
rect 17132 14764 17184 14816
rect 18512 14900 18564 14952
rect 18696 14900 18748 14952
rect 20076 14900 20128 14952
rect 22652 15104 22704 15156
rect 24216 15104 24268 15156
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 21364 14943 21416 14952
rect 21364 14909 21373 14943
rect 21373 14909 21407 14943
rect 21407 14909 21416 14943
rect 21364 14900 21416 14909
rect 21916 14968 21968 15020
rect 22376 14968 22428 15020
rect 26700 15036 26752 15088
rect 26976 15036 27028 15088
rect 27528 15036 27580 15088
rect 27804 15036 27856 15088
rect 22652 14900 22704 14952
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 25320 14900 25372 14952
rect 21916 14832 21968 14884
rect 22008 14832 22060 14884
rect 22192 14832 22244 14884
rect 26240 14832 26292 14884
rect 31484 14764 31536 14816
rect 32772 15011 32824 15020
rect 32772 14977 32781 15011
rect 32781 14977 32815 15011
rect 32815 14977 32824 15011
rect 32772 14968 32824 14977
rect 35992 15104 36044 15156
rect 38016 15104 38068 15156
rect 39580 15147 39632 15156
rect 39580 15113 39589 15147
rect 39589 15113 39623 15147
rect 39623 15113 39632 15147
rect 39580 15104 39632 15113
rect 43996 15104 44048 15156
rect 35440 15036 35492 15088
rect 33600 14900 33652 14952
rect 38200 15036 38252 15088
rect 37188 14900 37240 14952
rect 34612 14832 34664 14884
rect 43260 14968 43312 15020
rect 44272 15011 44324 15020
rect 44272 14977 44281 15011
rect 44281 14977 44315 15011
rect 44315 14977 44324 15011
rect 44272 14968 44324 14977
rect 42800 14900 42852 14952
rect 43076 14943 43128 14952
rect 43076 14909 43085 14943
rect 43085 14909 43119 14943
rect 43119 14909 43128 14943
rect 43076 14900 43128 14909
rect 43352 14832 43404 14884
rect 36084 14764 36136 14816
rect 36820 14807 36872 14816
rect 36820 14773 36829 14807
rect 36829 14773 36863 14807
rect 36863 14773 36872 14807
rect 36820 14764 36872 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 5172 14560 5224 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 14556 14560 14608 14612
rect 16028 14560 16080 14612
rect 7932 14492 7984 14544
rect 17132 14560 17184 14612
rect 19156 14560 19208 14612
rect 20076 14560 20128 14612
rect 11612 14356 11664 14408
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 22836 14492 22888 14544
rect 25228 14603 25280 14612
rect 25228 14569 25237 14603
rect 25237 14569 25271 14603
rect 25271 14569 25280 14603
rect 25228 14560 25280 14569
rect 25320 14560 25372 14612
rect 27160 14560 27212 14612
rect 25964 14492 26016 14544
rect 26516 14492 26568 14544
rect 13544 14424 13596 14476
rect 12532 14288 12584 14340
rect 14280 14356 14332 14408
rect 16488 14424 16540 14476
rect 19340 14424 19392 14476
rect 21088 14424 21140 14476
rect 22008 14424 22060 14476
rect 27436 14424 27488 14476
rect 27804 14467 27856 14476
rect 27804 14433 27813 14467
rect 27813 14433 27847 14467
rect 27847 14433 27856 14467
rect 27804 14424 27856 14433
rect 30472 14424 30524 14476
rect 35348 14560 35400 14612
rect 39948 14560 40000 14612
rect 43260 14603 43312 14612
rect 43260 14569 43269 14603
rect 43269 14569 43303 14603
rect 43303 14569 43312 14603
rect 43260 14560 43312 14569
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 15936 14356 15988 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 16212 14356 16264 14408
rect 16764 14356 16816 14408
rect 25412 14399 25464 14408
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 18880 14288 18932 14340
rect 21088 14288 21140 14340
rect 5724 14220 5776 14272
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 18236 14220 18288 14272
rect 18788 14220 18840 14272
rect 26240 14356 26292 14408
rect 31300 14356 31352 14408
rect 31668 14356 31720 14408
rect 26976 14288 27028 14340
rect 27252 14288 27304 14340
rect 35440 14399 35492 14408
rect 35440 14365 35449 14399
rect 35449 14365 35483 14399
rect 35483 14365 35492 14399
rect 35440 14356 35492 14365
rect 35716 14399 35768 14408
rect 35716 14365 35725 14399
rect 35725 14365 35759 14399
rect 35759 14365 35768 14399
rect 35716 14356 35768 14365
rect 36084 14356 36136 14408
rect 36820 14424 36872 14476
rect 43720 14467 43772 14476
rect 43720 14433 43729 14467
rect 43729 14433 43763 14467
rect 43763 14433 43772 14467
rect 43720 14424 43772 14433
rect 41604 14331 41656 14340
rect 41604 14297 41613 14331
rect 41613 14297 41647 14331
rect 41647 14297 41656 14331
rect 41604 14288 41656 14297
rect 42248 14288 42300 14340
rect 31300 14263 31352 14272
rect 31300 14229 31309 14263
rect 31309 14229 31343 14263
rect 31343 14229 31352 14263
rect 31300 14220 31352 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 5540 14016 5592 14068
rect 7288 14016 7340 14068
rect 12440 14016 12492 14068
rect 14464 14016 14516 14068
rect 15844 14016 15896 14068
rect 16120 14016 16172 14068
rect 7196 13880 7248 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 13084 13948 13136 14000
rect 13636 13948 13688 14000
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 13544 13880 13596 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 14188 13855 14240 13864
rect 11612 13744 11664 13796
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 14372 13855 14424 13864
rect 14372 13821 14381 13855
rect 14381 13821 14415 13855
rect 14415 13821 14424 13855
rect 14372 13812 14424 13821
rect 14556 13812 14608 13864
rect 15936 13948 15988 14000
rect 17224 14016 17276 14068
rect 18696 14016 18748 14068
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 18880 14016 18932 14068
rect 22560 14016 22612 14068
rect 22744 14059 22796 14068
rect 22744 14025 22753 14059
rect 22753 14025 22787 14059
rect 22787 14025 22796 14059
rect 22744 14016 22796 14025
rect 22836 14059 22888 14068
rect 22836 14025 22845 14059
rect 22845 14025 22879 14059
rect 22879 14025 22888 14059
rect 22836 14016 22888 14025
rect 30932 14016 30984 14068
rect 17132 13948 17184 14000
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 18052 13923 18104 13932
rect 12900 13744 12952 13796
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 18328 13923 18380 13932
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 6736 13676 6788 13728
rect 9588 13676 9640 13728
rect 11152 13676 11204 13728
rect 14464 13676 14516 13728
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17316 13812 17368 13864
rect 17224 13744 17276 13796
rect 18328 13889 18337 13923
rect 18337 13889 18371 13923
rect 18371 13889 18380 13923
rect 18328 13880 18380 13889
rect 20720 13948 20772 14000
rect 22376 13948 22428 14000
rect 24676 13948 24728 14000
rect 31116 13948 31168 14000
rect 35440 14016 35492 14068
rect 39948 14016 40000 14068
rect 41604 14016 41656 14068
rect 43352 14016 43404 14068
rect 43536 14016 43588 14068
rect 31576 13948 31628 14000
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 17040 13676 17092 13728
rect 17868 13676 17920 13728
rect 18972 13855 19024 13875
rect 18972 13823 18977 13855
rect 18977 13823 19011 13855
rect 19011 13823 19024 13855
rect 20076 13880 20128 13932
rect 22100 13923 22152 13932
rect 22100 13889 22127 13923
rect 22127 13889 22152 13923
rect 22100 13880 22152 13889
rect 23112 13880 23164 13932
rect 18880 13744 18932 13796
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 23480 13812 23532 13864
rect 22744 13744 22796 13796
rect 22836 13744 22888 13796
rect 29092 13880 29144 13932
rect 30012 13880 30064 13932
rect 30104 13880 30156 13932
rect 30932 13923 30984 13932
rect 30932 13889 30941 13923
rect 30941 13889 30975 13923
rect 30975 13889 30984 13923
rect 30932 13880 30984 13889
rect 29184 13812 29236 13864
rect 29736 13744 29788 13796
rect 30288 13855 30340 13864
rect 30288 13821 30297 13855
rect 30297 13821 30331 13855
rect 30331 13821 30340 13855
rect 30288 13812 30340 13821
rect 30656 13855 30708 13864
rect 30656 13821 30665 13855
rect 30665 13821 30699 13855
rect 30699 13821 30708 13855
rect 30656 13812 30708 13821
rect 30748 13855 30800 13864
rect 30748 13821 30757 13855
rect 30757 13821 30791 13855
rect 30791 13821 30800 13855
rect 30748 13812 30800 13821
rect 31024 13812 31076 13864
rect 31668 13880 31720 13932
rect 34796 13880 34848 13932
rect 35808 13923 35860 13932
rect 35808 13889 35817 13923
rect 35817 13889 35851 13923
rect 35851 13889 35860 13923
rect 35808 13880 35860 13889
rect 31484 13812 31536 13864
rect 36084 13812 36136 13864
rect 39028 13880 39080 13932
rect 43076 13880 43128 13932
rect 40132 13855 40184 13864
rect 40132 13821 40141 13855
rect 40141 13821 40175 13855
rect 40175 13821 40184 13855
rect 40132 13812 40184 13821
rect 40776 13855 40828 13864
rect 40776 13821 40785 13855
rect 40785 13821 40819 13855
rect 40819 13821 40828 13855
rect 40776 13812 40828 13821
rect 44088 13880 44140 13932
rect 30472 13744 30524 13796
rect 30932 13744 30984 13796
rect 22100 13676 22152 13728
rect 22468 13676 22520 13728
rect 22560 13676 22612 13728
rect 23388 13676 23440 13728
rect 23848 13676 23900 13728
rect 24768 13676 24820 13728
rect 26884 13676 26936 13728
rect 32956 13744 33008 13796
rect 31392 13676 31444 13728
rect 32680 13676 32732 13728
rect 34704 13719 34756 13728
rect 34704 13685 34713 13719
rect 34713 13685 34747 13719
rect 34747 13685 34756 13719
rect 34704 13676 34756 13685
rect 35900 13719 35952 13728
rect 35900 13685 35909 13719
rect 35909 13685 35943 13719
rect 35943 13685 35952 13719
rect 35900 13676 35952 13685
rect 36820 13676 36872 13728
rect 39580 13676 39632 13728
rect 43260 13719 43312 13728
rect 43260 13685 43269 13719
rect 43269 13685 43303 13719
rect 43303 13685 43312 13719
rect 43260 13676 43312 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7656 13472 7708 13524
rect 11980 13472 12032 13524
rect 12256 13472 12308 13524
rect 10324 13404 10376 13456
rect 13636 13472 13688 13524
rect 14372 13472 14424 13524
rect 5816 13336 5868 13388
rect 5908 13268 5960 13320
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 6736 13200 6788 13252
rect 6920 13132 6972 13184
rect 7196 13132 7248 13184
rect 11244 13336 11296 13388
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 14556 13404 14608 13456
rect 17040 13472 17092 13524
rect 17132 13515 17184 13524
rect 17132 13481 17141 13515
rect 17141 13481 17175 13515
rect 17175 13481 17184 13515
rect 17132 13472 17184 13481
rect 17224 13472 17276 13524
rect 12072 13268 12124 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 14096 13268 14148 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 17316 13404 17368 13456
rect 15108 13336 15160 13388
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 10140 13132 10192 13184
rect 11336 13200 11388 13252
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 11244 13132 11296 13184
rect 12256 13132 12308 13184
rect 15016 13268 15068 13320
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16580 13200 16632 13252
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 22284 13472 22336 13524
rect 23572 13472 23624 13524
rect 25412 13472 25464 13524
rect 26976 13472 27028 13524
rect 18052 13404 18104 13456
rect 20720 13447 20772 13456
rect 20720 13413 20729 13447
rect 20729 13413 20763 13447
rect 20763 13413 20772 13447
rect 20720 13404 20772 13413
rect 18512 13336 18564 13388
rect 21916 13336 21968 13388
rect 22560 13379 22612 13388
rect 22560 13345 22569 13379
rect 22569 13345 22603 13379
rect 22603 13345 22612 13379
rect 22560 13336 22612 13345
rect 18144 13268 18196 13320
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 23572 13336 23624 13388
rect 22744 13268 22796 13320
rect 23020 13311 23072 13320
rect 23020 13277 23029 13311
rect 23029 13277 23063 13311
rect 23063 13277 23072 13311
rect 23020 13268 23072 13277
rect 19340 13200 19392 13252
rect 21456 13200 21508 13252
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 23388 13268 23440 13320
rect 25596 13336 25648 13388
rect 27436 13379 27488 13388
rect 27436 13345 27445 13379
rect 27445 13345 27479 13379
rect 27479 13345 27488 13379
rect 27436 13336 27488 13345
rect 30748 13472 30800 13524
rect 31024 13515 31076 13524
rect 31024 13481 31033 13515
rect 31033 13481 31067 13515
rect 31067 13481 31076 13515
rect 31024 13472 31076 13481
rect 31208 13472 31260 13524
rect 31484 13472 31536 13524
rect 32956 13472 33008 13524
rect 30196 13404 30248 13456
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 17500 13132 17552 13184
rect 18052 13132 18104 13184
rect 22008 13175 22060 13184
rect 22008 13141 22017 13175
rect 22017 13141 22051 13175
rect 22051 13141 22060 13175
rect 22008 13132 22060 13141
rect 22100 13132 22152 13184
rect 22928 13132 22980 13184
rect 23664 13200 23716 13252
rect 24216 13311 24268 13320
rect 24216 13277 24225 13311
rect 24225 13277 24259 13311
rect 24259 13277 24268 13311
rect 24216 13268 24268 13277
rect 23940 13175 23992 13184
rect 23940 13141 23949 13175
rect 23949 13141 23983 13175
rect 23983 13141 23992 13175
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 29736 13311 29788 13320
rect 29736 13277 29745 13311
rect 29745 13277 29779 13311
rect 29779 13277 29788 13311
rect 29736 13268 29788 13277
rect 30104 13268 30156 13320
rect 32496 13379 32548 13388
rect 32496 13345 32505 13379
rect 32505 13345 32539 13379
rect 32539 13345 32548 13379
rect 32496 13336 32548 13345
rect 30380 13311 30432 13320
rect 30380 13277 30389 13311
rect 30389 13277 30423 13311
rect 30423 13277 30432 13311
rect 30380 13268 30432 13277
rect 30564 13311 30616 13320
rect 30564 13277 30573 13311
rect 30573 13277 30607 13311
rect 30607 13277 30616 13311
rect 30564 13268 30616 13277
rect 30656 13311 30708 13320
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 31392 13268 31444 13320
rect 31484 13311 31536 13320
rect 31484 13277 31493 13311
rect 31493 13277 31527 13311
rect 31527 13277 31536 13311
rect 31484 13268 31536 13277
rect 31668 13311 31720 13320
rect 31668 13277 31677 13311
rect 31677 13277 31711 13311
rect 31711 13277 31720 13311
rect 31668 13268 31720 13277
rect 27988 13200 28040 13252
rect 23940 13132 23992 13141
rect 26148 13132 26200 13184
rect 31760 13200 31812 13252
rect 29184 13175 29236 13184
rect 29184 13141 29193 13175
rect 29193 13141 29227 13175
rect 29227 13141 29236 13175
rect 29184 13132 29236 13141
rect 29552 13175 29604 13184
rect 29552 13141 29561 13175
rect 29561 13141 29595 13175
rect 29595 13141 29604 13175
rect 29552 13132 29604 13141
rect 30472 13132 30524 13184
rect 30932 13132 30984 13184
rect 35808 13472 35860 13524
rect 37556 13472 37608 13524
rect 39028 13472 39080 13524
rect 39120 13472 39172 13524
rect 40776 13472 40828 13524
rect 44088 13515 44140 13524
rect 44088 13481 44097 13515
rect 44097 13481 44131 13515
rect 44131 13481 44140 13515
rect 44088 13472 44140 13481
rect 36084 13336 36136 13388
rect 36176 13379 36228 13388
rect 36176 13345 36185 13379
rect 36185 13345 36219 13379
rect 36219 13345 36228 13379
rect 36176 13336 36228 13345
rect 38936 13336 38988 13388
rect 39120 13379 39172 13388
rect 39120 13345 39129 13379
rect 39129 13345 39163 13379
rect 39163 13345 39172 13379
rect 39120 13336 39172 13345
rect 39212 13336 39264 13388
rect 33324 13132 33376 13184
rect 36268 13200 36320 13252
rect 33968 13175 34020 13184
rect 33968 13141 33977 13175
rect 33977 13141 34011 13175
rect 34011 13141 34020 13175
rect 33968 13132 34020 13141
rect 34336 13132 34388 13184
rect 37556 13200 37608 13252
rect 38384 13200 38436 13252
rect 38568 13243 38620 13252
rect 38568 13209 38586 13243
rect 38586 13209 38620 13243
rect 38568 13200 38620 13209
rect 39304 13311 39356 13320
rect 39304 13277 39313 13311
rect 39313 13277 39347 13311
rect 39347 13277 39356 13311
rect 39304 13268 39356 13277
rect 39580 13268 39632 13320
rect 43260 13336 43312 13388
rect 38844 13200 38896 13252
rect 39672 13200 39724 13252
rect 43352 13200 43404 13252
rect 38660 13175 38712 13184
rect 38660 13141 38669 13175
rect 38669 13141 38703 13175
rect 38703 13141 38712 13175
rect 38660 13132 38712 13141
rect 39396 13132 39448 13184
rect 39488 13175 39540 13184
rect 39488 13141 39497 13175
rect 39497 13141 39531 13175
rect 39531 13141 39540 13175
rect 39488 13132 39540 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4620 12928 4672 12980
rect 6000 12928 6052 12980
rect 11428 12928 11480 12980
rect 12900 12928 12952 12980
rect 15384 12928 15436 12980
rect 16948 12928 17000 12980
rect 20904 12928 20956 12980
rect 4712 12860 4764 12912
rect 5724 12792 5776 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7656 12792 7708 12844
rect 9588 12860 9640 12912
rect 10232 12860 10284 12912
rect 10692 12860 10744 12912
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 6736 12724 6788 12776
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 8116 12724 8168 12776
rect 8576 12724 8628 12776
rect 10140 12724 10192 12776
rect 11888 12860 11940 12912
rect 13544 12860 13596 12912
rect 11520 12724 11572 12776
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 10968 12656 11020 12708
rect 12716 12724 12768 12776
rect 11796 12656 11848 12708
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 15476 12792 15528 12844
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 16396 12792 16448 12844
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18236 12792 18288 12801
rect 18788 12860 18840 12912
rect 18512 12792 18564 12844
rect 23020 12928 23072 12980
rect 23204 12928 23256 12980
rect 23756 12928 23808 12980
rect 24216 12928 24268 12980
rect 25504 12971 25556 12980
rect 25504 12937 25513 12971
rect 25513 12937 25547 12971
rect 25547 12937 25556 12971
rect 25504 12928 25556 12937
rect 14924 12656 14976 12708
rect 11244 12588 11296 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 15936 12656 15988 12708
rect 16028 12656 16080 12708
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 19984 12792 20036 12844
rect 20720 12792 20772 12844
rect 21916 12792 21968 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 19524 12767 19576 12776
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 22192 12792 22244 12844
rect 23388 12792 23440 12844
rect 19156 12656 19208 12708
rect 22836 12724 22888 12776
rect 22928 12724 22980 12776
rect 26240 12860 26292 12912
rect 26976 12971 27028 12980
rect 26976 12937 26985 12971
rect 26985 12937 27019 12971
rect 27019 12937 27028 12971
rect 26976 12928 27028 12937
rect 29552 12928 29604 12980
rect 30656 12928 30708 12980
rect 31300 12928 31352 12980
rect 31576 12928 31628 12980
rect 32772 12928 32824 12980
rect 36176 12928 36228 12980
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 25872 12835 25924 12844
rect 25872 12801 25881 12835
rect 25881 12801 25915 12835
rect 25915 12801 25924 12835
rect 25872 12792 25924 12801
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 26056 12767 26108 12776
rect 26056 12733 26065 12767
rect 26065 12733 26099 12767
rect 26099 12733 26108 12767
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 28816 12835 28868 12844
rect 28816 12801 28825 12835
rect 28825 12801 28859 12835
rect 28859 12801 28868 12835
rect 28816 12792 28868 12801
rect 29184 12835 29236 12844
rect 29184 12801 29193 12835
rect 29193 12801 29227 12835
rect 29227 12801 29236 12835
rect 29184 12792 29236 12801
rect 29920 12792 29972 12844
rect 30288 12792 30340 12844
rect 26056 12724 26108 12733
rect 26332 12656 26384 12708
rect 31208 12792 31260 12844
rect 32680 12903 32732 12912
rect 32680 12869 32689 12903
rect 32689 12869 32723 12903
rect 32723 12869 32732 12903
rect 32680 12860 32732 12869
rect 32312 12792 32364 12844
rect 32404 12835 32456 12844
rect 32404 12801 32413 12835
rect 32413 12801 32447 12835
rect 32447 12801 32456 12835
rect 32404 12792 32456 12801
rect 35900 12860 35952 12912
rect 32956 12835 33008 12844
rect 32956 12801 32965 12835
rect 32965 12801 32999 12835
rect 32999 12801 33008 12835
rect 32956 12792 33008 12801
rect 32864 12767 32916 12776
rect 32864 12733 32873 12767
rect 32873 12733 32907 12767
rect 32907 12733 32916 12767
rect 32864 12724 32916 12733
rect 16120 12588 16172 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 17132 12631 17184 12640
rect 17132 12597 17141 12631
rect 17141 12597 17175 12631
rect 17175 12597 17184 12631
rect 17132 12588 17184 12597
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 18144 12588 18196 12640
rect 18328 12588 18380 12640
rect 22192 12588 22244 12640
rect 23480 12588 23532 12640
rect 25596 12588 25648 12640
rect 26516 12588 26568 12640
rect 32404 12656 32456 12708
rect 33232 12792 33284 12844
rect 34336 12792 34388 12844
rect 34704 12792 34756 12844
rect 35716 12792 35768 12844
rect 34796 12724 34848 12776
rect 36084 12835 36136 12844
rect 36084 12801 36093 12835
rect 36093 12801 36127 12835
rect 36127 12801 36136 12835
rect 36084 12792 36136 12801
rect 38844 12928 38896 12980
rect 39212 12928 39264 12980
rect 39304 12928 39356 12980
rect 39488 12928 39540 12980
rect 40132 12928 40184 12980
rect 38568 12792 38620 12844
rect 39028 12792 39080 12844
rect 36268 12724 36320 12776
rect 37556 12767 37608 12776
rect 37556 12733 37565 12767
rect 37565 12733 37599 12767
rect 37599 12733 37608 12767
rect 37556 12724 37608 12733
rect 27160 12631 27212 12640
rect 27160 12597 27169 12631
rect 27169 12597 27203 12631
rect 27203 12597 27212 12631
rect 27160 12588 27212 12597
rect 27528 12631 27580 12640
rect 27528 12597 27537 12631
rect 27537 12597 27571 12631
rect 27571 12597 27580 12631
rect 27528 12588 27580 12597
rect 29000 12631 29052 12640
rect 29000 12597 29009 12631
rect 29009 12597 29043 12631
rect 29043 12597 29052 12631
rect 29000 12588 29052 12597
rect 31484 12588 31536 12640
rect 32128 12631 32180 12640
rect 32128 12597 32137 12631
rect 32137 12597 32171 12631
rect 32171 12597 32180 12631
rect 32128 12588 32180 12597
rect 32496 12588 32548 12640
rect 39580 12656 39632 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10324 12384 10376 12436
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 11612 12384 11664 12436
rect 10784 12316 10836 12368
rect 11704 12316 11756 12368
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 14832 12384 14884 12436
rect 15384 12384 15436 12436
rect 15844 12384 15896 12436
rect 17592 12384 17644 12436
rect 18696 12384 18748 12436
rect 19524 12384 19576 12436
rect 22100 12384 22152 12436
rect 23112 12384 23164 12436
rect 23572 12384 23624 12436
rect 12716 12316 12768 12368
rect 13820 12316 13872 12368
rect 6828 12112 6880 12164
rect 9772 12112 9824 12164
rect 9956 12155 10008 12164
rect 9956 12121 9965 12155
rect 9965 12121 9999 12155
rect 9999 12121 10008 12155
rect 9956 12112 10008 12121
rect 10600 12180 10652 12232
rect 11244 12180 11296 12232
rect 14004 12248 14056 12300
rect 13084 12180 13136 12232
rect 15108 12316 15160 12368
rect 15016 12248 15068 12300
rect 14096 12112 14148 12164
rect 5632 12044 5684 12096
rect 7656 12044 7708 12096
rect 10324 12044 10376 12096
rect 10416 12044 10468 12096
rect 11704 12044 11756 12096
rect 12532 12044 12584 12096
rect 14648 12044 14700 12096
rect 14740 12044 14792 12096
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 15752 12180 15804 12232
rect 16764 12180 16816 12232
rect 17776 12248 17828 12300
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 19432 12316 19484 12368
rect 19800 12359 19852 12368
rect 19800 12325 19809 12359
rect 19809 12325 19843 12359
rect 19843 12325 19852 12359
rect 19800 12316 19852 12325
rect 22468 12316 22520 12368
rect 26516 12384 26568 12436
rect 26608 12384 26660 12436
rect 27620 12384 27672 12436
rect 30564 12384 30616 12436
rect 18696 12180 18748 12232
rect 21916 12248 21968 12300
rect 23296 12248 23348 12300
rect 26332 12316 26384 12368
rect 25136 12248 25188 12300
rect 26056 12248 26108 12300
rect 26976 12248 27028 12300
rect 27068 12248 27120 12300
rect 27620 12248 27672 12300
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 21548 12180 21600 12232
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 29736 12248 29788 12300
rect 38200 12248 38252 12300
rect 18052 12112 18104 12164
rect 19156 12112 19208 12164
rect 16028 12044 16080 12096
rect 16212 12044 16264 12096
rect 16580 12044 16632 12096
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 19984 12112 20036 12164
rect 24308 12112 24360 12164
rect 20352 12044 20404 12096
rect 21732 12044 21784 12096
rect 21916 12044 21968 12096
rect 22652 12044 22704 12096
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 26240 12155 26292 12164
rect 26240 12121 26249 12155
rect 26249 12121 26283 12155
rect 26283 12121 26292 12155
rect 26240 12112 26292 12121
rect 27436 12112 27488 12164
rect 27620 12112 27672 12164
rect 29368 12223 29420 12232
rect 29368 12189 29377 12223
rect 29377 12189 29411 12223
rect 29411 12189 29420 12223
rect 29368 12180 29420 12189
rect 30104 12180 30156 12232
rect 30288 12180 30340 12232
rect 31116 12180 31168 12232
rect 33968 12180 34020 12232
rect 34520 12180 34572 12232
rect 34796 12180 34848 12232
rect 35072 12223 35124 12232
rect 35072 12189 35081 12223
rect 35081 12189 35115 12223
rect 35115 12189 35124 12223
rect 35072 12180 35124 12189
rect 40500 12112 40552 12164
rect 42524 12112 42576 12164
rect 34796 12044 34848 12096
rect 36084 12087 36136 12096
rect 36084 12053 36093 12087
rect 36093 12053 36127 12087
rect 36127 12053 36136 12087
rect 36084 12044 36136 12053
rect 39028 12044 39080 12096
rect 39672 12044 39724 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 10048 11840 10100 11892
rect 10692 11883 10744 11892
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 10876 11840 10928 11892
rect 9588 11704 9640 11756
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10416 11704 10468 11756
rect 5632 11636 5684 11688
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 10692 11704 10744 11756
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 11980 11840 12032 11892
rect 12348 11840 12400 11892
rect 12808 11840 12860 11892
rect 13084 11840 13136 11892
rect 10784 11636 10836 11688
rect 11428 11704 11480 11756
rect 12624 11704 12676 11756
rect 12716 11704 12768 11756
rect 10784 11500 10836 11552
rect 11060 11500 11112 11552
rect 11520 11568 11572 11620
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 12532 11500 12584 11552
rect 12716 11500 12768 11552
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 14556 11636 14608 11688
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 14096 11611 14148 11620
rect 14096 11577 14105 11611
rect 14105 11577 14139 11611
rect 14139 11577 14148 11611
rect 14096 11568 14148 11577
rect 15200 11636 15252 11688
rect 15568 11636 15620 11688
rect 15936 11636 15988 11688
rect 16764 11704 16816 11756
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 18972 11840 19024 11892
rect 22100 11883 22152 11892
rect 22100 11849 22109 11883
rect 22109 11849 22143 11883
rect 22143 11849 22152 11883
rect 22100 11840 22152 11849
rect 22468 11840 22520 11892
rect 24676 11840 24728 11892
rect 34428 11883 34480 11892
rect 34428 11849 34437 11883
rect 34437 11849 34471 11883
rect 34471 11849 34480 11883
rect 34428 11840 34480 11849
rect 34612 11883 34664 11892
rect 34612 11849 34639 11883
rect 34639 11849 34664 11883
rect 34612 11840 34664 11849
rect 35072 11840 35124 11892
rect 37556 11840 37608 11892
rect 16212 11636 16264 11688
rect 15660 11568 15712 11620
rect 16028 11568 16080 11620
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 20812 11636 20864 11688
rect 21088 11636 21140 11688
rect 22008 11636 22060 11688
rect 22560 11568 22612 11620
rect 23296 11704 23348 11756
rect 28816 11772 28868 11824
rect 24676 11747 24728 11756
rect 24676 11713 24685 11747
rect 24685 11713 24719 11747
rect 24719 11713 24728 11747
rect 24676 11704 24728 11713
rect 24952 11747 25004 11756
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 25596 11704 25648 11756
rect 27712 11704 27764 11756
rect 27436 11679 27488 11688
rect 27436 11645 27445 11679
rect 27445 11645 27479 11679
rect 27479 11645 27488 11679
rect 27436 11636 27488 11645
rect 27528 11679 27580 11688
rect 27528 11645 27537 11679
rect 27537 11645 27571 11679
rect 27571 11645 27580 11679
rect 27528 11636 27580 11645
rect 30748 11704 30800 11756
rect 31668 11704 31720 11756
rect 35348 11704 35400 11756
rect 32864 11636 32916 11688
rect 38660 11772 38712 11824
rect 36176 11679 36228 11688
rect 36176 11645 36185 11679
rect 36185 11645 36219 11679
rect 36219 11645 36228 11679
rect 36176 11636 36228 11645
rect 38476 11704 38528 11756
rect 24768 11568 24820 11620
rect 14648 11500 14700 11552
rect 22008 11500 22060 11552
rect 22468 11500 22520 11552
rect 22652 11500 22704 11552
rect 22836 11500 22888 11552
rect 23204 11500 23256 11552
rect 31576 11568 31628 11620
rect 32220 11568 32272 11620
rect 32956 11568 33008 11620
rect 29552 11500 29604 11552
rect 31300 11500 31352 11552
rect 36452 11568 36504 11620
rect 34704 11500 34756 11552
rect 38936 11500 38988 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7840 11296 7892 11348
rect 10968 11296 11020 11348
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 13084 11296 13136 11348
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7288 11024 7340 11076
rect 7656 11024 7708 11076
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 9680 11092 9732 11144
rect 10784 11092 10836 11144
rect 10968 11092 11020 11144
rect 11336 11160 11388 11212
rect 11888 11160 11940 11212
rect 9864 10956 9916 11008
rect 10416 10956 10468 11008
rect 10508 10956 10560 11008
rect 11336 11024 11388 11076
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 14556 11339 14608 11348
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 14648 11296 14700 11348
rect 15292 11296 15344 11348
rect 16028 11296 16080 11348
rect 18420 11296 18472 11348
rect 14740 11228 14792 11280
rect 19984 11296 20036 11348
rect 20444 11296 20496 11348
rect 21732 11296 21784 11348
rect 22284 11296 22336 11348
rect 24676 11296 24728 11348
rect 27252 11296 27304 11348
rect 29552 11339 29604 11348
rect 29552 11305 29561 11339
rect 29561 11305 29595 11339
rect 29595 11305 29604 11339
rect 29552 11296 29604 11305
rect 29920 11296 29972 11348
rect 32036 11296 32088 11348
rect 32588 11296 32640 11348
rect 32864 11296 32916 11348
rect 34704 11296 34756 11348
rect 34796 11296 34848 11348
rect 36452 11339 36504 11348
rect 36452 11305 36461 11339
rect 36461 11305 36495 11339
rect 36495 11305 36504 11339
rect 36452 11296 36504 11305
rect 38936 11339 38988 11348
rect 38936 11305 38945 11339
rect 38945 11305 38979 11339
rect 38979 11305 38988 11339
rect 38936 11296 38988 11305
rect 12532 11092 12584 11101
rect 12256 11024 12308 11076
rect 12992 11067 13044 11076
rect 12992 11033 13001 11067
rect 13001 11033 13035 11067
rect 13035 11033 13044 11067
rect 12992 11024 13044 11033
rect 13452 11092 13504 11144
rect 13544 11092 13596 11144
rect 13912 11024 13964 11076
rect 14188 11067 14240 11076
rect 14188 11033 14197 11067
rect 14197 11033 14231 11067
rect 14231 11033 14240 11067
rect 14188 11024 14240 11033
rect 14464 11092 14516 11144
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 15384 11203 15436 11212
rect 15384 11169 15393 11203
rect 15393 11169 15427 11203
rect 15427 11169 15436 11203
rect 15384 11160 15436 11169
rect 17224 11092 17276 11144
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18052 11160 18104 11212
rect 20260 11160 20312 11212
rect 16120 11024 16172 11076
rect 16764 11024 16816 11076
rect 17684 11024 17736 11076
rect 18420 11092 18472 11144
rect 18696 11092 18748 11144
rect 19248 11092 19300 11144
rect 19432 11092 19484 11144
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 20352 11092 20404 11144
rect 18144 11067 18196 11076
rect 18144 11033 18153 11067
rect 18153 11033 18187 11067
rect 18187 11033 18196 11067
rect 18144 11024 18196 11033
rect 21272 11092 21324 11144
rect 22744 11228 22796 11280
rect 23480 11228 23532 11280
rect 27620 11228 27672 11280
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 22100 11092 22152 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 22744 11092 22796 11144
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 12072 10956 12124 11008
rect 20628 11024 20680 11076
rect 20720 11024 20772 11076
rect 22192 11024 22244 11076
rect 19064 10999 19116 11008
rect 19064 10965 19073 10999
rect 19073 10965 19107 10999
rect 19107 10965 19116 10999
rect 19064 10956 19116 10965
rect 19432 10956 19484 11008
rect 24492 11092 24544 11144
rect 24952 11160 25004 11212
rect 27896 11135 27948 11144
rect 27896 11101 27905 11135
rect 27905 11101 27939 11135
rect 27939 11101 27948 11135
rect 27896 11092 27948 11101
rect 28632 11092 28684 11144
rect 29736 11135 29788 11144
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 29828 11092 29880 11101
rect 32680 11228 32732 11280
rect 31300 11203 31352 11212
rect 31300 11169 31309 11203
rect 31309 11169 31343 11203
rect 31343 11169 31352 11203
rect 31300 11160 31352 11169
rect 32588 11203 32640 11212
rect 32588 11169 32597 11203
rect 32597 11169 32631 11203
rect 32631 11169 32640 11203
rect 32588 11160 32640 11169
rect 33232 11160 33284 11212
rect 33784 11160 33836 11212
rect 31576 11135 31628 11144
rect 31576 11101 31585 11135
rect 31585 11101 31619 11135
rect 31619 11101 31628 11135
rect 31576 11092 31628 11101
rect 31668 11135 31720 11144
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 32036 11092 32088 11144
rect 32220 11092 32272 11144
rect 29460 11024 29512 11076
rect 30104 11024 30156 11076
rect 32496 11024 32548 11076
rect 22836 10956 22888 11008
rect 24308 10956 24360 11008
rect 25044 10956 25096 11008
rect 31116 10956 31168 11008
rect 31944 10956 31996 11008
rect 35348 11160 35400 11212
rect 41420 11228 41472 11280
rect 37280 11160 37332 11212
rect 38476 11160 38528 11212
rect 38660 11160 38712 11212
rect 42800 11160 42852 11212
rect 36268 11092 36320 11144
rect 37648 11092 37700 11144
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 38200 11092 38252 11144
rect 38568 11135 38620 11144
rect 38568 11101 38577 11135
rect 38577 11101 38611 11135
rect 38611 11101 38620 11135
rect 38568 11092 38620 11101
rect 39488 11135 39540 11144
rect 39488 11101 39497 11135
rect 39497 11101 39531 11135
rect 39531 11101 39540 11135
rect 39488 11092 39540 11101
rect 43996 11203 44048 11212
rect 43996 11169 44005 11203
rect 44005 11169 44039 11203
rect 44039 11169 44048 11203
rect 43996 11160 44048 11169
rect 44272 11135 44324 11144
rect 44272 11101 44281 11135
rect 44281 11101 44315 11135
rect 44315 11101 44324 11135
rect 44272 11092 44324 11101
rect 34612 11024 34664 11076
rect 35072 11024 35124 11076
rect 36544 10999 36596 11008
rect 36544 10965 36553 10999
rect 36553 10965 36587 10999
rect 36587 10965 36596 10999
rect 36544 10956 36596 10965
rect 37372 10999 37424 11008
rect 37372 10965 37381 10999
rect 37381 10965 37415 10999
rect 37415 10965 37424 10999
rect 37372 10956 37424 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 7472 10752 7524 10804
rect 12072 10752 12124 10804
rect 12164 10752 12216 10804
rect 12992 10752 13044 10804
rect 15384 10752 15436 10804
rect 16856 10752 16908 10804
rect 17224 10752 17276 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18328 10752 18380 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 21456 10752 21508 10804
rect 5724 10616 5776 10668
rect 7104 10616 7156 10668
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 4712 10548 4764 10600
rect 6736 10548 6788 10600
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 7472 10548 7524 10600
rect 11428 10616 11480 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 9588 10548 9640 10600
rect 10692 10480 10744 10532
rect 10784 10480 10836 10532
rect 11520 10480 11572 10532
rect 11796 10480 11848 10532
rect 11980 10480 12032 10532
rect 12072 10480 12124 10532
rect 4620 10412 4672 10464
rect 5632 10412 5684 10464
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 11888 10412 11940 10464
rect 12808 10684 12860 10736
rect 14188 10684 14240 10736
rect 14740 10684 14792 10736
rect 14832 10684 14884 10736
rect 12624 10616 12676 10668
rect 13084 10616 13136 10668
rect 13360 10616 13412 10668
rect 14740 10548 14792 10600
rect 16212 10616 16264 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17868 10616 17920 10668
rect 18236 10684 18288 10736
rect 19248 10727 19300 10736
rect 19248 10693 19257 10727
rect 19257 10693 19291 10727
rect 19291 10693 19300 10727
rect 19248 10684 19300 10693
rect 22100 10752 22152 10804
rect 22928 10752 22980 10804
rect 23112 10752 23164 10804
rect 24584 10752 24636 10804
rect 19064 10616 19116 10668
rect 16120 10548 16172 10600
rect 17500 10548 17552 10600
rect 17776 10591 17828 10600
rect 17776 10557 17785 10591
rect 17785 10557 17819 10591
rect 17819 10557 17828 10591
rect 17776 10548 17828 10557
rect 18328 10548 18380 10600
rect 19432 10548 19484 10600
rect 20720 10616 20772 10668
rect 22008 10727 22060 10736
rect 22008 10693 22017 10727
rect 22017 10693 22051 10727
rect 22051 10693 22060 10727
rect 22008 10684 22060 10693
rect 25872 10752 25924 10804
rect 27804 10752 27856 10804
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 21272 10548 21324 10600
rect 22100 10616 22152 10668
rect 21548 10548 21600 10600
rect 22284 10616 22336 10668
rect 22468 10480 22520 10532
rect 14096 10412 14148 10464
rect 17408 10412 17460 10464
rect 18052 10412 18104 10464
rect 19432 10412 19484 10464
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 23480 10616 23532 10668
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 25504 10659 25556 10668
rect 25504 10625 25513 10659
rect 25513 10625 25547 10659
rect 25547 10625 25556 10659
rect 25504 10616 25556 10625
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 27712 10616 27764 10668
rect 28632 10616 28684 10668
rect 29736 10752 29788 10804
rect 30288 10795 30340 10804
rect 30288 10761 30297 10795
rect 30297 10761 30331 10795
rect 30331 10761 30340 10795
rect 30288 10752 30340 10761
rect 30472 10752 30524 10804
rect 29000 10684 29052 10736
rect 24308 10523 24360 10532
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 25136 10548 25188 10600
rect 26332 10548 26384 10600
rect 27252 10548 27304 10600
rect 27436 10548 27488 10600
rect 28540 10548 28592 10600
rect 25044 10480 25096 10532
rect 29460 10727 29512 10736
rect 29460 10693 29469 10727
rect 29469 10693 29503 10727
rect 29503 10693 29512 10727
rect 29460 10684 29512 10693
rect 29552 10684 29604 10736
rect 31944 10752 31996 10804
rect 32220 10752 32272 10804
rect 34796 10752 34848 10804
rect 30748 10684 30800 10736
rect 31116 10684 31168 10736
rect 30380 10616 30432 10668
rect 30840 10659 30892 10668
rect 30840 10625 30849 10659
rect 30849 10625 30883 10659
rect 30883 10625 30892 10659
rect 30840 10616 30892 10625
rect 30012 10591 30064 10600
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 31668 10659 31720 10668
rect 31668 10625 31677 10659
rect 31677 10625 31711 10659
rect 31711 10625 31720 10659
rect 31668 10616 31720 10625
rect 31944 10659 31996 10668
rect 31944 10625 31953 10659
rect 31953 10625 31987 10659
rect 31987 10625 31996 10659
rect 31944 10616 31996 10625
rect 33784 10727 33836 10736
rect 33784 10693 33793 10727
rect 33793 10693 33827 10727
rect 33827 10693 33836 10727
rect 33784 10684 33836 10693
rect 35256 10795 35308 10804
rect 35256 10761 35265 10795
rect 35265 10761 35299 10795
rect 35299 10761 35308 10795
rect 35256 10752 35308 10761
rect 36268 10752 36320 10804
rect 37280 10752 37332 10804
rect 37372 10752 37424 10804
rect 39488 10752 39540 10804
rect 36544 10684 36596 10736
rect 37648 10684 37700 10736
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 32956 10616 33008 10668
rect 35072 10616 35124 10668
rect 35532 10616 35584 10668
rect 36084 10616 36136 10668
rect 37280 10659 37332 10668
rect 37280 10625 37289 10659
rect 37289 10625 37323 10659
rect 37323 10625 37332 10659
rect 37280 10616 37332 10625
rect 31484 10591 31536 10600
rect 31484 10557 31493 10591
rect 31493 10557 31527 10591
rect 31527 10557 31536 10591
rect 31484 10548 31536 10557
rect 32036 10548 32088 10600
rect 31208 10480 31260 10532
rect 28264 10455 28316 10464
rect 28264 10421 28273 10455
rect 28273 10421 28307 10455
rect 28307 10421 28316 10455
rect 28264 10412 28316 10421
rect 30472 10412 30524 10464
rect 30748 10412 30800 10464
rect 30840 10412 30892 10464
rect 31944 10480 31996 10532
rect 33508 10591 33560 10600
rect 33508 10557 33517 10591
rect 33517 10557 33551 10591
rect 33551 10557 33560 10591
rect 33508 10548 33560 10557
rect 36912 10591 36964 10600
rect 36912 10557 36921 10591
rect 36921 10557 36955 10591
rect 36955 10557 36964 10591
rect 36912 10548 36964 10557
rect 37188 10480 37240 10532
rect 38568 10480 38620 10532
rect 41420 10548 41472 10600
rect 32864 10455 32916 10464
rect 32864 10421 32873 10455
rect 32873 10421 32907 10455
rect 32907 10421 32916 10455
rect 32864 10412 32916 10421
rect 36176 10412 36228 10464
rect 37372 10412 37424 10464
rect 39028 10412 39080 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4712 10208 4764 10260
rect 10968 10251 11020 10260
rect 10048 10072 10100 10124
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 9864 10004 9916 10056
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 17960 10208 18012 10260
rect 21916 10208 21968 10260
rect 11796 10140 11848 10192
rect 12624 10140 12676 10192
rect 12072 10072 12124 10124
rect 13268 10072 13320 10124
rect 10784 10004 10836 10056
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11336 10004 11388 10056
rect 11520 10004 11572 10056
rect 14740 10004 14792 10056
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 18788 10140 18840 10192
rect 18236 10072 18288 10124
rect 22284 10208 22336 10260
rect 27804 10208 27856 10260
rect 22192 10140 22244 10192
rect 22468 10140 22520 10192
rect 22744 10140 22796 10192
rect 10692 9936 10744 9988
rect 15476 9936 15528 9988
rect 15844 10004 15896 10056
rect 15660 9936 15712 9988
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 19156 10004 19208 10056
rect 19800 10004 19852 10056
rect 19984 10004 20036 10056
rect 22100 10004 22152 10056
rect 22928 10004 22980 10056
rect 28264 10208 28316 10260
rect 28632 10208 28684 10260
rect 29276 10208 29328 10260
rect 29828 10208 29880 10260
rect 31024 10208 31076 10260
rect 31852 10208 31904 10260
rect 37280 10208 37332 10260
rect 38108 10208 38160 10260
rect 29736 10140 29788 10192
rect 28540 10072 28592 10124
rect 29276 10072 29328 10124
rect 31208 10072 31260 10124
rect 39028 10072 39080 10124
rect 28448 10004 28500 10056
rect 18788 9936 18840 9988
rect 10324 9868 10376 9920
rect 11428 9868 11480 9920
rect 16672 9868 16724 9920
rect 21916 9936 21968 9988
rect 22376 9979 22428 9988
rect 22376 9945 22385 9979
rect 22385 9945 22419 9979
rect 22419 9945 22428 9979
rect 22376 9936 22428 9945
rect 22468 9936 22520 9988
rect 28632 10047 28684 10056
rect 28632 10013 28641 10047
rect 28641 10013 28675 10047
rect 28675 10013 28684 10047
rect 28632 10004 28684 10013
rect 28908 10047 28960 10056
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10004 28960 10013
rect 30472 10004 30524 10056
rect 31760 10004 31812 10056
rect 37648 10004 37700 10056
rect 40868 9936 40920 9988
rect 19800 9868 19852 9920
rect 20628 9868 20680 9920
rect 22008 9868 22060 9920
rect 22928 9868 22980 9920
rect 26976 9868 27028 9920
rect 30748 9868 30800 9920
rect 31576 9868 31628 9920
rect 31760 9868 31812 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 5172 9664 5224 9716
rect 10232 9664 10284 9716
rect 10784 9664 10836 9716
rect 4804 9596 4856 9648
rect 5724 9596 5776 9648
rect 11152 9596 11204 9648
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 10324 9571 10376 9580
rect 10324 9537 10342 9571
rect 10342 9537 10376 9571
rect 10324 9528 10376 9537
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 4620 9392 4672 9444
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 11244 9460 11296 9512
rect 10968 9392 11020 9444
rect 12256 9528 12308 9580
rect 13268 9528 13320 9580
rect 13728 9596 13780 9648
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 14004 9596 14056 9648
rect 14188 9596 14240 9648
rect 14648 9596 14700 9648
rect 18328 9664 18380 9716
rect 20168 9664 20220 9716
rect 21272 9664 21324 9716
rect 14372 9528 14424 9580
rect 18052 9596 18104 9648
rect 21548 9596 21600 9648
rect 21916 9664 21968 9716
rect 23940 9664 23992 9716
rect 24676 9664 24728 9716
rect 27344 9664 27396 9716
rect 28908 9664 28960 9716
rect 31392 9664 31444 9716
rect 40868 9707 40920 9716
rect 40868 9673 40877 9707
rect 40877 9673 40911 9707
rect 40911 9673 40920 9707
rect 40868 9664 40920 9673
rect 16580 9528 16632 9580
rect 16672 9528 16724 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17408 9528 17460 9580
rect 17592 9528 17644 9580
rect 18604 9528 18656 9580
rect 18972 9528 19024 9580
rect 20352 9528 20404 9580
rect 23388 9596 23440 9648
rect 21916 9528 21968 9580
rect 22008 9528 22060 9580
rect 32864 9596 32916 9648
rect 42524 9639 42576 9648
rect 42524 9605 42533 9639
rect 42533 9605 42567 9639
rect 42567 9605 42576 9639
rect 42524 9596 42576 9605
rect 15844 9460 15896 9512
rect 14096 9392 14148 9444
rect 16304 9503 16356 9512
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 16488 9460 16540 9512
rect 20536 9460 20588 9512
rect 20720 9460 20772 9512
rect 21456 9460 21508 9512
rect 23664 9503 23716 9512
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 14188 9324 14240 9376
rect 22100 9392 22152 9444
rect 22652 9392 22704 9444
rect 22836 9392 22888 9444
rect 25228 9460 25280 9512
rect 26608 9460 26660 9512
rect 28540 9503 28592 9512
rect 28540 9469 28549 9503
rect 28549 9469 28583 9503
rect 28583 9469 28592 9503
rect 28540 9460 28592 9469
rect 28908 9571 28960 9580
rect 28908 9537 28917 9571
rect 28917 9537 28951 9571
rect 28951 9537 28960 9571
rect 28908 9528 28960 9537
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 29552 9528 29604 9580
rect 30656 9571 30708 9580
rect 30656 9537 30665 9571
rect 30665 9537 30699 9571
rect 30699 9537 30708 9571
rect 30656 9528 30708 9537
rect 30840 9571 30892 9580
rect 30840 9537 30849 9571
rect 30849 9537 30883 9571
rect 30883 9537 30892 9571
rect 30840 9528 30892 9537
rect 32036 9528 32088 9580
rect 27344 9392 27396 9444
rect 30012 9460 30064 9512
rect 31668 9503 31720 9512
rect 31668 9469 31677 9503
rect 31677 9469 31711 9503
rect 31711 9469 31720 9503
rect 31668 9460 31720 9469
rect 31760 9503 31812 9512
rect 31760 9469 31769 9503
rect 31769 9469 31803 9503
rect 31803 9469 31812 9503
rect 31760 9460 31812 9469
rect 21732 9324 21784 9376
rect 24400 9324 24452 9376
rect 24768 9324 24820 9376
rect 24860 9324 24912 9376
rect 25504 9324 25556 9376
rect 26148 9324 26200 9376
rect 28448 9367 28500 9376
rect 28448 9333 28457 9367
rect 28457 9333 28491 9367
rect 28491 9333 28500 9367
rect 28448 9324 28500 9333
rect 28816 9324 28868 9376
rect 30472 9392 30524 9444
rect 32220 9528 32272 9580
rect 33968 9435 34020 9444
rect 33968 9401 33977 9435
rect 33977 9401 34011 9435
rect 34011 9401 34020 9435
rect 33968 9392 34020 9401
rect 38568 9460 38620 9512
rect 41512 9503 41564 9512
rect 41512 9469 41521 9503
rect 41521 9469 41555 9503
rect 41555 9469 41564 9503
rect 41512 9460 41564 9469
rect 29644 9324 29696 9376
rect 30840 9324 30892 9376
rect 31208 9324 31260 9376
rect 31576 9324 31628 9376
rect 31760 9324 31812 9376
rect 31944 9324 31996 9376
rect 34060 9324 34112 9376
rect 34152 9367 34204 9376
rect 34152 9333 34161 9367
rect 34161 9333 34195 9367
rect 34195 9333 34204 9367
rect 34152 9324 34204 9333
rect 43720 9324 43772 9376
rect 44272 9324 44324 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2504 9120 2556 9172
rect 10416 9120 10468 9172
rect 10600 9120 10652 9172
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 11980 9120 12032 9172
rect 12532 9120 12584 9172
rect 12716 9120 12768 9172
rect 13636 9120 13688 9172
rect 14004 9120 14056 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 940 8916 992 8968
rect 9680 9052 9732 9104
rect 10048 9052 10100 9104
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 7380 8984 7432 9036
rect 7104 8848 7156 8900
rect 10508 8984 10560 9036
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 13176 9052 13228 9104
rect 14372 9120 14424 9172
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 9772 8891 9824 8900
rect 9772 8857 9781 8891
rect 9781 8857 9815 8891
rect 9815 8857 9824 8891
rect 9772 8848 9824 8857
rect 10416 8848 10468 8900
rect 10508 8891 10560 8900
rect 10508 8857 10517 8891
rect 10517 8857 10551 8891
rect 10551 8857 10560 8891
rect 10508 8848 10560 8857
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 16304 9120 16356 9172
rect 17132 9120 17184 9172
rect 17408 9120 17460 9172
rect 15568 9052 15620 9104
rect 17224 9052 17276 9104
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 12072 8780 12124 8832
rect 13360 8916 13412 8968
rect 13636 8916 13688 8968
rect 14188 8916 14240 8968
rect 14372 8916 14424 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 13268 8848 13320 8900
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14924 8916 14976 8968
rect 16028 8916 16080 8968
rect 16580 8984 16632 9036
rect 17592 9052 17644 9104
rect 17960 9095 18012 9104
rect 17960 9061 17969 9095
rect 17969 9061 18003 9095
rect 18003 9061 18012 9095
rect 17960 9052 18012 9061
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 14004 8780 14056 8832
rect 16948 8848 17000 8900
rect 17224 8959 17276 8968
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 17592 8916 17644 8968
rect 17316 8848 17368 8900
rect 18696 9120 18748 9172
rect 19340 9120 19392 9172
rect 19984 9120 20036 9172
rect 20168 9120 20220 9172
rect 20536 9120 20588 9172
rect 22284 9120 22336 9172
rect 22376 9120 22428 9172
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 24676 9120 24728 9172
rect 27804 9120 27856 9172
rect 30656 9120 30708 9172
rect 31484 9163 31536 9172
rect 31484 9129 31493 9163
rect 31493 9129 31527 9163
rect 31527 9129 31536 9163
rect 31484 9120 31536 9129
rect 36912 9120 36964 9172
rect 18236 9052 18288 9104
rect 18236 8916 18288 8968
rect 18788 9052 18840 9104
rect 22008 9052 22060 9104
rect 22468 9052 22520 9104
rect 22652 9052 22704 9104
rect 24768 9052 24820 9104
rect 17408 8780 17460 8832
rect 17592 8780 17644 8832
rect 18328 8780 18380 8832
rect 18604 8780 18656 8832
rect 19340 8848 19392 8900
rect 19984 8916 20036 8968
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 20628 8916 20680 8968
rect 21732 8959 21784 8968
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 23020 8984 23072 9036
rect 23480 8984 23532 9036
rect 30472 9052 30524 9104
rect 25228 8984 25280 9036
rect 26608 8984 26660 9036
rect 26976 9027 27028 9036
rect 26976 8993 26985 9027
rect 26985 8993 27019 9027
rect 27019 8993 27028 9027
rect 26976 8984 27028 8993
rect 27252 8984 27304 9036
rect 29736 8984 29788 9036
rect 31024 9052 31076 9104
rect 31576 9052 31628 9104
rect 26148 8959 26200 8968
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 27712 8916 27764 8968
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 29276 8916 29328 8968
rect 30380 8916 30432 8968
rect 31208 8984 31260 9036
rect 33140 8984 33192 9036
rect 33508 8984 33560 9036
rect 35348 8984 35400 9036
rect 31668 8916 31720 8968
rect 24952 8848 25004 8900
rect 28172 8891 28224 8900
rect 28172 8857 28181 8891
rect 28181 8857 28215 8891
rect 28215 8857 28224 8891
rect 28172 8848 28224 8857
rect 29184 8848 29236 8900
rect 30472 8848 30524 8900
rect 30656 8891 30708 8900
rect 30656 8857 30665 8891
rect 30665 8857 30699 8891
rect 30699 8857 30708 8891
rect 30656 8848 30708 8857
rect 20168 8780 20220 8832
rect 22652 8780 22704 8832
rect 23480 8780 23532 8832
rect 25872 8780 25924 8832
rect 26332 8780 26384 8832
rect 26884 8823 26936 8832
rect 26884 8789 26893 8823
rect 26893 8789 26927 8823
rect 26927 8789 26936 8823
rect 26884 8780 26936 8789
rect 29644 8780 29696 8832
rect 31116 8780 31168 8832
rect 34796 8848 34848 8900
rect 34520 8823 34572 8832
rect 34520 8789 34529 8823
rect 34529 8789 34563 8823
rect 34563 8789 34572 8823
rect 34520 8780 34572 8789
rect 35440 8848 35492 8900
rect 36084 8780 36136 8832
rect 37924 8916 37976 8968
rect 37740 8823 37792 8832
rect 37740 8789 37749 8823
rect 37749 8789 37783 8823
rect 37783 8789 37792 8823
rect 37740 8780 37792 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 10140 8576 10192 8628
rect 10232 8576 10284 8628
rect 11520 8576 11572 8628
rect 12164 8576 12216 8628
rect 12900 8576 12952 8628
rect 13176 8576 13228 8628
rect 14464 8576 14516 8628
rect 14556 8576 14608 8628
rect 17040 8576 17092 8628
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 17592 8576 17644 8628
rect 17960 8576 18012 8628
rect 7932 8440 7984 8492
rect 7380 8372 7432 8424
rect 8300 8372 8352 8424
rect 10324 8508 10376 8560
rect 14004 8508 14056 8560
rect 10140 8440 10192 8492
rect 10508 8440 10560 8492
rect 11888 8440 11940 8492
rect 11980 8440 12032 8492
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 13176 8440 13228 8492
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 13728 8440 13780 8492
rect 13912 8440 13964 8492
rect 11704 8372 11756 8424
rect 15660 8440 15712 8492
rect 16028 8440 16080 8492
rect 17500 8508 17552 8560
rect 18144 8508 18196 8560
rect 18328 8508 18380 8560
rect 17316 8440 17368 8492
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 18052 8372 18104 8424
rect 18328 8415 18380 8424
rect 18328 8381 18337 8415
rect 18337 8381 18371 8415
rect 18371 8381 18380 8415
rect 18328 8372 18380 8381
rect 18880 8372 18932 8424
rect 12532 8304 12584 8356
rect 13636 8304 13688 8356
rect 17224 8304 17276 8356
rect 18788 8304 18840 8356
rect 9956 8236 10008 8288
rect 11428 8236 11480 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 12072 8236 12124 8288
rect 13360 8236 13412 8288
rect 13452 8236 13504 8288
rect 17592 8236 17644 8288
rect 18236 8236 18288 8288
rect 20352 8576 20404 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 22008 8576 22060 8628
rect 23388 8576 23440 8628
rect 23664 8576 23716 8628
rect 24952 8576 25004 8628
rect 26884 8576 26936 8628
rect 28540 8576 28592 8628
rect 29736 8576 29788 8628
rect 30656 8576 30708 8628
rect 22468 8508 22520 8560
rect 21916 8483 21968 8492
rect 21916 8449 21925 8483
rect 21925 8449 21959 8483
rect 21959 8449 21968 8483
rect 21916 8440 21968 8449
rect 23480 8440 23532 8492
rect 21364 8415 21416 8424
rect 21364 8381 21373 8415
rect 21373 8381 21407 8415
rect 21407 8381 21416 8415
rect 21364 8372 21416 8381
rect 22192 8372 22244 8424
rect 22284 8304 22336 8356
rect 19524 8236 19576 8288
rect 20168 8236 20220 8288
rect 22100 8279 22152 8288
rect 22100 8245 22109 8279
rect 22109 8245 22143 8279
rect 22143 8245 22152 8279
rect 22100 8236 22152 8245
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 24032 8440 24084 8492
rect 28632 8508 28684 8560
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 25320 8372 25372 8424
rect 24952 8304 25004 8356
rect 26608 8372 26660 8424
rect 27068 8372 27120 8424
rect 28172 8372 28224 8424
rect 29552 8440 29604 8492
rect 30196 8440 30248 8492
rect 30380 8440 30432 8492
rect 30932 8508 30984 8560
rect 32220 8576 32272 8628
rect 34152 8576 34204 8628
rect 34520 8576 34572 8628
rect 35440 8576 35492 8628
rect 37740 8576 37792 8628
rect 41512 8576 41564 8628
rect 26332 8304 26384 8356
rect 29184 8372 29236 8424
rect 31208 8440 31260 8492
rect 31300 8440 31352 8492
rect 31944 8440 31996 8492
rect 43720 8508 43772 8560
rect 27160 8304 27212 8356
rect 28816 8304 28868 8356
rect 24584 8236 24636 8288
rect 25688 8279 25740 8288
rect 25688 8245 25697 8279
rect 25697 8245 25731 8279
rect 25731 8245 25740 8279
rect 25688 8236 25740 8245
rect 30840 8415 30892 8424
rect 30840 8381 30849 8415
rect 30849 8381 30883 8415
rect 30883 8381 30892 8415
rect 30840 8372 30892 8381
rect 31116 8372 31168 8424
rect 35532 8372 35584 8424
rect 36084 8483 36136 8492
rect 36084 8449 36093 8483
rect 36093 8449 36127 8483
rect 36127 8449 36136 8483
rect 36084 8440 36136 8449
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 38384 8440 38436 8492
rect 31484 8304 31536 8356
rect 33232 8304 33284 8356
rect 34060 8347 34112 8356
rect 34060 8313 34069 8347
rect 34069 8313 34103 8347
rect 34103 8313 34112 8347
rect 34060 8304 34112 8313
rect 34336 8304 34388 8356
rect 42800 8372 42852 8424
rect 43996 8415 44048 8424
rect 43996 8381 44005 8415
rect 44005 8381 44039 8415
rect 44039 8381 44048 8415
rect 43996 8372 44048 8381
rect 31392 8236 31444 8288
rect 31576 8279 31628 8288
rect 31576 8245 31585 8279
rect 31585 8245 31619 8279
rect 31619 8245 31628 8279
rect 31576 8236 31628 8245
rect 31944 8236 31996 8288
rect 36176 8279 36228 8288
rect 36176 8245 36185 8279
rect 36185 8245 36219 8279
rect 36219 8245 36228 8279
rect 36176 8236 36228 8245
rect 37924 8236 37976 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 6736 8032 6788 8084
rect 12256 8032 12308 8084
rect 11060 7964 11112 8016
rect 13268 8032 13320 8084
rect 13452 8032 13504 8084
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7196 7828 7248 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10692 7828 10744 7880
rect 11060 7828 11112 7880
rect 15660 7964 15712 8016
rect 16396 8032 16448 8084
rect 18236 8032 18288 8084
rect 18328 8032 18380 8084
rect 18880 8032 18932 8084
rect 19984 8032 20036 8084
rect 20628 8032 20680 8084
rect 21548 8032 21600 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 23480 8075 23532 8084
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 25872 8075 25924 8084
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 27712 8032 27764 8084
rect 28264 8075 28316 8084
rect 28264 8041 28273 8075
rect 28273 8041 28307 8075
rect 28307 8041 28316 8075
rect 28264 8032 28316 8041
rect 28816 8032 28868 8084
rect 11888 7896 11940 7948
rect 11428 7828 11480 7880
rect 12900 7828 12952 7880
rect 14924 7828 14976 7880
rect 15016 7828 15068 7880
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 17684 7896 17736 7948
rect 13084 7803 13136 7812
rect 13084 7769 13093 7803
rect 13093 7769 13127 7803
rect 13127 7769 13136 7803
rect 13084 7760 13136 7769
rect 13544 7760 13596 7812
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 15292 7760 15344 7812
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 15200 7692 15252 7744
rect 16488 7828 16540 7880
rect 17040 7828 17092 7880
rect 17592 7828 17644 7880
rect 18604 7896 18656 7948
rect 19984 7896 20036 7948
rect 20260 7896 20312 7948
rect 21916 7939 21968 7948
rect 21916 7905 21925 7939
rect 21925 7905 21959 7939
rect 21959 7905 21968 7939
rect 21916 7896 21968 7905
rect 15660 7692 15712 7744
rect 17040 7735 17092 7744
rect 17040 7701 17049 7735
rect 17049 7701 17083 7735
rect 17083 7701 17092 7735
rect 17040 7692 17092 7701
rect 17684 7692 17736 7744
rect 21824 7828 21876 7880
rect 30196 8007 30248 8016
rect 30196 7973 30205 8007
rect 30205 7973 30239 8007
rect 30239 7973 30248 8007
rect 30196 7964 30248 7973
rect 30840 7964 30892 8016
rect 31300 8032 31352 8084
rect 31576 8075 31628 8084
rect 31576 8041 31585 8075
rect 31585 8041 31619 8075
rect 31619 8041 31628 8075
rect 31576 8032 31628 8041
rect 38016 8032 38068 8084
rect 38384 8075 38436 8084
rect 38384 8041 38393 8075
rect 38393 8041 38427 8075
rect 38427 8041 38436 8075
rect 38384 8032 38436 8041
rect 43996 8032 44048 8084
rect 22192 7896 22244 7948
rect 24584 7896 24636 7948
rect 24676 7896 24728 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 27436 7896 27488 7948
rect 28908 7896 28960 7948
rect 29184 7896 29236 7948
rect 37924 7964 37976 8016
rect 37280 7896 37332 7948
rect 25688 7828 25740 7880
rect 22100 7760 22152 7812
rect 22652 7803 22704 7812
rect 22652 7769 22661 7803
rect 22661 7769 22695 7803
rect 22695 7769 22704 7803
rect 22652 7760 22704 7769
rect 18512 7692 18564 7744
rect 22744 7735 22796 7744
rect 22744 7701 22753 7735
rect 22753 7701 22787 7735
rect 22787 7701 22796 7735
rect 22744 7692 22796 7701
rect 24308 7692 24360 7744
rect 24860 7803 24912 7812
rect 24860 7769 24869 7803
rect 24869 7769 24903 7803
rect 24903 7769 24912 7803
rect 24860 7760 24912 7769
rect 29276 7828 29328 7880
rect 29828 7828 29880 7880
rect 30104 7828 30156 7880
rect 30196 7828 30248 7880
rect 31484 7828 31536 7880
rect 28448 7803 28500 7812
rect 28448 7769 28457 7803
rect 28457 7769 28491 7803
rect 28491 7769 28500 7803
rect 28448 7760 28500 7769
rect 29920 7760 29972 7812
rect 27528 7692 27580 7744
rect 27712 7692 27764 7744
rect 28632 7692 28684 7744
rect 29828 7692 29880 7744
rect 31760 7760 31812 7812
rect 33784 7760 33836 7812
rect 34336 7760 34388 7812
rect 35900 7760 35952 7812
rect 43352 7871 43404 7880
rect 43352 7837 43361 7871
rect 43361 7837 43395 7871
rect 43395 7837 43404 7871
rect 43352 7828 43404 7837
rect 38568 7803 38620 7812
rect 38568 7769 38577 7803
rect 38577 7769 38611 7803
rect 38611 7769 38620 7803
rect 38568 7760 38620 7769
rect 33416 7692 33468 7744
rect 35348 7692 35400 7744
rect 37004 7692 37056 7744
rect 37372 7692 37424 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 7196 7488 7248 7540
rect 7748 7488 7800 7540
rect 9956 7488 10008 7540
rect 7288 7352 7340 7404
rect 10048 7420 10100 7472
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 11428 7488 11480 7540
rect 12440 7488 12492 7540
rect 13360 7488 13412 7540
rect 15384 7488 15436 7540
rect 15936 7488 15988 7540
rect 19340 7488 19392 7540
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 21824 7488 21876 7540
rect 22744 7488 22796 7540
rect 24952 7488 25004 7540
rect 11612 7420 11664 7472
rect 18144 7420 18196 7472
rect 22468 7420 22520 7472
rect 25044 7420 25096 7472
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 26700 7488 26752 7540
rect 26976 7488 27028 7540
rect 27896 7488 27948 7540
rect 28264 7488 28316 7540
rect 28908 7488 28960 7540
rect 29276 7488 29328 7540
rect 6736 7284 6788 7336
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 7472 7284 7524 7293
rect 8208 7216 8260 7268
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 10876 7352 10928 7404
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 12348 7352 12400 7404
rect 14188 7352 14240 7404
rect 10508 7216 10560 7268
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12900 7284 12952 7336
rect 11060 7216 11112 7268
rect 11796 7216 11848 7268
rect 13176 7216 13228 7268
rect 13636 7216 13688 7268
rect 17960 7352 18012 7404
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 18788 7352 18840 7404
rect 20812 7352 20864 7404
rect 14924 7284 14976 7336
rect 14648 7216 14700 7268
rect 16028 7284 16080 7336
rect 22836 7395 22888 7404
rect 22836 7361 22844 7395
rect 22844 7361 22878 7395
rect 22878 7361 22888 7395
rect 22836 7352 22888 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 24676 7352 24728 7404
rect 25688 7395 25740 7404
rect 25688 7361 25697 7395
rect 25697 7361 25731 7395
rect 25731 7361 25740 7395
rect 25688 7352 25740 7361
rect 27160 7420 27212 7472
rect 26516 7395 26568 7404
rect 26516 7361 26525 7395
rect 26525 7361 26559 7395
rect 26559 7361 26568 7395
rect 26516 7352 26568 7361
rect 21456 7284 21508 7336
rect 22192 7259 22244 7268
rect 22192 7225 22201 7259
rect 22201 7225 22235 7259
rect 22235 7225 22244 7259
rect 22192 7216 22244 7225
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 25872 7327 25924 7336
rect 25872 7293 25881 7327
rect 25881 7293 25915 7327
rect 25915 7293 25924 7327
rect 25872 7284 25924 7293
rect 26792 7395 26844 7404
rect 26792 7361 26801 7395
rect 26801 7361 26835 7395
rect 26835 7361 26844 7395
rect 26792 7352 26844 7361
rect 27712 7352 27764 7404
rect 28724 7420 28776 7472
rect 30104 7488 30156 7540
rect 29460 7420 29512 7472
rect 30196 7420 30248 7472
rect 33140 7531 33192 7540
rect 33140 7497 33149 7531
rect 33149 7497 33183 7531
rect 33183 7497 33192 7531
rect 33140 7488 33192 7497
rect 33784 7488 33836 7540
rect 35992 7488 36044 7540
rect 31760 7420 31812 7472
rect 31852 7420 31904 7472
rect 35900 7420 35952 7472
rect 37372 7488 37424 7540
rect 37464 7531 37516 7540
rect 37464 7497 37473 7531
rect 37473 7497 37507 7531
rect 37507 7497 37516 7531
rect 37464 7488 37516 7497
rect 38568 7488 38620 7540
rect 27436 7284 27488 7336
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 10692 7148 10744 7200
rect 11428 7148 11480 7200
rect 19340 7148 19392 7200
rect 23480 7148 23532 7200
rect 25320 7148 25372 7200
rect 25596 7148 25648 7200
rect 25872 7148 25924 7200
rect 29000 7216 29052 7268
rect 29644 7352 29696 7404
rect 29920 7395 29972 7404
rect 29920 7361 29930 7395
rect 29930 7361 29964 7395
rect 29964 7361 29972 7395
rect 29920 7352 29972 7361
rect 31024 7352 31076 7404
rect 29460 7284 29512 7336
rect 29184 7216 29236 7268
rect 29552 7259 29604 7268
rect 29552 7225 29561 7259
rect 29561 7225 29595 7259
rect 29595 7225 29604 7259
rect 29552 7216 29604 7225
rect 29828 7327 29880 7336
rect 29828 7293 29837 7327
rect 29837 7293 29871 7327
rect 29871 7293 29880 7327
rect 29828 7284 29880 7293
rect 30748 7284 30800 7336
rect 31116 7284 31168 7336
rect 31576 7284 31628 7336
rect 35348 7327 35400 7336
rect 35348 7293 35357 7327
rect 35357 7293 35391 7327
rect 35391 7293 35400 7327
rect 35348 7284 35400 7293
rect 36176 7284 36228 7336
rect 38476 7420 38528 7472
rect 42800 7488 42852 7540
rect 43352 7531 43404 7540
rect 43352 7497 43361 7531
rect 43361 7497 43395 7531
rect 43395 7497 43404 7531
rect 43352 7488 43404 7497
rect 43812 7463 43864 7472
rect 43812 7429 43821 7463
rect 43821 7429 43855 7463
rect 43855 7429 43864 7463
rect 43812 7420 43864 7429
rect 43720 7352 43772 7404
rect 44088 7352 44140 7404
rect 38476 7284 38528 7336
rect 38936 7327 38988 7336
rect 38936 7293 38945 7327
rect 38945 7293 38979 7327
rect 38979 7293 38988 7327
rect 38936 7284 38988 7293
rect 30104 7216 30156 7268
rect 27068 7148 27120 7200
rect 29092 7148 29144 7200
rect 30472 7148 30524 7200
rect 30564 7191 30616 7200
rect 30564 7157 30573 7191
rect 30573 7157 30607 7191
rect 30607 7157 30616 7191
rect 30564 7148 30616 7157
rect 30840 7148 30892 7200
rect 31484 7148 31536 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10876 6944 10928 6996
rect 11244 6944 11296 6996
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2044 6808 2096 6860
rect 7472 6808 7524 6860
rect 13820 6944 13872 6996
rect 14924 6987 14976 6996
rect 14924 6953 14933 6987
rect 14933 6953 14967 6987
rect 14967 6953 14976 6987
rect 14924 6944 14976 6953
rect 12532 6876 12584 6928
rect 15016 6876 15068 6928
rect 7104 6740 7156 6792
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 10232 6740 10284 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 10968 6740 11020 6792
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 7288 6672 7340 6724
rect 9772 6672 9824 6724
rect 10692 6672 10744 6724
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11704 6740 11756 6792
rect 11888 6672 11940 6724
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 7656 6604 7708 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 11244 6604 11296 6656
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 12532 6672 12584 6724
rect 14004 6672 14056 6724
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 15200 6740 15252 6792
rect 15936 6740 15988 6792
rect 16028 6740 16080 6792
rect 16396 6740 16448 6792
rect 25044 6987 25096 6996
rect 25044 6953 25053 6987
rect 25053 6953 25087 6987
rect 25087 6953 25096 6987
rect 25044 6944 25096 6953
rect 26700 6944 26752 6996
rect 18880 6876 18932 6928
rect 20076 6876 20128 6928
rect 27712 6944 27764 6996
rect 30380 6944 30432 6996
rect 30564 6944 30616 6996
rect 19248 6808 19300 6860
rect 23480 6808 23532 6860
rect 24584 6808 24636 6860
rect 25596 6851 25648 6860
rect 25596 6817 25605 6851
rect 25605 6817 25639 6851
rect 25639 6817 25648 6851
rect 25596 6808 25648 6817
rect 26700 6851 26752 6860
rect 26700 6817 26718 6851
rect 26718 6817 26752 6851
rect 26700 6808 26752 6817
rect 27068 6851 27120 6860
rect 27068 6817 27077 6851
rect 27077 6817 27111 6851
rect 27111 6817 27120 6851
rect 27068 6808 27120 6817
rect 27160 6808 27212 6860
rect 27528 6851 27580 6860
rect 27528 6817 27537 6851
rect 27537 6817 27571 6851
rect 27571 6817 27580 6851
rect 27528 6808 27580 6817
rect 18236 6740 18288 6792
rect 17960 6672 18012 6724
rect 12716 6604 12768 6656
rect 13084 6604 13136 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 15292 6604 15344 6656
rect 15844 6604 15896 6656
rect 15936 6604 15988 6656
rect 17224 6604 17276 6656
rect 18052 6604 18104 6656
rect 18328 6715 18380 6724
rect 18328 6681 18337 6715
rect 18337 6681 18371 6715
rect 18371 6681 18380 6715
rect 18328 6672 18380 6681
rect 18604 6604 18656 6656
rect 25688 6604 25740 6656
rect 27804 6740 27856 6792
rect 27896 6740 27948 6792
rect 28816 6808 28868 6860
rect 28448 6740 28500 6792
rect 28908 6783 28960 6792
rect 28908 6749 28917 6783
rect 28917 6749 28951 6783
rect 28951 6749 28960 6783
rect 28908 6740 28960 6749
rect 29000 6783 29052 6792
rect 29000 6749 29009 6783
rect 29009 6749 29043 6783
rect 29043 6749 29052 6783
rect 29000 6740 29052 6749
rect 29460 6672 29512 6724
rect 29552 6672 29604 6724
rect 30104 6783 30156 6792
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30104 6740 30156 6749
rect 30840 6919 30892 6928
rect 30840 6885 30849 6919
rect 30849 6885 30883 6919
rect 30883 6885 30892 6919
rect 30840 6876 30892 6885
rect 31024 6944 31076 6996
rect 34336 6876 34388 6928
rect 30748 6740 30800 6792
rect 31116 6740 31168 6792
rect 31484 6783 31536 6792
rect 31484 6749 31493 6783
rect 31493 6749 31527 6783
rect 31527 6749 31536 6783
rect 31484 6740 31536 6749
rect 33416 6851 33468 6860
rect 33416 6817 33425 6851
rect 33425 6817 33459 6851
rect 33459 6817 33468 6851
rect 33416 6808 33468 6817
rect 35256 6944 35308 6996
rect 36084 6740 36136 6792
rect 37464 6851 37516 6860
rect 37464 6817 37473 6851
rect 37473 6817 37507 6851
rect 37507 6817 37516 6851
rect 37464 6808 37516 6817
rect 38200 6808 38252 6860
rect 37280 6783 37332 6792
rect 37280 6749 37289 6783
rect 37289 6749 37323 6783
rect 37323 6749 37332 6783
rect 37280 6740 37332 6749
rect 30840 6604 30892 6656
rect 35072 6715 35124 6724
rect 35072 6681 35081 6715
rect 35081 6681 35115 6715
rect 35115 6681 35124 6715
rect 35072 6672 35124 6681
rect 31300 6647 31352 6656
rect 31300 6613 31309 6647
rect 31309 6613 31343 6647
rect 31343 6613 31352 6647
rect 31300 6604 31352 6613
rect 32864 6604 32916 6656
rect 37004 6604 37056 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 3148 6400 3200 6452
rect 4804 6332 4856 6384
rect 8208 6332 8260 6384
rect 9864 6264 9916 6316
rect 11152 6264 11204 6316
rect 11244 6264 11296 6316
rect 11336 6264 11388 6316
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 10232 6196 10284 6248
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 12624 6400 12676 6452
rect 14556 6400 14608 6452
rect 14924 6443 14976 6452
rect 14924 6409 14933 6443
rect 14933 6409 14967 6443
rect 14967 6409 14976 6443
rect 14924 6400 14976 6409
rect 12164 6332 12216 6384
rect 12256 6307 12308 6316
rect 12256 6273 12265 6307
rect 12265 6273 12299 6307
rect 12299 6273 12308 6307
rect 12256 6264 12308 6273
rect 13636 6332 13688 6384
rect 14004 6332 14056 6384
rect 14188 6332 14240 6384
rect 15384 6400 15436 6452
rect 16672 6400 16724 6452
rect 14648 6264 14700 6316
rect 12992 6196 13044 6248
rect 15108 6264 15160 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 13636 6128 13688 6180
rect 8116 6060 8168 6112
rect 11152 6060 11204 6112
rect 12624 6060 12676 6112
rect 13360 6060 13412 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 13728 6060 13780 6112
rect 14832 6128 14884 6180
rect 14924 6128 14976 6180
rect 15936 6196 15988 6248
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17776 6400 17828 6452
rect 21916 6400 21968 6452
rect 22468 6443 22520 6452
rect 22468 6409 22477 6443
rect 22477 6409 22511 6443
rect 22511 6409 22520 6443
rect 22468 6400 22520 6409
rect 25688 6400 25740 6452
rect 27804 6400 27856 6452
rect 28816 6400 28868 6452
rect 35072 6400 35124 6452
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 17408 6264 17460 6316
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 17960 6264 18012 6316
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 27436 6375 27488 6384
rect 27436 6341 27445 6375
rect 27445 6341 27479 6375
rect 27479 6341 27488 6375
rect 27436 6332 27488 6341
rect 15844 6128 15896 6180
rect 16212 6128 16264 6180
rect 17132 6171 17184 6180
rect 17132 6137 17141 6171
rect 17141 6137 17175 6171
rect 17175 6137 17184 6171
rect 17132 6128 17184 6137
rect 14372 6060 14424 6112
rect 15108 6060 15160 6112
rect 16948 6060 17000 6112
rect 17316 6060 17368 6112
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 17868 6128 17920 6180
rect 17960 6171 18012 6180
rect 17960 6137 17969 6171
rect 17969 6137 18003 6171
rect 18003 6137 18012 6171
rect 17960 6128 18012 6137
rect 20168 6196 20220 6248
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 22560 6196 22612 6248
rect 26516 6264 26568 6316
rect 28908 6307 28960 6316
rect 28908 6273 28917 6307
rect 28917 6273 28951 6307
rect 28951 6273 28960 6307
rect 28908 6264 28960 6273
rect 29092 6264 29144 6316
rect 38200 6264 38252 6316
rect 37004 6196 37056 6248
rect 38936 6196 38988 6248
rect 18052 6060 18104 6112
rect 18788 6060 18840 6112
rect 21180 6128 21232 6180
rect 22928 6060 22980 6112
rect 29000 6128 29052 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6920 5856 6972 5908
rect 12900 5899 12952 5908
rect 12900 5865 12909 5899
rect 12909 5865 12943 5899
rect 12943 5865 12952 5899
rect 12900 5856 12952 5865
rect 13360 5856 13412 5908
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 12440 5652 12492 5704
rect 12900 5584 12952 5636
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 10784 5516 10836 5568
rect 12256 5516 12308 5568
rect 12992 5516 13044 5568
rect 13176 5627 13228 5636
rect 13176 5593 13185 5627
rect 13185 5593 13219 5627
rect 13219 5593 13228 5627
rect 13176 5584 13228 5593
rect 13636 5856 13688 5908
rect 14556 5856 14608 5908
rect 15752 5856 15804 5908
rect 16028 5856 16080 5908
rect 17224 5856 17276 5908
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 18512 5856 18564 5908
rect 19340 5856 19392 5908
rect 19432 5856 19484 5908
rect 23296 5856 23348 5908
rect 24676 5856 24728 5908
rect 32864 5856 32916 5908
rect 18696 5788 18748 5840
rect 16948 5720 17000 5772
rect 18604 5720 18656 5772
rect 24584 5831 24636 5840
rect 24584 5797 24593 5831
rect 24593 5797 24627 5831
rect 24627 5797 24636 5831
rect 24584 5788 24636 5797
rect 22100 5763 22152 5772
rect 22100 5729 22109 5763
rect 22109 5729 22143 5763
rect 22143 5729 22152 5763
rect 25228 5763 25280 5772
rect 22100 5720 22152 5729
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 14096 5652 14148 5704
rect 15016 5652 15068 5704
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 15752 5652 15804 5704
rect 14188 5516 14240 5568
rect 15660 5516 15712 5568
rect 16212 5652 16264 5704
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 16764 5652 16816 5704
rect 17684 5652 17736 5704
rect 18052 5695 18104 5704
rect 18052 5661 18061 5695
rect 18061 5661 18095 5695
rect 18095 5661 18104 5695
rect 18052 5652 18104 5661
rect 18144 5695 18196 5704
rect 18144 5661 18153 5695
rect 18153 5661 18187 5695
rect 18187 5661 18196 5695
rect 18144 5652 18196 5661
rect 18236 5584 18288 5636
rect 16672 5516 16724 5568
rect 19432 5652 19484 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 20444 5584 20496 5636
rect 20536 5584 20588 5636
rect 20904 5584 20956 5636
rect 23480 5652 23532 5704
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 32772 5720 32824 5772
rect 33140 5720 33192 5772
rect 24676 5652 24728 5704
rect 23388 5584 23440 5636
rect 26056 5652 26108 5704
rect 33324 5584 33376 5636
rect 22560 5516 22612 5568
rect 22836 5516 22888 5568
rect 23756 5516 23808 5568
rect 26424 5516 26476 5568
rect 33048 5516 33100 5568
rect 34152 5559 34204 5568
rect 34152 5525 34161 5559
rect 34161 5525 34195 5559
rect 34195 5525 34204 5559
rect 34152 5516 34204 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 7196 5312 7248 5364
rect 9956 5312 10008 5364
rect 10508 5312 10560 5364
rect 12072 5312 12124 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 8208 5176 8260 5228
rect 6552 5108 6604 5160
rect 9128 5176 9180 5228
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 14372 5312 14424 5364
rect 14924 5312 14976 5364
rect 15568 5312 15620 5364
rect 32312 5312 32364 5364
rect 10232 5176 10284 5228
rect 10048 5108 10100 5160
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 11060 5176 11112 5228
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 13728 5244 13780 5296
rect 13912 5244 13964 5296
rect 14556 5244 14608 5296
rect 12624 5176 12676 5228
rect 13268 5176 13320 5228
rect 8116 4972 8168 5024
rect 10324 4972 10376 5024
rect 10968 4972 11020 5024
rect 11888 5083 11940 5092
rect 11888 5049 11897 5083
rect 11897 5049 11931 5083
rect 11931 5049 11940 5083
rect 11888 5040 11940 5049
rect 12164 5040 12216 5092
rect 13912 5040 13964 5092
rect 14188 5176 14240 5228
rect 15108 5244 15160 5296
rect 16672 5244 16724 5296
rect 26516 5244 26568 5296
rect 15200 5176 15252 5228
rect 14648 5108 14700 5160
rect 15752 5108 15804 5160
rect 23388 5176 23440 5228
rect 25228 5176 25280 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 30932 5176 30984 5228
rect 29000 5151 29052 5160
rect 29000 5117 29009 5151
rect 29009 5117 29043 5151
rect 29043 5117 29052 5151
rect 29000 5108 29052 5117
rect 31208 5219 31260 5228
rect 31208 5185 31217 5219
rect 31217 5185 31251 5219
rect 31251 5185 31260 5219
rect 31208 5176 31260 5185
rect 33232 5244 33284 5296
rect 33784 5244 33836 5296
rect 22836 5040 22888 5092
rect 26056 5040 26108 5092
rect 31116 5040 31168 5092
rect 22560 5015 22612 5024
rect 22560 4981 22569 5015
rect 22569 4981 22603 5015
rect 22603 4981 22612 5015
rect 22560 4972 22612 4981
rect 23020 4972 23072 5024
rect 23664 4972 23716 5024
rect 25596 4972 25648 5024
rect 27068 4972 27120 5024
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 30656 4972 30708 5024
rect 32772 5176 32824 5228
rect 31576 5040 31628 5092
rect 32128 5040 32180 5092
rect 32036 4972 32088 5024
rect 33324 4972 33376 5024
rect 34612 5015 34664 5024
rect 34612 4981 34621 5015
rect 34621 4981 34655 5015
rect 34655 4981 34664 5015
rect 34612 4972 34664 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 11336 4768 11388 4820
rect 11428 4768 11480 4820
rect 11796 4768 11848 4820
rect 13084 4768 13136 4820
rect 13360 4768 13412 4820
rect 13820 4768 13872 4820
rect 15568 4768 15620 4820
rect 19156 4768 19208 4820
rect 23388 4768 23440 4820
rect 29368 4811 29420 4820
rect 29368 4777 29377 4811
rect 29377 4777 29411 4811
rect 29411 4777 29420 4811
rect 29368 4768 29420 4777
rect 30656 4811 30708 4820
rect 30656 4777 30665 4811
rect 30665 4777 30699 4811
rect 30699 4777 30708 4811
rect 30656 4768 30708 4777
rect 7840 4564 7892 4616
rect 9680 4564 9732 4616
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 10508 4564 10560 4616
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 11060 4539 11112 4548
rect 11060 4505 11090 4539
rect 11090 4505 11112 4539
rect 11612 4564 11664 4616
rect 12532 4564 12584 4616
rect 12716 4564 12768 4616
rect 13452 4632 13504 4684
rect 11060 4496 11112 4505
rect 11336 4496 11388 4548
rect 13268 4564 13320 4616
rect 13912 4632 13964 4684
rect 14188 4632 14240 4684
rect 15016 4675 15068 4684
rect 15016 4641 15025 4675
rect 15025 4641 15059 4675
rect 15059 4641 15068 4675
rect 15016 4632 15068 4641
rect 15752 4700 15804 4752
rect 18972 4700 19024 4752
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 15568 4564 15620 4616
rect 17132 4564 17184 4616
rect 18604 4564 18656 4616
rect 17868 4496 17920 4548
rect 16396 4428 16448 4480
rect 18144 4428 18196 4480
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 19340 4496 19392 4548
rect 22284 4564 22336 4616
rect 23020 4607 23072 4616
rect 23020 4573 23029 4607
rect 23029 4573 23063 4607
rect 23063 4573 23072 4607
rect 23020 4564 23072 4573
rect 23940 4700 23992 4752
rect 28908 4700 28960 4752
rect 24032 4632 24084 4684
rect 23756 4607 23808 4616
rect 23756 4573 23765 4607
rect 23765 4573 23799 4607
rect 23799 4573 23808 4607
rect 23756 4564 23808 4573
rect 24400 4607 24452 4616
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 26240 4564 26292 4616
rect 22836 4428 22888 4480
rect 23112 4471 23164 4480
rect 23112 4437 23121 4471
rect 23121 4437 23155 4471
rect 23155 4437 23164 4471
rect 23112 4428 23164 4437
rect 25412 4496 25464 4548
rect 28356 4632 28408 4684
rect 27620 4607 27672 4616
rect 27620 4573 27629 4607
rect 27629 4573 27663 4607
rect 27663 4573 27672 4607
rect 27620 4564 27672 4573
rect 29184 4496 29236 4548
rect 32036 4632 32088 4684
rect 32772 4632 32824 4684
rect 34612 4700 34664 4752
rect 34152 4564 34204 4616
rect 34612 4564 34664 4616
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 8208 4156 8260 4208
rect 9864 4156 9916 4208
rect 7196 4020 7248 4072
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 8116 4020 8168 4072
rect 10140 4088 10192 4140
rect 9680 4020 9732 4072
rect 10416 4020 10468 4072
rect 11336 4088 11388 4140
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12256 4156 12308 4208
rect 12072 4088 12124 4097
rect 11428 4020 11480 4072
rect 11612 4020 11664 4072
rect 12348 4063 12400 4072
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 12716 4020 12768 4072
rect 12900 4020 12952 4072
rect 11980 3995 12032 4004
rect 11980 3961 11989 3995
rect 11989 3961 12023 3995
rect 12023 3961 12032 3995
rect 13452 4020 13504 4072
rect 14924 4224 14976 4276
rect 14372 4156 14424 4208
rect 14280 4088 14332 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 17960 4224 18012 4276
rect 18972 4224 19024 4276
rect 23112 4224 23164 4276
rect 24676 4224 24728 4276
rect 16212 4156 16264 4208
rect 11980 3952 12032 3961
rect 10600 3884 10652 3936
rect 12164 3884 12216 3936
rect 13084 3952 13136 4004
rect 13544 3884 13596 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 15752 4088 15804 4140
rect 16120 4088 16172 4140
rect 16396 4088 16448 4140
rect 17040 4088 17092 4140
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 15660 3952 15712 4004
rect 15936 3884 15988 3936
rect 16488 3952 16540 4004
rect 17408 4020 17460 4072
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 17500 3995 17552 4004
rect 17500 3961 17509 3995
rect 17509 3961 17543 3995
rect 17543 3961 17552 3995
rect 17500 3952 17552 3961
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17316 3884 17368 3936
rect 21640 4199 21692 4208
rect 21640 4165 21649 4199
rect 21649 4165 21683 4199
rect 21683 4165 21692 4199
rect 21640 4156 21692 4165
rect 22836 4156 22888 4208
rect 23204 4156 23256 4208
rect 31852 4224 31904 4276
rect 34612 4224 34664 4276
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18328 4131 18380 4140
rect 18328 4097 18337 4131
rect 18337 4097 18371 4131
rect 18371 4097 18380 4131
rect 18328 4088 18380 4097
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 18604 4088 18656 4140
rect 18880 4088 18932 4140
rect 19156 4088 19208 4140
rect 19432 4088 19484 4140
rect 19984 4088 20036 4140
rect 20168 4088 20220 4140
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 19340 4020 19392 4072
rect 23848 4020 23900 4072
rect 18972 3995 19024 4004
rect 18972 3961 18981 3995
rect 18981 3961 19015 3995
rect 19015 3961 19024 3995
rect 18972 3952 19024 3961
rect 22284 3952 22336 4004
rect 23480 3952 23532 4004
rect 23572 3995 23624 4004
rect 23572 3961 23581 3995
rect 23581 3961 23615 3995
rect 23615 3961 23624 3995
rect 23572 3952 23624 3961
rect 23664 3995 23716 4004
rect 23664 3961 23673 3995
rect 23673 3961 23707 3995
rect 23707 3961 23716 3995
rect 23664 3952 23716 3961
rect 18420 3884 18472 3936
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 22468 3884 22520 3936
rect 23296 3927 23348 3936
rect 23296 3893 23305 3927
rect 23305 3893 23339 3927
rect 23339 3893 23348 3927
rect 23296 3884 23348 3893
rect 24584 4131 24636 4140
rect 24584 4097 24593 4131
rect 24593 4097 24627 4131
rect 24627 4097 24636 4131
rect 24584 4088 24636 4097
rect 29184 4156 29236 4208
rect 36084 4156 36136 4208
rect 24492 3952 24544 4004
rect 28908 4088 28960 4140
rect 33048 4088 33100 4140
rect 34796 4088 34848 4140
rect 37096 4131 37148 4140
rect 37096 4097 37105 4131
rect 37105 4097 37139 4131
rect 37139 4097 37148 4131
rect 37096 4088 37148 4097
rect 25412 3952 25464 4004
rect 27528 3952 27580 4004
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 30932 4063 30984 4072
rect 30932 4029 30941 4063
rect 30941 4029 30975 4063
rect 30975 4029 30984 4063
rect 30932 4020 30984 4029
rect 36820 4063 36872 4072
rect 36820 4029 36829 4063
rect 36829 4029 36863 4063
rect 36863 4029 36872 4063
rect 36820 4020 36872 4029
rect 24860 3884 24912 3936
rect 26056 3884 26108 3936
rect 27620 3884 27672 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8208 3680 8260 3732
rect 9312 3680 9364 3732
rect 9864 3680 9916 3732
rect 10968 3680 11020 3732
rect 11336 3612 11388 3664
rect 11704 3612 11756 3664
rect 12164 3612 12216 3664
rect 12256 3655 12308 3664
rect 12256 3621 12265 3655
rect 12265 3621 12299 3655
rect 12299 3621 12308 3655
rect 12256 3612 12308 3621
rect 12716 3680 12768 3732
rect 13728 3680 13780 3732
rect 14464 3680 14516 3732
rect 15752 3723 15804 3732
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 9496 3476 9548 3528
rect 9680 3476 9732 3528
rect 11520 3476 11572 3528
rect 12072 3476 12124 3528
rect 10232 3340 10284 3392
rect 10968 3340 11020 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 12348 3544 12400 3596
rect 13360 3612 13412 3664
rect 14924 3612 14976 3664
rect 16396 3680 16448 3732
rect 18788 3680 18840 3732
rect 18880 3680 18932 3732
rect 22192 3680 22244 3732
rect 22836 3680 22888 3732
rect 22928 3680 22980 3732
rect 23940 3723 23992 3732
rect 23940 3689 23949 3723
rect 23949 3689 23983 3723
rect 23983 3689 23992 3723
rect 23940 3680 23992 3689
rect 24492 3680 24544 3732
rect 24860 3680 24912 3732
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 12532 3476 12584 3528
rect 16488 3544 16540 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 22468 3612 22520 3664
rect 23572 3655 23624 3664
rect 23572 3621 23581 3655
rect 23581 3621 23615 3655
rect 23615 3621 23624 3655
rect 23572 3612 23624 3621
rect 29000 3680 29052 3732
rect 29460 3680 29512 3732
rect 36820 3680 36872 3732
rect 20168 3544 20220 3596
rect 13360 3497 13412 3528
rect 12256 3408 12308 3460
rect 12716 3408 12768 3460
rect 13360 3476 13391 3497
rect 13391 3476 13412 3497
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 13728 3476 13780 3528
rect 14188 3476 14240 3528
rect 14556 3476 14608 3528
rect 14832 3476 14884 3528
rect 13176 3408 13228 3460
rect 13912 3408 13964 3460
rect 14464 3451 14516 3460
rect 14464 3417 14473 3451
rect 14473 3417 14507 3451
rect 14507 3417 14516 3451
rect 14464 3408 14516 3417
rect 16212 3476 16264 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 18236 3476 18288 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 20812 3476 20864 3528
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 15752 3340 15804 3392
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 16304 3340 16356 3392
rect 20996 3408 21048 3460
rect 22284 3408 22336 3460
rect 23204 3476 23256 3528
rect 24400 3544 24452 3596
rect 27620 3544 27672 3596
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 23480 3408 23532 3460
rect 26700 3519 26752 3528
rect 26700 3485 26709 3519
rect 26709 3485 26743 3519
rect 26743 3485 26752 3519
rect 26700 3476 26752 3485
rect 36544 3476 36596 3528
rect 19432 3383 19484 3392
rect 19432 3349 19441 3383
rect 19441 3349 19475 3383
rect 19475 3349 19484 3383
rect 19432 3340 19484 3349
rect 22560 3340 22612 3392
rect 27528 3408 27580 3460
rect 29184 3340 29236 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 9496 3136 9548 3188
rect 9312 3068 9364 3120
rect 8116 3000 8168 3052
rect 11520 3136 11572 3188
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 13360 3136 13412 3188
rect 13912 3136 13964 3188
rect 14740 3136 14792 3188
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 12992 3068 13044 3120
rect 16304 3136 16356 3188
rect 16580 3136 16632 3188
rect 19248 3136 19300 3188
rect 19340 3136 19392 3188
rect 19432 3136 19484 3188
rect 20168 3136 20220 3188
rect 16028 3068 16080 3120
rect 15660 3000 15712 3052
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 15936 3000 15988 3052
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 13452 2932 13504 2984
rect 15476 2932 15528 2984
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 8668 2864 8720 2916
rect 13176 2864 13228 2916
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 10692 2839 10744 2848
rect 10692 2805 10701 2839
rect 10701 2805 10735 2839
rect 10735 2805 10744 2839
rect 10692 2796 10744 2805
rect 20996 3068 21048 3120
rect 22468 3068 22520 3120
rect 23480 3136 23532 3188
rect 23572 3136 23624 3188
rect 24860 3136 24912 3188
rect 25412 3068 25464 3120
rect 26056 3068 26108 3120
rect 29276 3068 29328 3120
rect 31208 3136 31260 3188
rect 36544 3179 36596 3188
rect 36544 3145 36553 3179
rect 36553 3145 36587 3179
rect 36587 3145 36596 3179
rect 36544 3136 36596 3145
rect 22192 3041 22244 3052
rect 22192 3007 22201 3041
rect 22201 3007 22235 3041
rect 22235 3007 22244 3041
rect 22192 3000 22244 3007
rect 18972 2907 19024 2916
rect 18972 2873 18981 2907
rect 18981 2873 19015 2907
rect 19015 2873 19024 2907
rect 18972 2864 19024 2873
rect 22928 3000 22980 3052
rect 22284 2839 22336 2848
rect 22284 2805 22293 2839
rect 22293 2805 22327 2839
rect 22327 2805 22336 2839
rect 22284 2796 22336 2805
rect 24400 3000 24452 3052
rect 27620 3000 27672 3052
rect 23480 2975 23532 2984
rect 23480 2941 23489 2975
rect 23489 2941 23523 2975
rect 23523 2941 23532 2975
rect 23480 2932 23532 2941
rect 28816 2975 28868 2984
rect 28816 2941 28825 2975
rect 28825 2941 28859 2975
rect 28859 2941 28868 2975
rect 28816 2932 28868 2941
rect 43260 2864 43312 2916
rect 24860 2796 24912 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2044 2592 2096 2644
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 18972 2592 19024 2644
rect 26700 2592 26752 2644
rect 43260 2635 43312 2644
rect 43260 2601 43269 2635
rect 43269 2601 43303 2635
rect 43303 2601 43312 2635
rect 43260 2592 43312 2601
rect 10692 2456 10744 2508
rect 28816 2456 28868 2508
rect 20 2388 72 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 24860 2388 24912 2440
rect 26148 2388 26200 2440
rect 43168 2388 43220 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 6458 47077 6514 47877
rect 14830 47077 14886 47877
rect 23846 47077 23902 47877
rect 32218 47077 32274 47877
rect 41234 47077 41290 47877
rect 1398 45656 1454 45665
rect 1398 45591 1454 45600
rect 1412 45490 1440 45591
rect 6472 45490 6500 47077
rect 14844 45558 14872 47077
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 14832 45552 14884 45558
rect 23860 45554 23888 47077
rect 32232 45558 32260 47077
rect 23860 45526 23980 45554
rect 14832 45494 14884 45500
rect 23952 45490 23980 45526
rect 32220 45552 32272 45558
rect 32220 45494 32272 45500
rect 41248 45490 41276 47077
rect 1400 45484 1452 45490
rect 1400 45426 1452 45432
rect 6460 45484 6512 45490
rect 6460 45426 6512 45432
rect 23940 45484 23992 45490
rect 23940 45426 23992 45432
rect 41236 45484 41288 45490
rect 41236 45426 41288 45432
rect 5908 45280 5960 45286
rect 5908 45222 5960 45228
rect 7288 45280 7340 45286
rect 7288 45222 7340 45228
rect 15108 45280 15160 45286
rect 15108 45222 15160 45228
rect 24308 45280 24360 45286
rect 24308 45222 24360 45228
rect 32312 45280 32364 45286
rect 32312 45222 32364 45228
rect 41328 45280 41380 45286
rect 41328 45222 41380 45228
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 5920 45014 5948 45222
rect 5908 45008 5960 45014
rect 5908 44950 5960 44956
rect 6644 44940 6696 44946
rect 6644 44882 6696 44888
rect 6092 44736 6144 44742
rect 6092 44678 6144 44684
rect 6104 44538 6132 44678
rect 6092 44532 6144 44538
rect 6092 44474 6144 44480
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 6656 42770 6684 44882
rect 7300 44402 7328 45222
rect 15120 45082 15148 45222
rect 15108 45076 15160 45082
rect 15108 45018 15160 45024
rect 16120 45008 16172 45014
rect 16172 44956 16528 44962
rect 16120 44950 16528 44956
rect 16132 44946 16528 44950
rect 16132 44940 16540 44946
rect 16132 44934 16488 44940
rect 16488 44882 16540 44888
rect 9864 44872 9916 44878
rect 9864 44814 9916 44820
rect 12440 44872 12492 44878
rect 12440 44814 12492 44820
rect 14096 44872 14148 44878
rect 14096 44814 14148 44820
rect 15844 44872 15896 44878
rect 15844 44814 15896 44820
rect 16028 44872 16080 44878
rect 16028 44814 16080 44820
rect 16120 44872 16172 44878
rect 16120 44814 16172 44820
rect 7288 44396 7340 44402
rect 7288 44338 7340 44344
rect 6920 44192 6972 44198
rect 6920 44134 6972 44140
rect 6932 43722 6960 44134
rect 7012 43852 7064 43858
rect 7012 43794 7064 43800
rect 6920 43716 6972 43722
rect 6920 43658 6972 43664
rect 6644 42764 6696 42770
rect 6644 42706 6696 42712
rect 5540 42696 5592 42702
rect 5540 42638 5592 42644
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5552 37262 5580 42638
rect 6656 41414 6684 42706
rect 7024 42226 7052 43794
rect 7012 42220 7064 42226
rect 7012 42162 7064 42168
rect 6564 41386 6684 41414
rect 940 37256 992 37262
rect 940 37198 992 37204
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 952 36825 980 37198
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1780 36718 1808 37198
rect 2136 37120 2188 37126
rect 2136 37062 2188 37068
rect 1768 36712 1820 36718
rect 1768 36654 1820 36660
rect 940 27464 992 27470
rect 940 27406 992 27412
rect 952 27305 980 27406
rect 1584 27328 1636 27334
rect 938 27296 994 27305
rect 1584 27270 1636 27276
rect 938 27231 994 27240
rect 1596 26586 1624 27270
rect 1584 26580 1636 26586
rect 1584 26522 1636 26528
rect 1780 18834 1808 36654
rect 2148 36650 2176 37062
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 6368 36712 6420 36718
rect 6368 36654 6420 36660
rect 2136 36644 2188 36650
rect 2136 36586 2188 36592
rect 2228 36576 2280 36582
rect 2228 36518 2280 36524
rect 2240 35698 2268 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36378 4660 36654
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 5828 36106 5856 36518
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 4068 36100 4120 36106
rect 4068 36042 4120 36048
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 4080 35834 4108 36042
rect 5724 36032 5776 36038
rect 5724 35974 5776 35980
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 5540 35760 5592 35766
rect 5540 35702 5592 35708
rect 2228 35692 2280 35698
rect 2228 35634 2280 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 5552 35290 5580 35702
rect 5632 35488 5684 35494
rect 5632 35430 5684 35436
rect 5540 35284 5592 35290
rect 5540 35226 5592 35232
rect 5448 35216 5500 35222
rect 5448 35158 5500 35164
rect 5080 35080 5132 35086
rect 5080 35022 5132 35028
rect 5092 34542 5120 35022
rect 5460 34542 5488 35158
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5080 34536 5132 34542
rect 5080 34478 5132 34484
rect 5448 34536 5500 34542
rect 5448 34478 5500 34484
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5552 34202 5580 35022
rect 5644 34746 5672 35430
rect 5632 34740 5684 34746
rect 5632 34682 5684 34688
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5172 33516 5224 33522
rect 5172 33458 5224 33464
rect 3884 33448 3936 33454
rect 3884 33390 3936 33396
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 3896 32910 3924 33390
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33390
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 3884 32904 3936 32910
rect 3884 32846 3936 32852
rect 3896 31890 3924 32846
rect 5184 32298 5212 33458
rect 5552 32910 5580 33798
rect 5736 32910 5764 35974
rect 6104 35834 6132 36110
rect 6092 35828 6144 35834
rect 6092 35770 6144 35776
rect 6380 35442 6408 36654
rect 6012 35414 6408 35442
rect 6012 34746 6040 35414
rect 6092 35284 6144 35290
rect 6092 35226 6144 35232
rect 6104 34746 6132 35226
rect 6380 34762 6408 35414
rect 6000 34740 6052 34746
rect 6000 34682 6052 34688
rect 6092 34740 6144 34746
rect 6380 34734 6500 34762
rect 6092 34682 6144 34688
rect 6104 34134 6132 34682
rect 6184 34672 6236 34678
rect 6184 34614 6236 34620
rect 6092 34128 6144 34134
rect 6092 34070 6144 34076
rect 6196 33998 6224 34614
rect 6472 34610 6500 34734
rect 6368 34604 6420 34610
rect 6368 34546 6420 34552
rect 6460 34604 6512 34610
rect 6460 34546 6512 34552
rect 6380 33998 6408 34546
rect 6184 33992 6236 33998
rect 6184 33934 6236 33940
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6380 33658 6408 33934
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5828 33114 5856 33254
rect 5816 33108 5868 33114
rect 5816 33050 5868 33056
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3884 31884 3936 31890
rect 3884 31826 3936 31832
rect 3896 30938 3924 31826
rect 5184 31754 5212 32234
rect 5816 32224 5868 32230
rect 5816 32166 5868 32172
rect 5828 31890 5856 32166
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 6196 31754 6224 32370
rect 6564 31754 6592 41386
rect 7104 39976 7156 39982
rect 7104 39918 7156 39924
rect 7116 39642 7144 39918
rect 7104 39636 7156 39642
rect 7104 39578 7156 39584
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 6736 38412 6788 38418
rect 6736 38354 6788 38360
rect 6748 37942 6776 38354
rect 7024 38282 7052 38694
rect 7012 38276 7064 38282
rect 7012 38218 7064 38224
rect 6736 37936 6788 37942
rect 6736 37878 6788 37884
rect 6748 36854 6776 37878
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 6932 37466 6960 37742
rect 6920 37460 6972 37466
rect 6920 37402 6972 37408
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 6748 36242 6776 36790
rect 6736 36236 6788 36242
rect 6736 36178 6788 36184
rect 6748 35154 6776 36178
rect 7196 36100 7248 36106
rect 7196 36042 7248 36048
rect 7208 35834 7236 36042
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 6920 35692 6972 35698
rect 6920 35634 6972 35640
rect 6736 35148 6788 35154
rect 6736 35090 6788 35096
rect 6736 34944 6788 34950
rect 6736 34886 6788 34892
rect 6748 34746 6776 34886
rect 6644 34740 6696 34746
rect 6644 34682 6696 34688
rect 6736 34740 6788 34746
rect 6736 34682 6788 34688
rect 6656 34610 6684 34682
rect 6644 34604 6696 34610
rect 6644 34546 6696 34552
rect 6932 33096 6960 35634
rect 6840 33068 7144 33096
rect 6840 32842 6868 33068
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 6828 32836 6880 32842
rect 6828 32778 6880 32784
rect 6932 31890 6960 32914
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 5172 31748 5224 31754
rect 6196 31726 6316 31754
rect 5172 31690 5224 31696
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3884 30932 3936 30938
rect 3884 30874 3936 30880
rect 3896 29850 3924 30874
rect 5184 30734 5212 31690
rect 6288 31482 6316 31726
rect 6380 31726 6592 31754
rect 6276 31476 6328 31482
rect 6276 31418 6328 31424
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3884 29844 3936 29850
rect 3884 29786 3936 29792
rect 5184 29646 5212 30670
rect 5448 30048 5500 30054
rect 5448 29990 5500 29996
rect 5460 29850 5488 29990
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 5172 29640 5224 29646
rect 5172 29582 5224 29588
rect 4068 29572 4120 29578
rect 4068 29514 4120 29520
rect 4080 29306 4108 29514
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 5460 29238 5488 29786
rect 5552 29238 5580 31282
rect 6000 31136 6052 31142
rect 6000 31078 6052 31084
rect 6012 30938 6040 31078
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 6092 30728 6144 30734
rect 6092 30670 6144 30676
rect 5644 30394 5672 30670
rect 5816 30660 5868 30666
rect 5816 30602 5868 30608
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 5724 30184 5776 30190
rect 5724 30126 5776 30132
rect 5736 29578 5764 30126
rect 5828 30054 5856 30602
rect 6104 30394 6132 30670
rect 6092 30388 6144 30394
rect 6092 30330 6144 30336
rect 6000 30184 6052 30190
rect 6000 30126 6052 30132
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 6012 29714 6040 30126
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5724 29572 5776 29578
rect 5724 29514 5776 29520
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 5448 29232 5500 29238
rect 5448 29174 5500 29180
rect 5540 29232 5592 29238
rect 5540 29174 5592 29180
rect 6196 28966 6224 29446
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5552 28082 5580 28562
rect 6092 28416 6144 28422
rect 6092 28358 6144 28364
rect 6104 28082 6132 28358
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5816 28076 5868 28082
rect 5816 28018 5868 28024
rect 6092 28076 6144 28082
rect 6380 28064 6408 31726
rect 6932 31142 6960 31826
rect 6920 31136 6972 31142
rect 6920 31078 6972 31084
rect 6932 30190 6960 31078
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 6552 29572 6604 29578
rect 6552 29514 6604 29520
rect 6564 28626 6592 29514
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6092 28018 6144 28024
rect 6288 28036 6408 28064
rect 5356 27872 5408 27878
rect 5828 27860 5856 28018
rect 5908 27872 5960 27878
rect 5828 27832 5908 27860
rect 5356 27814 5408 27820
rect 5908 27814 5960 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5368 27674 5396 27814
rect 5356 27668 5408 27674
rect 5356 27610 5408 27616
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 6288 26450 6316 28036
rect 6368 27940 6420 27946
rect 6368 27882 6420 27888
rect 6380 27674 6408 27882
rect 6368 27668 6420 27674
rect 6368 27610 6420 27616
rect 6932 27538 6960 30126
rect 6920 27532 6972 27538
rect 6920 27474 6972 27480
rect 6644 27464 6696 27470
rect 6644 27406 6696 27412
rect 6656 26926 6684 27406
rect 6644 26920 6696 26926
rect 6644 26862 6696 26868
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 5736 26042 5764 26386
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5828 25362 5856 25774
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 6196 25362 6224 25638
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6288 22094 6316 26386
rect 6656 25838 6684 26862
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6288 22066 6408 22094
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1780 9042 1808 18770
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 18426 2268 18566
rect 3160 18426 3188 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 16250 2820 17614
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 3344 15910 3372 18022
rect 3712 17882 3740 18158
rect 4632 18086 4660 18702
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4724 18358 4752 18566
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 4724 17678 4752 18294
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17338 4384 17478
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4724 16998 4752 17614
rect 5092 17338 5120 18702
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6104 17746 6132 18090
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6196 17610 6224 18022
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4724 16250 4752 16934
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 15570 3372 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3344 15026 3372 15506
rect 4724 15434 4752 16186
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15706 5396 15982
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15094 3832 15302
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 4724 15026 4752 15370
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13258 4108 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4632 12986 4660 13806
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12918 4752 14962
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14618 5212 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5552 14074 5580 14962
rect 5644 14958 5672 15846
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5736 14278 5764 16050
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6012 15706 6040 15982
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6380 14890 6408 22066
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6932 19514 6960 21286
rect 7024 19854 7052 32438
rect 7116 31754 7144 33068
rect 7196 32836 7248 32842
rect 7196 32778 7248 32784
rect 7208 32570 7236 32778
rect 7196 32564 7248 32570
rect 7196 32506 7248 32512
rect 7300 32502 7328 44338
rect 8208 44192 8260 44198
rect 8208 44134 8260 44140
rect 8220 43858 8248 44134
rect 8208 43852 8260 43858
rect 8208 43794 8260 43800
rect 9876 43790 9904 44814
rect 10508 44804 10560 44810
rect 10508 44746 10560 44752
rect 11796 44804 11848 44810
rect 11796 44746 11848 44752
rect 10520 44538 10548 44746
rect 10508 44532 10560 44538
rect 10508 44474 10560 44480
rect 11808 44198 11836 44746
rect 12072 44736 12124 44742
rect 12072 44678 12124 44684
rect 12084 44538 12112 44678
rect 12072 44532 12124 44538
rect 12072 44474 12124 44480
rect 11980 44328 12032 44334
rect 11980 44270 12032 44276
rect 12072 44328 12124 44334
rect 12072 44270 12124 44276
rect 11796 44192 11848 44198
rect 11796 44134 11848 44140
rect 9864 43784 9916 43790
rect 9864 43726 9916 43732
rect 8484 43648 8536 43654
rect 8536 43608 8708 43636
rect 8484 43590 8536 43596
rect 7380 42152 7432 42158
rect 7380 42094 7432 42100
rect 7392 41818 7420 42094
rect 7380 41812 7432 41818
rect 7380 41754 7432 41760
rect 8484 41472 8536 41478
rect 8484 41414 8536 41420
rect 8312 41386 8524 41414
rect 7840 38888 7892 38894
rect 7840 38830 7892 38836
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 7392 35086 7420 35974
rect 7564 35692 7616 35698
rect 7564 35634 7616 35640
rect 7656 35692 7708 35698
rect 7656 35634 7708 35640
rect 7472 35216 7524 35222
rect 7472 35158 7524 35164
rect 7380 35080 7432 35086
rect 7380 35022 7432 35028
rect 7484 34746 7512 35158
rect 7576 35018 7604 35634
rect 7668 35290 7696 35634
rect 7656 35284 7708 35290
rect 7656 35226 7708 35232
rect 7564 35012 7616 35018
rect 7564 34954 7616 34960
rect 7472 34740 7524 34746
rect 7472 34682 7524 34688
rect 7288 32496 7340 32502
rect 7288 32438 7340 32444
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7196 32020 7248 32026
rect 7196 31962 7248 31968
rect 7104 31748 7156 31754
rect 7104 31690 7156 31696
rect 7116 31346 7144 31690
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7208 30802 7236 31962
rect 7380 31408 7432 31414
rect 7380 31350 7432 31356
rect 7196 30796 7248 30802
rect 7196 30738 7248 30744
rect 7392 30666 7420 31350
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 7380 30660 7432 30666
rect 7380 30602 7432 30608
rect 7392 30394 7420 30602
rect 7576 30394 7604 30670
rect 7380 30388 7432 30394
rect 7380 30330 7432 30336
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 7392 29646 7420 30330
rect 7564 30116 7616 30122
rect 7564 30058 7616 30064
rect 7380 29640 7432 29646
rect 7576 29628 7604 30058
rect 7668 29866 7696 32302
rect 7760 32026 7788 37062
rect 7748 32020 7800 32026
rect 7748 31962 7800 31968
rect 7748 31748 7800 31754
rect 7748 31690 7800 31696
rect 7760 31142 7788 31690
rect 7748 31136 7800 31142
rect 7748 31078 7800 31084
rect 7748 30660 7800 30666
rect 7852 30648 7880 38830
rect 8208 38820 8260 38826
rect 8208 38762 8260 38768
rect 8220 37330 8248 38762
rect 8208 37324 8260 37330
rect 8208 37266 8260 37272
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8220 36378 8248 36722
rect 8312 36718 8340 41386
rect 8484 40520 8536 40526
rect 8484 40462 8536 40468
rect 8496 39846 8524 40462
rect 8576 40384 8628 40390
rect 8576 40326 8628 40332
rect 8588 40186 8616 40326
rect 8576 40180 8628 40186
rect 8576 40122 8628 40128
rect 8680 39930 8708 43608
rect 8852 42628 8904 42634
rect 8852 42570 8904 42576
rect 8864 42294 8892 42570
rect 8944 42560 8996 42566
rect 8944 42502 8996 42508
rect 9496 42560 9548 42566
rect 9496 42502 9548 42508
rect 8852 42288 8904 42294
rect 8852 42230 8904 42236
rect 8956 41818 8984 42502
rect 9508 42294 9536 42502
rect 9876 42362 9904 43726
rect 10876 43716 10928 43722
rect 10876 43658 10928 43664
rect 10888 43450 10916 43658
rect 10968 43648 11020 43654
rect 10968 43590 11020 43596
rect 10876 43444 10928 43450
rect 10876 43386 10928 43392
rect 10876 43308 10928 43314
rect 10796 43268 10876 43296
rect 10796 42809 10824 43268
rect 10876 43250 10928 43256
rect 10980 43194 11008 43590
rect 10888 43166 11008 43194
rect 10782 42800 10838 42809
rect 10782 42735 10838 42744
rect 10140 42696 10192 42702
rect 10140 42638 10192 42644
rect 10048 42560 10100 42566
rect 10048 42502 10100 42508
rect 9864 42356 9916 42362
rect 9864 42298 9916 42304
rect 9496 42288 9548 42294
rect 9496 42230 9548 42236
rect 8944 41812 8996 41818
rect 8944 41754 8996 41760
rect 9876 41682 9904 42298
rect 9588 41676 9640 41682
rect 9588 41618 9640 41624
rect 9864 41676 9916 41682
rect 9864 41618 9916 41624
rect 9600 41414 9628 41618
rect 9680 41472 9732 41478
rect 9680 41414 9732 41420
rect 9508 41386 9628 41414
rect 9692 41386 9812 41414
rect 9404 40452 9456 40458
rect 9404 40394 9456 40400
rect 8760 40384 8812 40390
rect 8760 40326 8812 40332
rect 8772 40186 8800 40326
rect 9416 40186 9444 40394
rect 8760 40180 8812 40186
rect 8760 40122 8812 40128
rect 9404 40180 9456 40186
rect 9404 40122 9456 40128
rect 9220 40044 9272 40050
rect 9220 39986 9272 39992
rect 9128 39976 9180 39982
rect 8680 39902 8800 39930
rect 9128 39918 9180 39924
rect 8484 39840 8536 39846
rect 8484 39782 8536 39788
rect 8668 39840 8720 39846
rect 8668 39782 8720 39788
rect 8496 39506 8524 39782
rect 8484 39500 8536 39506
rect 8484 39442 8536 39448
rect 8680 39438 8708 39782
rect 8668 39432 8720 39438
rect 8668 39374 8720 39380
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 8404 37942 8432 38490
rect 8392 37936 8444 37942
rect 8392 37878 8444 37884
rect 8404 37754 8432 37878
rect 8404 37726 8524 37754
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8404 37262 8432 37606
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8300 36712 8352 36718
rect 8352 36672 8432 36700
rect 8300 36654 8352 36660
rect 8208 36372 8260 36378
rect 8208 36314 8260 36320
rect 8220 34898 8248 36314
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8128 34870 8248 34898
rect 8024 33448 8076 33454
rect 8024 33390 8076 33396
rect 8036 32570 8064 33390
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 8024 32428 8076 32434
rect 8024 32370 8076 32376
rect 8036 31958 8064 32370
rect 8024 31952 8076 31958
rect 8024 31894 8076 31900
rect 8128 31414 8156 34870
rect 8312 34746 8340 35090
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 8404 33658 8432 36672
rect 8496 36174 8524 37726
rect 8668 36576 8720 36582
rect 8668 36518 8720 36524
rect 8680 36310 8708 36518
rect 8668 36304 8720 36310
rect 8668 36246 8720 36252
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 8484 35216 8536 35222
rect 8484 35158 8536 35164
rect 8496 34610 8524 35158
rect 8668 34944 8720 34950
rect 8668 34886 8720 34892
rect 8680 34746 8708 34886
rect 8668 34740 8720 34746
rect 8668 34682 8720 34688
rect 8484 34604 8536 34610
rect 8484 34546 8536 34552
rect 8668 34536 8720 34542
rect 8668 34478 8720 34484
rect 8392 33652 8444 33658
rect 8392 33594 8444 33600
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 8312 31754 8340 33050
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 8496 32314 8524 32778
rect 8404 32298 8524 32314
rect 8392 32292 8524 32298
rect 8444 32286 8524 32292
rect 8392 32234 8444 32240
rect 8484 32224 8536 32230
rect 8484 32166 8536 32172
rect 8496 31804 8524 32166
rect 8576 31816 8628 31822
rect 8496 31776 8576 31804
rect 8300 31748 8352 31754
rect 8300 31690 8352 31696
rect 8392 31748 8444 31754
rect 8392 31690 8444 31696
rect 8404 31634 8432 31690
rect 8312 31606 8432 31634
rect 8116 31408 8168 31414
rect 8116 31350 8168 31356
rect 8312 31210 8340 31606
rect 8496 31482 8524 31776
rect 8576 31758 8628 31764
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8588 31346 8616 31622
rect 8680 31346 8708 34478
rect 8772 31754 8800 39902
rect 9036 38888 9088 38894
rect 9036 38830 9088 38836
rect 9048 38418 9076 38830
rect 9036 38412 9088 38418
rect 9036 38354 9088 38360
rect 8944 37800 8996 37806
rect 8944 37742 8996 37748
rect 8956 37466 8984 37742
rect 8944 37460 8996 37466
rect 8944 37402 8996 37408
rect 8852 36304 8904 36310
rect 8852 36246 8904 36252
rect 8864 35086 8892 36246
rect 8852 35080 8904 35086
rect 8852 35022 8904 35028
rect 8944 35080 8996 35086
rect 8944 35022 8996 35028
rect 8956 34762 8984 35022
rect 8864 34734 8984 34762
rect 8864 34610 8892 34734
rect 8852 34604 8904 34610
rect 8852 34546 8904 34552
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8852 34468 8904 34474
rect 8852 34410 8904 34416
rect 8864 33998 8892 34410
rect 8852 33992 8904 33998
rect 8852 33934 8904 33940
rect 8956 33862 8984 34546
rect 9036 34400 9088 34406
rect 9036 34342 9088 34348
rect 9048 33998 9076 34342
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 9140 33114 9168 39918
rect 9232 38962 9260 39986
rect 9508 39982 9536 41386
rect 9680 40384 9732 40390
rect 9680 40326 9732 40332
rect 9692 40050 9720 40326
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9496 39976 9548 39982
rect 9496 39918 9548 39924
rect 9404 39500 9456 39506
rect 9404 39442 9456 39448
rect 9220 38956 9272 38962
rect 9220 38898 9272 38904
rect 9220 38276 9272 38282
rect 9220 38218 9272 38224
rect 9232 37398 9260 38218
rect 9416 37874 9444 39442
rect 9508 38894 9536 39918
rect 9588 39296 9640 39302
rect 9588 39238 9640 39244
rect 9600 39098 9628 39238
rect 9588 39092 9640 39098
rect 9588 39034 9640 39040
rect 9496 38888 9548 38894
rect 9496 38830 9548 38836
rect 9600 38554 9628 39034
rect 9588 38548 9640 38554
rect 9588 38490 9640 38496
rect 9692 38350 9720 39986
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 9404 37868 9456 37874
rect 9404 37810 9456 37816
rect 9220 37392 9272 37398
rect 9220 37334 9272 37340
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9416 36242 9444 36654
rect 9404 36236 9456 36242
rect 9404 36178 9456 36184
rect 9416 35086 9444 36178
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9416 34746 9444 35022
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9312 34400 9364 34406
rect 9312 34342 9364 34348
rect 9324 34202 9352 34342
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9784 33386 9812 41386
rect 9876 40934 9904 41618
rect 10060 41614 10088 42502
rect 10152 41818 10180 42638
rect 10140 41812 10192 41818
rect 10140 41754 10192 41760
rect 10048 41608 10100 41614
rect 10048 41550 10100 41556
rect 10508 41540 10560 41546
rect 10508 41482 10560 41488
rect 10520 41274 10548 41482
rect 10508 41268 10560 41274
rect 10508 41210 10560 41216
rect 9864 40928 9916 40934
rect 9864 40870 9916 40876
rect 9876 40594 9904 40870
rect 9864 40588 9916 40594
rect 9864 40530 9916 40536
rect 10796 40390 10824 42735
rect 10888 41138 10916 43166
rect 10968 42696 11020 42702
rect 10968 42638 11020 42644
rect 10980 42362 11008 42638
rect 10968 42356 11020 42362
rect 10968 42298 11020 42304
rect 11808 42294 11836 44134
rect 11992 43382 12020 44270
rect 12084 43858 12112 44270
rect 12072 43852 12124 43858
rect 12072 43794 12124 43800
rect 11980 43376 12032 43382
rect 11980 43318 12032 43324
rect 11980 42696 12032 42702
rect 11980 42638 12032 42644
rect 11796 42288 11848 42294
rect 11796 42230 11848 42236
rect 11244 42152 11296 42158
rect 11244 42094 11296 42100
rect 10876 41132 10928 41138
rect 10876 41074 10928 41080
rect 10888 40458 10916 41074
rect 10876 40452 10928 40458
rect 10876 40394 10928 40400
rect 10784 40384 10836 40390
rect 10784 40326 10836 40332
rect 10888 39370 10916 40394
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 10980 39914 11008 40326
rect 10968 39908 11020 39914
rect 10968 39850 11020 39856
rect 11060 39908 11112 39914
rect 11060 39850 11112 39856
rect 9864 39364 9916 39370
rect 9864 39306 9916 39312
rect 10876 39364 10928 39370
rect 10876 39306 10928 39312
rect 9876 39098 9904 39306
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 10888 38978 10916 39306
rect 10980 39098 11008 39850
rect 10968 39092 11020 39098
rect 10968 39034 11020 39040
rect 10888 38950 11008 38978
rect 10980 38894 11008 38950
rect 10968 38888 11020 38894
rect 10968 38830 11020 38836
rect 10876 38276 10928 38282
rect 10876 38218 10928 38224
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9968 38010 9996 38150
rect 9956 38004 10008 38010
rect 9956 37946 10008 37952
rect 10888 37330 10916 38218
rect 10980 37874 11008 38830
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 10876 37324 10928 37330
rect 10876 37266 10928 37272
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 9876 36310 9904 36654
rect 10704 36310 10732 37062
rect 10980 36786 11008 37810
rect 11072 37398 11100 39850
rect 11060 37392 11112 37398
rect 11060 37334 11112 37340
rect 11060 37120 11112 37126
rect 11060 37062 11112 37068
rect 10968 36780 11020 36786
rect 10968 36722 11020 36728
rect 11072 36582 11100 37062
rect 11060 36576 11112 36582
rect 11060 36518 11112 36524
rect 9864 36304 9916 36310
rect 9864 36246 9916 36252
rect 10692 36304 10744 36310
rect 10692 36246 10744 36252
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 11072 34678 11100 35022
rect 11060 34672 11112 34678
rect 11060 34614 11112 34620
rect 10784 34400 10836 34406
rect 10784 34342 10836 34348
rect 10796 34066 10824 34342
rect 10784 34060 10836 34066
rect 10784 34002 10836 34008
rect 9772 33380 9824 33386
rect 9772 33322 9824 33328
rect 9128 33108 9180 33114
rect 9128 33050 9180 33056
rect 9312 32836 9364 32842
rect 9312 32778 9364 32784
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 9140 31822 9168 32370
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 8772 31726 8984 31754
rect 8576 31340 8628 31346
rect 8576 31282 8628 31288
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 8312 30938 8340 31146
rect 8300 30932 8352 30938
rect 8300 30874 8352 30880
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 7800 30620 7880 30648
rect 7748 30602 7800 30608
rect 7852 30394 7880 30620
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7668 29838 7880 29866
rect 7944 29850 7972 30534
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 8036 29850 8064 30126
rect 7656 29640 7708 29646
rect 7576 29600 7656 29628
rect 7380 29582 7432 29588
rect 7708 29588 7788 29594
rect 7656 29582 7788 29588
rect 7668 29566 7788 29582
rect 7760 29306 7788 29566
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 7116 28150 7144 28698
rect 7208 28626 7236 29174
rect 7196 28620 7248 28626
rect 7196 28562 7248 28568
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 7196 28484 7248 28490
rect 7196 28426 7248 28432
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 7116 27334 7144 28086
rect 7208 28014 7236 28426
rect 7484 28422 7512 28562
rect 7760 28422 7788 29242
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 7484 28082 7512 28358
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7380 27872 7432 27878
rect 7380 27814 7432 27820
rect 7760 27826 7788 28358
rect 7852 28150 7880 29838
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8220 29646 8248 30670
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8680 29306 8708 31282
rect 8956 29714 8984 31726
rect 9036 31680 9088 31686
rect 9036 31622 9088 31628
rect 9048 31482 9076 31622
rect 9036 31476 9088 31482
rect 9036 31418 9088 31424
rect 9140 31346 9168 31758
rect 9324 31754 9352 32778
rect 9784 32366 9812 33322
rect 9772 32360 9824 32366
rect 9772 32302 9824 32308
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10980 32026 11008 32166
rect 11256 32026 11284 42094
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 11532 41138 11560 41958
rect 11808 41614 11836 42230
rect 11992 42022 12020 42638
rect 11980 42016 12032 42022
rect 11980 41958 12032 41964
rect 11992 41818 12020 41958
rect 11980 41812 12032 41818
rect 11980 41754 12032 41760
rect 11796 41608 11848 41614
rect 11796 41550 11848 41556
rect 11888 41608 11940 41614
rect 11888 41550 11940 41556
rect 11900 41274 11928 41550
rect 12084 41414 12112 43794
rect 12452 43314 12480 44814
rect 13452 44736 13504 44742
rect 13452 44678 13504 44684
rect 13464 44538 13492 44678
rect 13452 44532 13504 44538
rect 13452 44474 13504 44480
rect 12900 44328 12952 44334
rect 12900 44270 12952 44276
rect 13084 44328 13136 44334
rect 13084 44270 13136 44276
rect 12912 43994 12940 44270
rect 12900 43988 12952 43994
rect 12900 43930 12952 43936
rect 12532 43648 12584 43654
rect 12532 43590 12584 43596
rect 12544 43450 12572 43590
rect 12532 43444 12584 43450
rect 12532 43386 12584 43392
rect 12440 43308 12492 43314
rect 12440 43250 12492 43256
rect 12624 43240 12676 43246
rect 12624 43182 12676 43188
rect 12532 43104 12584 43110
rect 12532 43046 12584 43052
rect 12164 42152 12216 42158
rect 12164 42094 12216 42100
rect 12176 41818 12204 42094
rect 12164 41812 12216 41818
rect 12164 41754 12216 41760
rect 12544 41732 12572 43046
rect 12636 42906 12664 43182
rect 13096 43110 13124 44270
rect 14108 43994 14136 44814
rect 14648 44736 14700 44742
rect 14648 44678 14700 44684
rect 14660 44402 14688 44678
rect 15856 44538 15884 44814
rect 16040 44742 16068 44814
rect 16028 44736 16080 44742
rect 16028 44678 16080 44684
rect 15844 44532 15896 44538
rect 15844 44474 15896 44480
rect 14648 44396 14700 44402
rect 14648 44338 14700 44344
rect 14464 44192 14516 44198
rect 14464 44134 14516 44140
rect 14096 43988 14148 43994
rect 14096 43930 14148 43936
rect 14188 43920 14240 43926
rect 14188 43862 14240 43868
rect 13176 43784 13228 43790
rect 13176 43726 13228 43732
rect 13912 43784 13964 43790
rect 13912 43726 13964 43732
rect 13084 43104 13136 43110
rect 13084 43046 13136 43052
rect 12624 42900 12676 42906
rect 12624 42842 12676 42848
rect 11992 41386 12112 41414
rect 12452 41704 12572 41732
rect 11888 41268 11940 41274
rect 11888 41210 11940 41216
rect 11520 41132 11572 41138
rect 11520 41074 11572 41080
rect 11900 40390 11928 41210
rect 11888 40384 11940 40390
rect 11888 40326 11940 40332
rect 11888 39840 11940 39846
rect 11888 39782 11940 39788
rect 11900 39506 11928 39782
rect 11888 39500 11940 39506
rect 11888 39442 11940 39448
rect 11520 39296 11572 39302
rect 11520 39238 11572 39244
rect 11532 38962 11560 39238
rect 11520 38956 11572 38962
rect 11520 38898 11572 38904
rect 11336 38888 11388 38894
rect 11336 38830 11388 38836
rect 11348 37890 11376 38830
rect 11428 38344 11480 38350
rect 11428 38286 11480 38292
rect 11440 38010 11468 38286
rect 11428 38004 11480 38010
rect 11428 37946 11480 37952
rect 11348 37862 11468 37890
rect 11440 37330 11468 37862
rect 11428 37324 11480 37330
rect 11428 37266 11480 37272
rect 11336 34060 11388 34066
rect 11336 34002 11388 34008
rect 11348 32230 11376 34002
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 11348 32026 11376 32166
rect 10968 32020 11020 32026
rect 10968 31962 11020 31968
rect 11244 32020 11296 32026
rect 11244 31962 11296 31968
rect 11336 32020 11388 32026
rect 11336 31962 11388 31968
rect 11256 31822 11284 31962
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 9588 31748 9640 31754
rect 9588 31690 9640 31696
rect 9128 31340 9180 31346
rect 9128 31282 9180 31288
rect 9324 30258 9352 31690
rect 9600 31482 9628 31690
rect 9588 31476 9640 31482
rect 9588 31418 9640 31424
rect 10506 30832 10562 30841
rect 10506 30767 10562 30776
rect 10520 30734 10548 30767
rect 10508 30728 10560 30734
rect 10508 30670 10560 30676
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8852 29504 8904 29510
rect 8852 29446 8904 29452
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8760 28416 8812 28422
rect 8760 28358 8812 28364
rect 7840 28144 7892 28150
rect 7840 28086 7892 28092
rect 8772 28082 8800 28358
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 7840 27940 7892 27946
rect 7840 27882 7892 27888
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 7852 27826 7880 27882
rect 7392 27402 7420 27814
rect 7760 27798 7880 27826
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 7852 26042 7880 27798
rect 8220 27402 8248 27814
rect 8404 27674 8432 27882
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 8496 27062 8524 27814
rect 8484 27056 8536 27062
rect 8484 26998 8536 27004
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8588 26586 8616 26862
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7852 25294 7880 25978
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7944 25498 7972 25774
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7760 21350 7788 22510
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 8312 21010 8340 25094
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8128 19990 8156 20334
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7024 19446 7052 19654
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7024 17898 7052 19382
rect 6932 17870 7052 17898
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6472 17338 6500 17546
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6564 16998 6592 17546
rect 6932 17202 6960 17870
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7024 17134 7052 17682
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 16182 6592 16934
rect 6828 16516 6880 16522
rect 6828 16458 6880 16464
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6748 15162 6776 15438
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 5736 12850 5764 14214
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5828 12850 5856 13330
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12730 5856 12786
rect 5644 12702 5856 12730
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5644 12102 5672 12702
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11694 5672 12038
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 9178 2544 9522
rect 4632 9450 4660 10406
rect 4724 10266 4752 10542
rect 5644 10470 5672 11630
rect 5724 10668 5776 10674
rect 5920 10656 5948 13262
rect 6012 12986 6040 13262
rect 6748 13258 6776 13670
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 5776 10628 5948 10656
rect 5724 10610 5776 10616
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9722 5212 9998
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5736 9654 5764 10610
rect 6748 10606 6776 12718
rect 6840 12170 6868 16458
rect 7024 16454 7052 17070
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 15570 7052 16390
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7208 13938 7236 19926
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7392 18426 7420 19110
rect 7852 18630 7880 19654
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7944 18970 7972 19246
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7668 17746 7696 18566
rect 7852 18222 7880 18566
rect 8312 18290 8340 18770
rect 8496 18358 8524 19314
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8036 17270 8064 17478
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8680 16046 8708 17478
rect 8864 16674 8892 29446
rect 9508 29306 9536 30194
rect 10416 29776 10468 29782
rect 10416 29718 10468 29724
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9232 28762 9260 29106
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9036 28620 9088 28626
rect 9036 28562 9088 28568
rect 9048 28218 9076 28562
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 9324 27470 9352 29038
rect 10428 28762 10456 29718
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 11072 29306 11100 29582
rect 11256 29510 11284 31758
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 11060 29300 11112 29306
rect 11060 29242 11112 29248
rect 10416 28756 10468 28762
rect 10416 28698 10468 28704
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9600 28218 9628 28358
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9404 28144 9456 28150
rect 9404 28086 9456 28092
rect 9312 27464 9364 27470
rect 9312 27406 9364 27412
rect 9416 26518 9444 28086
rect 9496 28076 9548 28082
rect 9680 28076 9732 28082
rect 9548 28036 9680 28064
rect 9496 28018 9548 28024
rect 9680 28018 9732 28024
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 9404 26512 9456 26518
rect 9404 26454 9456 26460
rect 9508 26382 9536 28018
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9600 26926 9628 27338
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9048 25906 9076 26318
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9508 25838 9536 26318
rect 9600 25974 9628 26862
rect 9692 26586 9720 27406
rect 10336 27130 10364 28018
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 11164 27674 11192 27814
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 11440 26926 11468 37266
rect 11532 34610 11560 38898
rect 11992 38894 12020 41386
rect 12256 40520 12308 40526
rect 12256 40462 12308 40468
rect 12268 40186 12296 40462
rect 12256 40180 12308 40186
rect 12256 40122 12308 40128
rect 12072 39976 12124 39982
rect 12072 39918 12124 39924
rect 12084 39098 12112 39918
rect 12072 39092 12124 39098
rect 12072 39034 12124 39040
rect 11980 38888 12032 38894
rect 11980 38830 12032 38836
rect 12452 38570 12480 41704
rect 12636 41614 12664 42842
rect 13096 42158 13124 43046
rect 13188 42906 13216 43726
rect 13820 43648 13872 43654
rect 13820 43590 13872 43596
rect 13176 42900 13228 42906
rect 13176 42842 13228 42848
rect 13832 42702 13860 43590
rect 13924 43450 13952 43726
rect 13912 43444 13964 43450
rect 13912 43386 13964 43392
rect 13910 42800 13966 42809
rect 13910 42735 13966 42744
rect 13924 42702 13952 42735
rect 13820 42696 13872 42702
rect 13820 42638 13872 42644
rect 13912 42696 13964 42702
rect 13912 42638 13964 42644
rect 14004 42696 14056 42702
rect 14004 42638 14056 42644
rect 13268 42288 13320 42294
rect 13268 42230 13320 42236
rect 13084 42152 13136 42158
rect 13084 42094 13136 42100
rect 12900 41676 12952 41682
rect 12900 41618 12952 41624
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 12532 41540 12584 41546
rect 12532 41482 12584 41488
rect 12544 40458 12572 41482
rect 12912 40526 12940 41618
rect 13280 41546 13308 42230
rect 13360 42152 13412 42158
rect 13360 42094 13412 42100
rect 13372 41818 13400 42094
rect 14016 42022 14044 42638
rect 14096 42560 14148 42566
rect 14096 42502 14148 42508
rect 14108 42158 14136 42502
rect 14096 42152 14148 42158
rect 14096 42094 14148 42100
rect 14004 42016 14056 42022
rect 14004 41958 14056 41964
rect 13360 41812 13412 41818
rect 13360 41754 13412 41760
rect 13268 41540 13320 41546
rect 13268 41482 13320 41488
rect 14016 41070 14044 41958
rect 14004 41064 14056 41070
rect 14004 41006 14056 41012
rect 13728 40928 13780 40934
rect 13728 40870 13780 40876
rect 12900 40520 12952 40526
rect 12900 40462 12952 40468
rect 13544 40520 13596 40526
rect 13544 40462 13596 40468
rect 12532 40452 12584 40458
rect 12532 40394 12584 40400
rect 12544 39030 12572 40394
rect 12808 39976 12860 39982
rect 12808 39918 12860 39924
rect 12624 39296 12676 39302
rect 12624 39238 12676 39244
rect 12532 39024 12584 39030
rect 12532 38966 12584 38972
rect 12360 38542 12480 38570
rect 12256 37256 12308 37262
rect 12256 37198 12308 37204
rect 12268 36922 12296 37198
rect 12256 36916 12308 36922
rect 12256 36858 12308 36864
rect 12164 36712 12216 36718
rect 12164 36654 12216 36660
rect 12072 36576 12124 36582
rect 12072 36518 12124 36524
rect 12084 35698 12112 36518
rect 12176 36106 12204 36654
rect 12164 36100 12216 36106
rect 12164 36042 12216 36048
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12256 35148 12308 35154
rect 12256 35090 12308 35096
rect 12268 34950 12296 35090
rect 12256 34944 12308 34950
rect 12256 34886 12308 34892
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 11612 34400 11664 34406
rect 11612 34342 11664 34348
rect 11624 33998 11652 34342
rect 12360 34184 12388 38542
rect 12544 38350 12572 38966
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12636 36786 12664 39238
rect 12820 39098 12848 39918
rect 12808 39092 12860 39098
rect 12808 39034 12860 39040
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12728 38486 12756 38898
rect 12912 38758 12940 40462
rect 13360 39840 13412 39846
rect 13360 39782 13412 39788
rect 13372 39098 13400 39782
rect 13556 39642 13584 40462
rect 13740 40186 13768 40870
rect 13728 40180 13780 40186
rect 13728 40122 13780 40128
rect 14016 39846 14044 41006
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 13544 39636 13596 39642
rect 13544 39578 13596 39584
rect 13360 39092 13412 39098
rect 13360 39034 13412 39040
rect 12900 38752 12952 38758
rect 12900 38694 12952 38700
rect 12716 38480 12768 38486
rect 12716 38422 12768 38428
rect 13372 38350 13400 39034
rect 13556 38894 13584 39578
rect 14016 39438 14044 39782
rect 14004 39432 14056 39438
rect 14004 39374 14056 39380
rect 14016 39030 14044 39374
rect 14004 39024 14056 39030
rect 14004 38966 14056 38972
rect 13544 38888 13596 38894
rect 13544 38830 13596 38836
rect 13728 38752 13780 38758
rect 13728 38694 13780 38700
rect 13740 38350 13768 38694
rect 12900 38344 12952 38350
rect 12900 38286 12952 38292
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 12912 37874 12940 38286
rect 13740 38010 13768 38286
rect 13728 38004 13780 38010
rect 13728 37946 13780 37952
rect 12900 37868 12952 37874
rect 12900 37810 12952 37816
rect 13360 37868 13412 37874
rect 13360 37810 13412 37816
rect 12912 37194 12940 37810
rect 12992 37664 13044 37670
rect 12992 37606 13044 37612
rect 13004 37330 13032 37606
rect 12992 37324 13044 37330
rect 12992 37266 13044 37272
rect 13372 37262 13400 37810
rect 14016 37806 14044 38966
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 12900 37188 12952 37194
rect 12900 37130 12952 37136
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12452 35834 12480 35974
rect 12440 35828 12492 35834
rect 12440 35770 12492 35776
rect 12636 35086 12664 36722
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 12808 35488 12860 35494
rect 12808 35430 12860 35436
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 12268 34156 12388 34184
rect 12268 33998 12296 34156
rect 12348 34060 12400 34066
rect 12348 34002 12400 34008
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 11808 33862 11836 33934
rect 11980 33924 12032 33930
rect 11980 33866 12032 33872
rect 11796 33856 11848 33862
rect 11796 33798 11848 33804
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11624 32434 11652 33458
rect 11704 32768 11756 32774
rect 11704 32710 11756 32716
rect 11716 32434 11744 32710
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11704 32428 11756 32434
rect 11704 32370 11756 32376
rect 11624 30138 11652 32370
rect 11808 31754 11836 33798
rect 11992 33658 12020 33866
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 11886 33552 11942 33561
rect 12084 33538 12112 33934
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 11992 33522 12112 33538
rect 11886 33487 11888 33496
rect 11940 33487 11942 33496
rect 11980 33516 12112 33522
rect 11888 33458 11940 33464
rect 12032 33510 12112 33516
rect 11980 33458 12032 33464
rect 12176 33386 12204 33798
rect 12268 33522 12296 33798
rect 12360 33674 12388 34002
rect 12544 33998 12572 34546
rect 12636 34134 12664 34614
rect 12820 34610 12848 35430
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 13084 34604 13136 34610
rect 13084 34546 13136 34552
rect 12728 34202 12756 34546
rect 12716 34196 12768 34202
rect 12716 34138 12768 34144
rect 12624 34128 12676 34134
rect 12624 34070 12676 34076
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12440 33856 12492 33862
rect 12440 33798 12492 33804
rect 12452 33674 12480 33798
rect 12360 33646 12480 33674
rect 12256 33516 12308 33522
rect 12256 33458 12308 33464
rect 12164 33380 12216 33386
rect 12164 33322 12216 33328
rect 12072 33312 12124 33318
rect 12072 33254 12124 33260
rect 12084 33114 12112 33254
rect 12268 33130 12296 33458
rect 12452 33386 12480 33646
rect 12440 33380 12492 33386
rect 12440 33322 12492 33328
rect 12072 33108 12124 33114
rect 12268 33102 12480 33130
rect 12072 33050 12124 33056
rect 12452 32978 12480 33102
rect 12440 32972 12492 32978
rect 12440 32914 12492 32920
rect 12544 32858 12572 33934
rect 12728 33658 12756 34138
rect 12820 33930 12848 34546
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 12900 34196 12952 34202
rect 12900 34138 12952 34144
rect 12808 33924 12860 33930
rect 12808 33866 12860 33872
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 12624 33516 12676 33522
rect 12912 33504 12940 34138
rect 13004 34066 13032 34342
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 13004 33522 13032 34002
rect 13096 33930 13124 34546
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13084 33924 13136 33930
rect 13084 33866 13136 33872
rect 12676 33476 12940 33504
rect 12992 33516 13044 33522
rect 12624 33458 12676 33464
rect 12992 33458 13044 33464
rect 13096 33402 13124 33866
rect 13004 33374 13124 33402
rect 12900 33312 12952 33318
rect 12900 33254 12952 33260
rect 12624 33108 12676 33114
rect 12624 33050 12676 33056
rect 12452 32830 12572 32858
rect 12452 31822 12480 32830
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 11808 31726 11928 31754
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11716 30734 11744 31622
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 11624 30110 11744 30138
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11624 29646 11652 29990
rect 11520 29640 11572 29646
rect 11520 29582 11572 29588
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11532 28762 11560 29582
rect 11520 28756 11572 28762
rect 11520 28698 11572 28704
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11624 28150 11652 28494
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 25498 9168 25638
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 9508 25362 9536 25774
rect 9600 25498 9628 25910
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9692 25362 9720 26522
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 9784 26042 9812 26250
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 10612 25906 10640 26250
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10704 25498 10732 25638
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 11072 25362 11100 25774
rect 11716 25362 11744 30110
rect 11808 29646 11836 31282
rect 11900 31226 11928 31726
rect 11980 31748 12032 31754
rect 11980 31690 12032 31696
rect 11992 31482 12020 31690
rect 11980 31476 12032 31482
rect 11980 31418 12032 31424
rect 11900 31198 12020 31226
rect 11992 30598 12020 31198
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29646 11928 29990
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 9496 25356 9548 25362
rect 9496 25298 9548 25304
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 11072 24274 11100 25298
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11348 24750 11376 25162
rect 11716 24954 11744 25298
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11808 23118 11836 29582
rect 11992 28558 12020 30534
rect 12084 30394 12112 30670
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 12176 30326 12204 31758
rect 12346 30696 12402 30705
rect 12346 30631 12402 30640
rect 12440 30660 12492 30666
rect 12360 30598 12388 30631
rect 12440 30602 12492 30608
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12164 30320 12216 30326
rect 12164 30262 12216 30268
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 12268 28506 12296 30126
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11900 23866 11928 24074
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11992 23746 12020 28494
rect 12268 28478 12388 28506
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 12256 28416 12308 28422
rect 12256 28358 12308 28364
rect 12084 28150 12112 28358
rect 12268 28218 12296 28358
rect 12256 28212 12308 28218
rect 12256 28154 12308 28160
rect 12072 28144 12124 28150
rect 12072 28086 12124 28092
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12084 26042 12112 26182
rect 12072 26036 12124 26042
rect 12072 25978 12124 25984
rect 12360 25838 12388 28478
rect 12452 28218 12480 30602
rect 12544 29850 12572 31894
rect 12636 31346 12664 33050
rect 12912 32910 12940 33254
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 13004 31754 13032 33374
rect 13188 33318 13216 33934
rect 13280 33386 13308 36314
rect 13372 35834 13400 37198
rect 13452 37120 13504 37126
rect 13452 37062 13504 37068
rect 13636 37120 13688 37126
rect 13636 37062 13688 37068
rect 13464 36922 13492 37062
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13452 36032 13504 36038
rect 13452 35974 13504 35980
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13464 34746 13492 35974
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13360 34536 13412 34542
rect 13360 34478 13412 34484
rect 13268 33380 13320 33386
rect 13268 33322 13320 33328
rect 13176 33312 13228 33318
rect 13176 33254 13228 33260
rect 12820 31726 13032 31754
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12820 30274 12848 31726
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 13188 30870 13216 31214
rect 13084 30864 13136 30870
rect 13084 30806 13136 30812
rect 13176 30864 13228 30870
rect 13176 30806 13228 30812
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12912 30394 12940 30670
rect 12992 30592 13044 30598
rect 12990 30560 12992 30569
rect 13044 30560 13046 30569
rect 12990 30495 13046 30504
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12990 30288 13046 30297
rect 12728 30258 12940 30274
rect 12716 30252 12940 30258
rect 12768 30246 12940 30252
rect 12716 30194 12768 30200
rect 12624 30116 12676 30122
rect 12624 30058 12676 30064
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12636 29646 12664 30058
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12440 27396 12492 27402
rect 12440 27338 12492 27344
rect 12452 27062 12480 27338
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 12452 25974 12480 26998
rect 12544 26518 12572 27950
rect 12636 27538 12664 28018
rect 12820 27674 12848 28494
rect 12808 27668 12860 27674
rect 12808 27610 12860 27616
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 12532 26512 12584 26518
rect 12532 26454 12584 26460
rect 12636 26450 12664 27474
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12452 25294 12480 25910
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12452 24138 12480 25230
rect 12912 24410 12940 30246
rect 12990 30223 12992 30232
rect 13044 30223 13046 30232
rect 12992 30194 13044 30200
rect 12992 29504 13044 29510
rect 12992 29446 13044 29452
rect 13004 28082 13032 29446
rect 13096 29238 13124 30806
rect 13188 30326 13216 30806
rect 13176 30320 13228 30326
rect 13176 30262 13228 30268
rect 13084 29232 13136 29238
rect 13084 29174 13136 29180
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 13004 27554 13032 27814
rect 13096 27674 13124 28018
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 13004 27526 13124 27554
rect 13096 27470 13124 27526
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12440 24132 12492 24138
rect 12440 24074 12492 24080
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 11900 23718 12020 23746
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 22778 10088 22918
rect 10520 22778 10548 23054
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10612 22234 10640 22918
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10888 21978 10916 22578
rect 11152 22092 11204 22098
rect 11440 22094 11468 22918
rect 11808 22234 11836 23054
rect 11900 22642 11928 23718
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11796 22228 11848 22234
rect 11796 22170 11848 22176
rect 11152 22034 11204 22040
rect 11256 22066 11468 22094
rect 10888 21962 11008 21978
rect 10876 21956 11008 21962
rect 10928 21950 11008 21956
rect 10876 21898 10928 21904
rect 10980 21842 11008 21950
rect 11060 21888 11112 21894
rect 10980 21836 11060 21842
rect 10980 21830 11112 21836
rect 10980 21814 11100 21830
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9508 19378 9536 19858
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9508 18970 9536 19314
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18426 9260 18702
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9048 17610 9076 18294
rect 9508 17882 9536 18906
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9048 17354 9076 17546
rect 8956 17338 9076 17354
rect 8944 17332 9076 17338
rect 8996 17326 9076 17332
rect 8944 17274 8996 17280
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8956 16794 8984 17070
rect 9048 16794 9076 17326
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8864 16646 9076 16674
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8312 15570 8340 15982
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15026 8340 15506
rect 9048 15094 9076 16646
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9324 16182 9352 16526
rect 9600 16250 9628 20742
rect 10520 19334 10548 21490
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10612 20058 10640 20198
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10980 19786 11008 21814
rect 11164 19922 11192 22034
rect 11256 20330 11284 22066
rect 11992 20602 12020 22510
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12268 21894 12296 22034
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12452 21690 12480 21898
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10980 19666 11008 19722
rect 11152 19712 11204 19718
rect 10980 19660 11152 19666
rect 10980 19654 11204 19660
rect 10980 19638 11192 19654
rect 11072 19378 11100 19638
rect 11256 19514 11284 20266
rect 11992 20058 12020 20538
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11060 19372 11112 19378
rect 10140 19304 10192 19310
rect 10520 19306 10732 19334
rect 11060 19314 11112 19320
rect 10140 19246 10192 19252
rect 10152 18426 10180 19246
rect 10704 18766 10732 19306
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10336 17338 10364 17546
rect 10704 17490 10732 18702
rect 10796 18426 10824 18838
rect 10888 18426 10916 18906
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17610 10824 18022
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10704 17462 10824 17490
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10612 16794 10640 16934
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9680 16176 9732 16182
rect 10796 16153 10824 17462
rect 9680 16118 9732 16124
rect 10782 16144 10838 16153
rect 9692 15094 9720 16118
rect 10782 16079 10838 16088
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10520 15162 10548 15370
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 6932 12850 6960 13126
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 1768 9036 1820 9042
rect 1820 8996 1992 9024
rect 1768 8978 1820 8984
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1964 6866 1992 8996
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 2650 2084 6802
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6458 3188 6598
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 4816 6390 4844 9590
rect 6748 9042 6776 10542
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8090 6776 8978
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6748 7342 6776 8026
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 4804 6384 4856 6390
rect 4802 6352 4804 6361
rect 4856 6352 4858 6361
rect 4802 6287 4858 6296
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 6840 5710 6868 12106
rect 7208 10674 7236 13126
rect 7300 12782 7328 14010
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7668 13530 7696 13874
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7944 13394 7972 14486
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7668 12102 7696 12786
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7116 8906 7144 10610
rect 7300 10606 7328 11018
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7392 9042 7420 11086
rect 7484 10810 7512 11086
rect 7668 11082 7696 12038
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7852 11354 7880 11630
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7944 11150 7972 13330
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8128 12782 8156 13126
rect 8588 12782 8616 13126
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7484 10606 7512 10746
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7392 8922 7420 8978
rect 7104 8900 7156 8906
rect 7392 8894 7512 8922
rect 7104 8842 7156 8848
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 5914 6960 7142
rect 7116 6798 7144 7890
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7546 7236 7822
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5166 6592 5510
rect 7208 5370 7236 7482
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6730 7328 7346
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7392 6254 7420 8366
rect 7484 7342 7512 8894
rect 7760 7546 7788 10406
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8498 7972 8774
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7484 6866 7512 7278
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 8220 6798 8248 7210
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7668 6254 7696 6598
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 7852 4622 7880 6598
rect 8208 6384 8260 6390
rect 8206 6352 8208 6361
rect 8312 6372 8340 8366
rect 8260 6352 8340 6372
rect 8262 6344 8340 6352
rect 8206 6287 8262 6296
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5574 8156 6054
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5030 8156 5510
rect 8220 5234 8248 6287
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4078 7236 4422
rect 8128 4078 8156 4966
rect 8220 4214 8248 5170
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8128 3058 8156 4014
rect 8220 3738 8248 4150
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8772 3126 8800 14826
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 12918 9628 13670
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9600 11762 9628 12854
rect 10152 12782 10180 13126
rect 10232 12912 10284 12918
rect 10336 12900 10364 13398
rect 10284 12872 10364 12900
rect 10232 12854 10284 12860
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10336 12442 10364 12872
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9600 10606 9628 11698
rect 9692 11150 9720 11698
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9680 9104 9732 9110
rect 9784 9092 9812 12106
rect 9968 11880 9996 12106
rect 10336 12102 10364 12378
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10046 11928 10102 11937
rect 9968 11872 10046 11880
rect 9968 11852 10048 11872
rect 9862 11248 9918 11257
rect 9862 11183 9864 11192
rect 9916 11183 9918 11192
rect 9864 11154 9916 11160
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10062 9904 10950
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9732 9064 9812 9092
rect 9680 9046 9732 9052
rect 9784 8906 9812 9064
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9784 6730 9812 8842
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9876 6474 9904 9998
rect 9968 8294 9996 11852
rect 10100 11863 10102 11872
rect 10048 11834 10100 11840
rect 10428 11762 10456 12038
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 10060 10130 10088 11319
rect 10336 10996 10364 11698
rect 10416 11008 10468 11014
rect 10336 10976 10416 10996
rect 10508 11008 10560 11014
rect 10468 10976 10470 10985
rect 10336 10968 10414 10976
rect 10508 10950 10560 10956
rect 10414 10911 10470 10920
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10060 9110 10088 10066
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7546 9996 7686
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10060 7478 10088 8910
rect 10152 8634 10180 9454
rect 10244 8634 10272 9658
rect 10336 9586 10364 9862
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9178 10456 9454
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10520 9042 10548 10950
rect 10612 9178 10640 12174
rect 10704 11898 10732 12854
rect 10796 12374 10824 16079
rect 11072 15434 11100 19314
rect 11256 18630 11284 19450
rect 12084 19446 12112 20334
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11624 18834 11652 19382
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 16250 11744 16458
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11808 15706 11836 18158
rect 11900 17882 11928 18634
rect 12360 18426 12388 20402
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11900 17338 11928 17818
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 13802 11652 14350
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10980 12714 11008 12786
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10888 11898 10916 12378
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10704 10538 10732 11698
rect 10784 11688 10836 11694
rect 10836 11648 10916 11676
rect 10784 11630 10836 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11234 10824 11494
rect 10888 11393 10916 11648
rect 10874 11384 10930 11393
rect 10980 11354 11008 12650
rect 11072 11558 11100 12786
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10874 11319 10930 11328
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10796 11206 10916 11234
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10538 10824 11086
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10796 10062 10824 10474
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9178 10732 9930
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10782 9072 10838 9081
rect 10508 9036 10560 9042
rect 10782 9007 10784 9016
rect 10508 8978 10560 8984
rect 10836 9007 10838 9016
rect 10784 8978 10836 8984
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10152 7886 10180 8434
rect 10336 7970 10364 8502
rect 10244 7942 10364 7970
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10244 7018 10272 7942
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10152 6990 10272 7018
rect 9876 6446 9996 6474
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9140 4146 9168 5170
rect 9692 4622 9720 5170
rect 9876 4622 9904 6258
rect 9968 5370 9996 6446
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4622 10088 5102
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9692 4078 9720 4558
rect 9876 4214 9904 4558
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9324 3126 9352 3674
rect 9692 3534 9720 4014
rect 9876 3738 9904 4150
rect 10152 4146 10180 6990
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6254 10272 6734
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5234 10272 6190
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9508 3194 9536 3470
rect 10244 3398 10272 5170
rect 10336 5030 10364 7822
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10428 4321 10456 8842
rect 10520 8498 10548 8842
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10520 7274 10548 7822
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10520 6984 10548 7210
rect 10612 7177 10640 7346
rect 10704 7206 10732 7822
rect 10888 7410 10916 11206
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10980 10266 11008 11086
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10692 7200 10744 7206
rect 10598 7168 10654 7177
rect 10692 7142 10744 7148
rect 10598 7103 10654 7112
rect 10888 7002 10916 7346
rect 10876 6996 10928 7002
rect 10520 6956 10640 6984
rect 10506 6896 10562 6905
rect 10506 6831 10562 6840
rect 10520 6798 10548 6831
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10520 4622 10548 5306
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10414 4312 10470 4321
rect 10414 4247 10470 4256
rect 10428 4078 10456 4247
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10612 3942 10640 6956
rect 10876 6938 10928 6944
rect 10980 6798 11008 9386
rect 11072 8022 11100 9998
rect 11164 9654 11192 13670
rect 11624 13394 11652 13738
rect 11992 13530 12020 17070
rect 12360 15502 12388 18362
rect 12452 18290 12480 18566
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12452 17814 12480 18226
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12452 17134 12480 17750
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 16794 12480 17070
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12452 16114 12480 16730
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12084 15162 12112 15302
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 13870 12296 14758
rect 12452 14074 12480 15302
rect 12636 14414 12664 24006
rect 12912 23866 12940 24346
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 13004 23662 13032 24686
rect 13096 24342 13124 27406
rect 13280 26586 13308 33322
rect 13372 32910 13400 34478
rect 13452 33992 13504 33998
rect 13452 33934 13504 33940
rect 13464 33561 13492 33934
rect 13450 33552 13506 33561
rect 13450 33487 13506 33496
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13544 30864 13596 30870
rect 13544 30806 13596 30812
rect 13556 30734 13584 30806
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 13372 30297 13400 30534
rect 13648 30394 13676 37062
rect 14016 36786 14044 37742
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 14016 36242 14044 36722
rect 14004 36236 14056 36242
rect 14004 36178 14056 36184
rect 14096 36032 14148 36038
rect 14096 35974 14148 35980
rect 14108 35834 14136 35974
rect 14096 35828 14148 35834
rect 14096 35770 14148 35776
rect 14200 33998 14228 43862
rect 14476 43790 14504 44134
rect 14464 43784 14516 43790
rect 14464 43726 14516 43732
rect 14660 43314 14688 44338
rect 14924 44328 14976 44334
rect 14924 44270 14976 44276
rect 14936 43790 14964 44270
rect 16132 43858 16160 44814
rect 16856 44804 16908 44810
rect 16856 44746 16908 44752
rect 16120 43852 16172 43858
rect 16120 43794 16172 43800
rect 14924 43784 14976 43790
rect 14924 43726 14976 43732
rect 15568 43716 15620 43722
rect 15568 43658 15620 43664
rect 15580 43450 15608 43658
rect 15568 43444 15620 43450
rect 15568 43386 15620 43392
rect 16132 43314 16160 43794
rect 16868 43790 16896 44746
rect 17868 44736 17920 44742
rect 17868 44678 17920 44684
rect 19156 44736 19208 44742
rect 19156 44678 19208 44684
rect 19984 44736 20036 44742
rect 19984 44678 20036 44684
rect 17880 44402 17908 44678
rect 19168 44402 19196 44678
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19996 44538 20024 44678
rect 19984 44532 20036 44538
rect 19984 44474 20036 44480
rect 20076 44464 20128 44470
rect 20076 44406 20128 44412
rect 20628 44464 20680 44470
rect 20628 44406 20680 44412
rect 17868 44396 17920 44402
rect 17868 44338 17920 44344
rect 18512 44396 18564 44402
rect 18512 44338 18564 44344
rect 19156 44396 19208 44402
rect 19156 44338 19208 44344
rect 17132 44328 17184 44334
rect 17132 44270 17184 44276
rect 17316 44328 17368 44334
rect 17316 44270 17368 44276
rect 17144 43994 17172 44270
rect 17132 43988 17184 43994
rect 17132 43930 17184 43936
rect 17328 43926 17356 44270
rect 17776 43988 17828 43994
rect 17776 43930 17828 43936
rect 17316 43920 17368 43926
rect 17316 43862 17368 43868
rect 16856 43784 16908 43790
rect 16856 43726 16908 43732
rect 14648 43308 14700 43314
rect 14648 43250 14700 43256
rect 16120 43308 16172 43314
rect 16120 43250 16172 43256
rect 14462 42800 14518 42809
rect 14660 42770 14688 43250
rect 14832 43240 14884 43246
rect 14832 43182 14884 43188
rect 14462 42735 14518 42744
rect 14556 42764 14608 42770
rect 14476 42090 14504 42735
rect 14556 42706 14608 42712
rect 14648 42764 14700 42770
rect 14648 42706 14700 42712
rect 14568 42090 14596 42706
rect 14660 42294 14688 42706
rect 14844 42362 14872 43182
rect 15016 43104 15068 43110
rect 15016 43046 15068 43052
rect 16764 43104 16816 43110
rect 16764 43046 16816 43052
rect 14924 42560 14976 42566
rect 14924 42502 14976 42508
rect 14832 42356 14884 42362
rect 14832 42298 14884 42304
rect 14648 42288 14700 42294
rect 14648 42230 14700 42236
rect 14936 42226 14964 42502
rect 15028 42226 15056 43046
rect 15200 42628 15252 42634
rect 15200 42570 15252 42576
rect 15212 42362 15240 42570
rect 15200 42356 15252 42362
rect 15200 42298 15252 42304
rect 16672 42356 16724 42362
rect 16672 42298 16724 42304
rect 14924 42220 14976 42226
rect 14924 42162 14976 42168
rect 15016 42220 15068 42226
rect 15016 42162 15068 42168
rect 15568 42220 15620 42226
rect 15568 42162 15620 42168
rect 14464 42084 14516 42090
rect 14464 42026 14516 42032
rect 14556 42084 14608 42090
rect 14556 42026 14608 42032
rect 15028 41546 15056 42162
rect 15580 41818 15608 42162
rect 15568 41812 15620 41818
rect 15568 41754 15620 41760
rect 16684 41614 16712 42298
rect 16776 42294 16804 43046
rect 16868 42702 16896 43726
rect 17788 43450 17816 43930
rect 17776 43444 17828 43450
rect 17776 43386 17828 43392
rect 17684 43308 17736 43314
rect 17684 43250 17736 43256
rect 17316 43240 17368 43246
rect 17316 43182 17368 43188
rect 17224 43104 17276 43110
rect 17224 43046 17276 43052
rect 17236 42838 17264 43046
rect 17328 42906 17356 43182
rect 17316 42900 17368 42906
rect 17316 42842 17368 42848
rect 17224 42832 17276 42838
rect 17224 42774 17276 42780
rect 16856 42696 16908 42702
rect 16856 42638 16908 42644
rect 16764 42288 16816 42294
rect 16764 42230 16816 42236
rect 16776 41614 16804 42230
rect 15476 41608 15528 41614
rect 15476 41550 15528 41556
rect 16672 41608 16724 41614
rect 16672 41550 16724 41556
rect 16764 41608 16816 41614
rect 16764 41550 16816 41556
rect 15016 41540 15068 41546
rect 15016 41482 15068 41488
rect 15488 41070 15516 41550
rect 16868 41414 16896 42638
rect 17040 42560 17092 42566
rect 17040 42502 17092 42508
rect 17052 41614 17080 42502
rect 17696 42362 17724 43250
rect 17684 42356 17736 42362
rect 17684 42298 17736 42304
rect 17408 42220 17460 42226
rect 17408 42162 17460 42168
rect 17316 42152 17368 42158
rect 17316 42094 17368 42100
rect 17328 41818 17356 42094
rect 17316 41812 17368 41818
rect 17316 41754 17368 41760
rect 17040 41608 17092 41614
rect 17040 41550 17092 41556
rect 17316 41472 17368 41478
rect 17420 41460 17448 42162
rect 17592 41608 17644 41614
rect 17592 41550 17644 41556
rect 17368 41432 17448 41460
rect 17316 41414 17368 41420
rect 16684 41386 16896 41414
rect 14280 41064 14332 41070
rect 14280 41006 14332 41012
rect 15476 41064 15528 41070
rect 15476 41006 15528 41012
rect 15568 41064 15620 41070
rect 15568 41006 15620 41012
rect 14292 40730 14320 41006
rect 14280 40724 14332 40730
rect 14280 40666 14332 40672
rect 15108 40520 15160 40526
rect 15108 40462 15160 40468
rect 15120 39846 15148 40462
rect 15488 40050 15516 41006
rect 15476 40044 15528 40050
rect 15476 39986 15528 39992
rect 15108 39840 15160 39846
rect 15108 39782 15160 39788
rect 15292 39092 15344 39098
rect 15292 39034 15344 39040
rect 14740 38888 14792 38894
rect 14740 38830 14792 38836
rect 14752 38554 14780 38830
rect 14740 38548 14792 38554
rect 14740 38490 14792 38496
rect 15304 38282 15332 39034
rect 15292 38276 15344 38282
rect 15292 38218 15344 38224
rect 15304 37942 15332 38218
rect 15292 37936 15344 37942
rect 15292 37878 15344 37884
rect 15292 37800 15344 37806
rect 15292 37742 15344 37748
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 15212 36922 15240 37062
rect 15304 36922 15332 37742
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15292 36916 15344 36922
rect 15292 36858 15344 36864
rect 15200 36100 15252 36106
rect 15200 36042 15252 36048
rect 15212 35834 15240 36042
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15580 35290 15608 41006
rect 16120 40928 16172 40934
rect 16120 40870 16172 40876
rect 16132 40594 16160 40870
rect 16120 40588 16172 40594
rect 16120 40530 16172 40536
rect 16684 40526 16712 41386
rect 16672 40520 16724 40526
rect 16672 40462 16724 40468
rect 16028 40452 16080 40458
rect 16028 40394 16080 40400
rect 16856 40452 16908 40458
rect 16856 40394 16908 40400
rect 15752 39840 15804 39846
rect 15752 39782 15804 39788
rect 15764 39642 15792 39782
rect 15752 39636 15804 39642
rect 15752 39578 15804 39584
rect 16040 39370 16068 40394
rect 16868 40118 16896 40394
rect 17224 40384 17276 40390
rect 17224 40326 17276 40332
rect 17236 40118 17264 40326
rect 16856 40112 16908 40118
rect 16856 40054 16908 40060
rect 17224 40112 17276 40118
rect 17224 40054 17276 40060
rect 16120 39976 16172 39982
rect 16120 39918 16172 39924
rect 16212 39976 16264 39982
rect 16212 39918 16264 39924
rect 16132 39506 16160 39918
rect 16120 39500 16172 39506
rect 16120 39442 16172 39448
rect 16028 39364 16080 39370
rect 16028 39306 16080 39312
rect 16028 37664 16080 37670
rect 16028 37606 16080 37612
rect 16040 37330 16068 37606
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 16132 37210 16160 39442
rect 16040 37194 16160 37210
rect 16028 37188 16160 37194
rect 16080 37182 16160 37188
rect 16028 37130 16080 37136
rect 16040 36854 16068 37130
rect 16028 36848 16080 36854
rect 16028 36790 16080 36796
rect 15936 35760 15988 35766
rect 15936 35702 15988 35708
rect 14280 35284 14332 35290
rect 14280 35226 14332 35232
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 13820 33856 13872 33862
rect 13820 33798 13872 33804
rect 13832 33658 13860 33798
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13820 33312 13872 33318
rect 13820 33254 13872 33260
rect 13832 33046 13860 33254
rect 13820 33040 13872 33046
rect 13820 32982 13872 32988
rect 14200 32910 14228 33934
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14004 31476 14056 31482
rect 14004 31418 14056 31424
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30394 13768 31214
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13832 30938 13860 31078
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13636 30388 13688 30394
rect 13636 30330 13688 30336
rect 13728 30388 13780 30394
rect 13728 30330 13780 30336
rect 13358 30288 13414 30297
rect 13832 30274 13860 30670
rect 13912 30592 13964 30598
rect 13910 30560 13912 30569
rect 13964 30560 13966 30569
rect 13910 30495 13966 30504
rect 13358 30223 13414 30232
rect 13740 30246 13860 30274
rect 13360 30048 13412 30054
rect 13360 29990 13412 29996
rect 13372 29850 13400 29990
rect 13360 29844 13412 29850
rect 13360 29786 13412 29792
rect 13740 29238 13768 30246
rect 14016 30190 14044 31418
rect 14292 31346 14320 35226
rect 14832 34944 14884 34950
rect 14832 34886 14884 34892
rect 15752 34944 15804 34950
rect 15752 34886 15804 34892
rect 14740 34536 14792 34542
rect 14740 34478 14792 34484
rect 14752 34202 14780 34478
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14476 32978 14504 33934
rect 14556 33108 14608 33114
rect 14556 33050 14608 33056
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14200 30802 14228 31282
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14292 30938 14320 31078
rect 14384 30938 14412 31622
rect 14476 31482 14504 32914
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 14568 31414 14596 33050
rect 14648 32360 14700 32366
rect 14648 32302 14700 32308
rect 14660 31498 14688 32302
rect 14660 31470 14780 31498
rect 14556 31408 14608 31414
rect 14556 31350 14608 31356
rect 14648 31408 14700 31414
rect 14648 31350 14700 31356
rect 14556 31136 14608 31142
rect 14556 31078 14608 31084
rect 14568 30938 14596 31078
rect 14280 30932 14332 30938
rect 14280 30874 14332 30880
rect 14372 30932 14424 30938
rect 14372 30874 14424 30880
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14188 30796 14240 30802
rect 14188 30738 14240 30744
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 14094 30696 14150 30705
rect 14094 30631 14096 30640
rect 14148 30631 14150 30640
rect 14096 30602 14148 30608
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 13832 29850 13860 30126
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 14292 29510 14320 30738
rect 14660 30666 14688 31350
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 13452 29232 13504 29238
rect 13452 29174 13504 29180
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13084 24336 13136 24342
rect 13084 24278 13136 24284
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13004 23186 13032 23598
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13004 22574 13032 23122
rect 13464 22642 13492 29174
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13740 25906 13768 26862
rect 13832 26246 13860 27950
rect 13924 27674 13952 28018
rect 13912 27668 13964 27674
rect 13912 27610 13964 27616
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14660 26790 14688 27406
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13832 25838 13860 26182
rect 13924 26042 13952 26318
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13832 24818 13860 25774
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 13924 25498 13952 25638
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 14108 25294 14136 26182
rect 14568 26042 14596 26182
rect 14556 26036 14608 26042
rect 14556 25978 14608 25984
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14384 25498 14412 25774
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14752 25294 14780 31470
rect 14844 31346 14872 34886
rect 15660 34740 15712 34746
rect 15660 34682 15712 34688
rect 15672 34202 15700 34682
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14936 33658 14964 33934
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15672 32978 15700 34138
rect 15764 33658 15792 34886
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 15752 33652 15804 33658
rect 15752 33594 15804 33600
rect 15856 33522 15884 33934
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 15948 33402 15976 35702
rect 16224 35290 16252 39918
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 16592 38654 16620 39238
rect 16408 38626 16620 38654
rect 16408 36582 16436 38626
rect 16948 38344 17000 38350
rect 17328 38298 17356 41414
rect 17604 41138 17632 41550
rect 17592 41132 17644 41138
rect 17592 41074 17644 41080
rect 17604 40730 17632 41074
rect 17592 40724 17644 40730
rect 17592 40666 17644 40672
rect 17408 40520 17460 40526
rect 17408 40462 17460 40468
rect 17684 40520 17736 40526
rect 17684 40462 17736 40468
rect 17420 40118 17448 40462
rect 17408 40112 17460 40118
rect 17408 40054 17460 40060
rect 17696 39506 17724 40462
rect 17684 39500 17736 39506
rect 17684 39442 17736 39448
rect 17500 38888 17552 38894
rect 17500 38830 17552 38836
rect 16948 38286 17000 38292
rect 16488 38276 16540 38282
rect 16488 38218 16540 38224
rect 16500 37398 16528 38218
rect 16672 37732 16724 37738
rect 16672 37674 16724 37680
rect 16488 37392 16540 37398
rect 16488 37334 16540 37340
rect 16396 36576 16448 36582
rect 16396 36518 16448 36524
rect 16212 35284 16264 35290
rect 16212 35226 16264 35232
rect 16212 34944 16264 34950
rect 16212 34886 16264 34892
rect 16224 34746 16252 34886
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 15856 33374 15976 33402
rect 16028 33380 16080 33386
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15672 32434 15700 32914
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15856 32230 15884 33374
rect 16028 33322 16080 33328
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15948 32842 15976 33254
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15752 31952 15804 31958
rect 15752 31894 15804 31900
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15108 31680 15160 31686
rect 15108 31622 15160 31628
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 14844 30802 14872 31282
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14936 28762 14964 31282
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 15028 30938 15056 31078
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 15120 29306 15148 31622
rect 15212 30326 15240 31826
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15304 31346 15332 31758
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15488 31210 15516 31758
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15580 31414 15608 31690
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 15764 31346 15792 31894
rect 15856 31346 15884 32166
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15384 31136 15436 31142
rect 15384 31078 15436 31084
rect 15396 30802 15424 31078
rect 15384 30796 15436 30802
rect 15384 30738 15436 30744
rect 15200 30320 15252 30326
rect 15200 30262 15252 30268
rect 15396 29714 15424 30738
rect 15672 30734 15700 31214
rect 15764 30870 15792 31282
rect 16040 31278 16068 33322
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16316 32026 16344 32370
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 16408 31958 16436 36518
rect 16500 36174 16528 37334
rect 16684 36922 16712 37674
rect 16960 37262 16988 38286
rect 17236 38270 17356 38298
rect 17236 37890 17264 38270
rect 17316 38208 17368 38214
rect 17368 38156 17448 38162
rect 17316 38150 17448 38156
rect 17328 38134 17448 38150
rect 17236 37874 17356 37890
rect 17420 37874 17448 38134
rect 17040 37868 17092 37874
rect 17040 37810 17092 37816
rect 17236 37868 17368 37874
rect 17236 37862 17316 37868
rect 17052 37466 17080 37810
rect 17040 37460 17092 37466
rect 17040 37402 17092 37408
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 16948 37256 17000 37262
rect 16948 37198 17000 37204
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16500 34678 16528 36110
rect 16684 35680 16712 36722
rect 16764 36032 16816 36038
rect 16764 35974 16816 35980
rect 16776 35834 16804 35974
rect 16868 35834 16896 37198
rect 16960 36242 16988 37198
rect 17052 36786 17080 37402
rect 17236 36854 17264 37862
rect 17316 37810 17368 37816
rect 17408 37868 17460 37874
rect 17408 37810 17460 37816
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 17328 36922 17356 37130
rect 17316 36916 17368 36922
rect 17316 36858 17368 36864
rect 17132 36848 17184 36854
rect 17132 36790 17184 36796
rect 17224 36848 17276 36854
rect 17224 36790 17276 36796
rect 17040 36780 17092 36786
rect 17040 36722 17092 36728
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 16764 35828 16816 35834
rect 16764 35770 16816 35776
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 16764 35692 16816 35698
rect 16684 35652 16764 35680
rect 16764 35634 16816 35640
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16580 34672 16632 34678
rect 16580 34614 16632 34620
rect 16592 32570 16620 34614
rect 16580 32564 16632 32570
rect 16580 32506 16632 32512
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16592 31754 16620 32506
rect 16592 31726 16712 31754
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 14924 28756 14976 28762
rect 14924 28698 14976 28704
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14936 27334 14964 28562
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 14936 27130 14964 27270
rect 14924 27124 14976 27130
rect 14924 27066 14976 27072
rect 15120 26518 15148 27474
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 15580 24954 15608 30126
rect 16040 29730 16068 31214
rect 16500 30666 16528 31282
rect 16488 30660 16540 30666
rect 16488 30602 16540 30608
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 15948 29702 16068 29730
rect 16592 29714 16620 30126
rect 16580 29708 16632 29714
rect 15660 28144 15712 28150
rect 15660 28086 15712 28092
rect 15672 27674 15700 28086
rect 15844 27872 15896 27878
rect 15844 27814 15896 27820
rect 15660 27668 15712 27674
rect 15660 27610 15712 27616
rect 15672 26858 15700 27610
rect 15856 27470 15884 27814
rect 15948 27470 15976 29702
rect 16580 29650 16632 29656
rect 16028 29572 16080 29578
rect 16028 29514 16080 29520
rect 16040 29306 16068 29514
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 16396 28552 16448 28558
rect 16396 28494 16448 28500
rect 16408 28218 16436 28494
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 15660 26852 15712 26858
rect 15660 26794 15712 26800
rect 15672 25974 15700 26794
rect 16408 26450 16436 27406
rect 16592 27334 16620 29650
rect 16684 28558 16712 31726
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16684 28014 16712 28494
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16684 27470 16712 27950
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16592 26926 16620 27270
rect 16776 27130 16804 35634
rect 16868 35154 16896 35770
rect 16960 35154 16988 36178
rect 16856 35148 16908 35154
rect 16856 35090 16908 35096
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 16868 34746 16896 35090
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17144 34610 17172 36790
rect 17512 36242 17540 38830
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 17788 38010 17816 38150
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17316 35012 17368 35018
rect 17316 34954 17368 34960
rect 17328 34746 17356 34954
rect 17316 34740 17368 34746
rect 17316 34682 17368 34688
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17144 34490 17172 34546
rect 16960 34462 17172 34490
rect 16960 29306 16988 34462
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 17144 30802 17172 33390
rect 17236 33318 17264 34546
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 17316 33448 17368 33454
rect 17316 33390 17368 33396
rect 17224 33312 17276 33318
rect 17224 33254 17276 33260
rect 17236 33114 17264 33254
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17222 32872 17278 32881
rect 17222 32807 17224 32816
rect 17276 32807 17278 32816
rect 17224 32778 17276 32784
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17236 29714 17264 32778
rect 17328 31890 17356 33390
rect 17604 33114 17632 33866
rect 17592 33108 17644 33114
rect 17592 33050 17644 33056
rect 17604 32230 17632 33050
rect 17880 32910 17908 44338
rect 17960 44328 18012 44334
rect 17960 44270 18012 44276
rect 17972 43314 18000 44270
rect 18420 43648 18472 43654
rect 18420 43590 18472 43596
rect 17960 43308 18012 43314
rect 17960 43250 18012 43256
rect 17972 42022 18000 43250
rect 18432 43246 18460 43590
rect 18144 43240 18196 43246
rect 18144 43182 18196 43188
rect 18420 43240 18472 43246
rect 18420 43182 18472 43188
rect 18156 42906 18184 43182
rect 18144 42900 18196 42906
rect 18144 42842 18196 42848
rect 18328 42628 18380 42634
rect 18328 42570 18380 42576
rect 18340 42362 18368 42570
rect 18524 42378 18552 44338
rect 18604 44192 18656 44198
rect 18604 44134 18656 44140
rect 18616 43858 18644 44134
rect 18604 43852 18656 43858
rect 18604 43794 18656 43800
rect 19064 43784 19116 43790
rect 19064 43726 19116 43732
rect 19076 43246 19104 43726
rect 19064 43240 19116 43246
rect 19064 43182 19116 43188
rect 19168 43092 19196 44338
rect 19432 44328 19484 44334
rect 19432 44270 19484 44276
rect 19444 44146 19472 44270
rect 19260 44118 19472 44146
rect 19260 43790 19288 44118
rect 20088 43858 20116 44406
rect 20640 44198 20668 44406
rect 20628 44192 20680 44198
rect 20628 44134 20680 44140
rect 20536 43988 20588 43994
rect 20536 43930 20588 43936
rect 20076 43852 20128 43858
rect 20076 43794 20128 43800
rect 19248 43784 19300 43790
rect 19248 43726 19300 43732
rect 19076 43064 19196 43092
rect 18604 42764 18656 42770
rect 18604 42706 18656 42712
rect 18432 42362 18552 42378
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 18420 42356 18552 42362
rect 18472 42350 18552 42356
rect 18420 42298 18472 42304
rect 18144 42084 18196 42090
rect 18144 42026 18196 42032
rect 17960 42016 18012 42022
rect 17960 41958 18012 41964
rect 17972 41478 18000 41958
rect 18156 41546 18184 42026
rect 18432 41818 18460 42298
rect 18420 41812 18472 41818
rect 18420 41754 18472 41760
rect 18144 41540 18196 41546
rect 18144 41482 18196 41488
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 18156 41138 18184 41482
rect 18616 41414 18644 42706
rect 18788 42220 18840 42226
rect 18788 42162 18840 42168
rect 18800 41682 18828 42162
rect 18972 42016 19024 42022
rect 18972 41958 19024 41964
rect 18984 41818 19012 41958
rect 18972 41812 19024 41818
rect 18972 41754 19024 41760
rect 19076 41698 19104 43064
rect 19260 42770 19288 43726
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 20088 43246 20116 43794
rect 20548 43246 20576 43930
rect 20640 43790 20668 44134
rect 20628 43784 20680 43790
rect 20628 43726 20680 43732
rect 20812 43784 20864 43790
rect 20812 43726 20864 43732
rect 20640 43314 20668 43726
rect 20824 43382 20852 43726
rect 20996 43648 21048 43654
rect 20996 43590 21048 43596
rect 21008 43450 21036 43590
rect 20996 43444 21048 43450
rect 20996 43386 21048 43392
rect 20812 43376 20864 43382
rect 20812 43318 20864 43324
rect 20628 43308 20680 43314
rect 20628 43250 20680 43256
rect 20076 43240 20128 43246
rect 20536 43240 20588 43246
rect 20076 43182 20128 43188
rect 20272 43200 20536 43228
rect 19248 42764 19300 42770
rect 19248 42706 19300 42712
rect 19156 42560 19208 42566
rect 19156 42502 19208 42508
rect 19168 42362 19196 42502
rect 19260 42362 19288 42706
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19156 42356 19208 42362
rect 19156 42298 19208 42304
rect 19248 42356 19300 42362
rect 19248 42298 19300 42304
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 19352 41818 19380 42094
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 18788 41676 18840 41682
rect 18788 41618 18840 41624
rect 18984 41670 19104 41698
rect 18524 41386 18644 41414
rect 18144 41132 18196 41138
rect 18144 41074 18196 41080
rect 17960 41064 18012 41070
rect 17960 41006 18012 41012
rect 17972 40730 18000 41006
rect 17960 40724 18012 40730
rect 17960 40666 18012 40672
rect 17960 40520 18012 40526
rect 17960 40462 18012 40468
rect 17972 39642 18000 40462
rect 17960 39636 18012 39642
rect 17960 39578 18012 39584
rect 18156 39302 18184 41074
rect 18524 40050 18552 41386
rect 18788 40520 18840 40526
rect 18788 40462 18840 40468
rect 18512 40044 18564 40050
rect 18512 39986 18564 39992
rect 18420 39908 18472 39914
rect 18420 39850 18472 39856
rect 18432 39506 18460 39850
rect 18524 39506 18552 39986
rect 18800 39982 18828 40462
rect 18788 39976 18840 39982
rect 18788 39918 18840 39924
rect 18420 39500 18472 39506
rect 18420 39442 18472 39448
rect 18512 39500 18564 39506
rect 18512 39442 18564 39448
rect 18880 39432 18932 39438
rect 18880 39374 18932 39380
rect 18144 39296 18196 39302
rect 18144 39238 18196 39244
rect 18156 38826 18184 39238
rect 18892 39098 18920 39374
rect 18880 39092 18932 39098
rect 18880 39034 18932 39040
rect 18144 38820 18196 38826
rect 18144 38762 18196 38768
rect 17960 38276 18012 38282
rect 17960 38218 18012 38224
rect 17972 38010 18000 38218
rect 17960 38004 18012 38010
rect 17960 37946 18012 37952
rect 18052 35488 18104 35494
rect 18052 35430 18104 35436
rect 18064 34542 18092 35430
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 17868 32904 17920 32910
rect 17972 32881 18000 34138
rect 17868 32846 17920 32852
rect 17958 32872 18014 32881
rect 17958 32807 18014 32816
rect 17972 32502 18000 32807
rect 17960 32496 18012 32502
rect 17960 32438 18012 32444
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 18052 32224 18104 32230
rect 18052 32166 18104 32172
rect 17316 31884 17368 31890
rect 17316 31826 17368 31832
rect 17328 30938 17356 31826
rect 17316 30932 17368 30938
rect 17316 30874 17368 30880
rect 17328 30376 17356 30874
rect 17328 30348 17448 30376
rect 17316 30048 17368 30054
rect 17316 29990 17368 29996
rect 17224 29708 17276 29714
rect 17052 29668 17224 29696
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 17052 29186 17080 29668
rect 17224 29650 17276 29656
rect 17328 29578 17356 29990
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 16868 29158 17080 29186
rect 17132 29164 17184 29170
rect 16868 28098 16896 29158
rect 17132 29106 17184 29112
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 16960 28762 16988 28970
rect 16948 28756 17000 28762
rect 16948 28698 17000 28704
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 28218 16988 28358
rect 17144 28218 17172 29106
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 16868 28070 16988 28098
rect 16960 27606 16988 28070
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17052 27674 17080 28018
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 15856 26042 15884 26386
rect 16592 26314 16620 26862
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15568 24948 15620 24954
rect 15568 24890 15620 24896
rect 15672 24886 15700 25910
rect 16592 25906 16620 26250
rect 16776 25974 16804 27066
rect 16960 26314 16988 27542
rect 17144 27130 17172 27814
rect 17236 27674 17264 27814
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 17420 26518 17448 30348
rect 18064 30258 18092 32166
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18052 30116 18104 30122
rect 18052 30058 18104 30064
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17972 29646 18000 29990
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17512 29306 17540 29446
rect 17880 29306 17908 29446
rect 18064 29306 18092 30058
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17512 28082 17540 28902
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17972 28218 18000 28358
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 18064 27538 18092 28562
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 18064 26994 18092 27338
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17960 26852 18012 26858
rect 17960 26794 18012 26800
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 16592 24818 16620 25842
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13832 24562 13860 24618
rect 13832 24534 13952 24562
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 21554 12940 22374
rect 13464 22234 13492 22578
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13556 22098 13584 23598
rect 13832 23322 13860 23598
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13556 21622 13584 22034
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13096 21146 13124 21490
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13924 20942 13952 24534
rect 14108 24410 14136 24686
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15764 24410 15792 24550
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 14556 24200 14608 24206
rect 14740 24200 14792 24206
rect 14556 24142 14608 24148
rect 14660 24148 14740 24154
rect 14660 24142 14792 24148
rect 14568 23866 14596 24142
rect 14660 24126 14780 24142
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14384 21622 14412 23258
rect 14476 23050 14504 23462
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14372 21616 14424 21622
rect 14372 21558 14424 21564
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 19922 13124 20198
rect 13740 20058 13768 20402
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14292 20058 14320 20334
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14476 19938 14504 22986
rect 14660 22982 14688 24126
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15120 23322 15148 23734
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15304 23186 15332 24006
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 20602 14596 20742
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 14384 19910 14504 19938
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18426 12848 18566
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 13004 17882 13032 18702
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13464 17746 13492 19382
rect 14384 18358 14412 19910
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 14384 17678 14412 18294
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12912 16046 12940 17138
rect 13096 16794 13124 17478
rect 13464 17202 13492 17478
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 14384 17134 14412 17478
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13096 16250 13124 16730
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 12728 14618 12756 15982
rect 12912 15570 12940 15982
rect 13556 15706 13584 15982
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13648 15638 13676 15846
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13938 12572 14282
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 14006 13124 14214
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13556 13938 13584 14418
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11256 13190 11284 13330
rect 11428 13320 11480 13326
rect 12072 13320 12124 13326
rect 11428 13262 11480 13268
rect 11794 13288 11850 13297
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11348 12866 11376 13194
rect 11440 12986 11468 13262
rect 12072 13262 12124 13268
rect 11794 13223 11796 13232
rect 11848 13223 11850 13232
rect 11796 13194 11848 13200
rect 11886 13016 11942 13025
rect 11428 12980 11480 12986
rect 11886 12951 11942 12960
rect 11428 12922 11480 12928
rect 11900 12918 11928 12951
rect 11888 12912 11940 12918
rect 11348 12838 11468 12866
rect 11888 12854 11940 12860
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12322 11284 12582
rect 11256 12294 11376 12322
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11256 9602 11284 12174
rect 11348 11529 11376 12294
rect 11440 11762 11468 12838
rect 11520 12776 11572 12782
rect 11572 12736 11652 12764
rect 11520 12718 11572 12724
rect 11624 12442 11652 12736
rect 11796 12708 11848 12714
rect 11716 12668 11796 12696
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11334 11520 11390 11529
rect 11334 11455 11390 11464
rect 11348 11218 11376 11455
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11334 11112 11390 11121
rect 11334 11047 11336 11056
rect 11388 11047 11390 11056
rect 11336 11018 11388 11024
rect 11348 10062 11376 11018
rect 11440 10674 11468 11698
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11440 9926 11468 10610
rect 11532 10538 11560 11562
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11532 10062 11560 10474
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11256 9574 11376 9602
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7426 11100 7822
rect 11164 7546 11192 9454
rect 11256 9178 11284 9454
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11072 7398 11192 7426
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 6254 10732 6666
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5234 10824 5510
rect 11072 5234 11100 7210
rect 11164 6798 11192 7398
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11256 7002 11284 7346
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11164 6322 11192 6734
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6322 11284 6598
rect 11348 6322 11376 9574
rect 11518 9208 11574 9217
rect 11518 9143 11520 9152
rect 11572 9143 11574 9152
rect 11520 9114 11572 9120
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8809 11560 8910
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11532 8634 11560 8735
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 7886 11468 8230
rect 11428 7880 11480 7886
rect 11624 7834 11652 12378
rect 11716 12374 11744 12668
rect 11796 12650 11848 12656
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11898 11744 12038
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11900 11218 11928 12854
rect 11978 12744 12034 12753
rect 11978 12679 12034 12688
rect 11992 12442 12020 12679
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11980 11892 12032 11898
rect 12084 11880 12112 13262
rect 12268 13190 12296 13466
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12032 11852 12112 11880
rect 11980 11834 12032 11840
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12084 11354 12112 11630
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10810 12112 10950
rect 12176 10810 12204 11630
rect 12268 11082 12296 13126
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11716 9761 11744 10610
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11808 10198 11836 10474
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11702 9752 11758 9761
rect 11702 9687 11758 9696
rect 11900 8498 11928 10406
rect 11992 10305 12020 10474
rect 11978 10296 12034 10305
rect 11978 10231 12034 10240
rect 11992 9178 12020 10231
rect 12084 10130 12112 10474
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12162 9752 12218 9761
rect 12162 9687 12218 9696
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 8498 12020 9114
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11704 8424 11756 8430
rect 12084 8378 12112 8774
rect 12176 8634 12204 9687
rect 12268 9586 12296 11018
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11704 8366 11756 8372
rect 11428 7822 11480 7828
rect 11532 7806 11652 7834
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7546 11468 7686
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6798 11468 7142
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11164 6118 11192 6258
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10980 3738 11008 4966
rect 11072 4554 11100 5170
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11060 3392 11112 3398
rect 11164 3380 11192 6054
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11256 4826 11284 5170
rect 11440 4826 11468 6734
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11348 4554 11376 4762
rect 11532 4706 11560 7806
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7478 11652 7686
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11716 7256 11744 8366
rect 11992 8350 12112 8378
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7954 11928 8230
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11624 7228 11744 7256
rect 11796 7268 11848 7274
rect 11624 5692 11652 7228
rect 11796 7210 11848 7216
rect 11702 7168 11758 7177
rect 11808 7154 11836 7210
rect 11758 7126 11836 7154
rect 11702 7103 11758 7112
rect 11716 6798 11744 7103
rect 11704 6792 11756 6798
rect 11756 6752 11836 6780
rect 11704 6734 11756 6740
rect 11624 5664 11744 5692
rect 11440 4678 11560 4706
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4146 11376 4490
rect 11440 4185 11468 4678
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11426 4176 11482 4185
rect 11336 4140 11388 4146
rect 11426 4111 11482 4120
rect 11336 4082 11388 4088
rect 11348 3670 11376 4082
rect 11440 4078 11468 4111
rect 11624 4078 11652 4558
rect 11428 4072 11480 4078
rect 11612 4072 11664 4078
rect 11428 4014 11480 4020
rect 11532 4032 11612 4060
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11532 3534 11560 4032
rect 11612 4014 11664 4020
rect 11716 3670 11744 5664
rect 11808 4826 11836 6752
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6497 11928 6666
rect 11886 6488 11942 6497
rect 11886 6423 11942 6432
rect 11886 5536 11942 5545
rect 11886 5471 11942 5480
rect 11900 5098 11928 5471
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11900 5001 11928 5034
rect 11886 4992 11942 5001
rect 11886 4927 11942 4936
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11992 4010 12020 8350
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 5370 12112 8230
rect 12176 7342 12204 8570
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12268 8090 12296 8434
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12360 7410 12388 11834
rect 12452 7546 12480 13874
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11558 12572 12038
rect 12636 11762 12664 13874
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12912 12986 12940 13738
rect 13648 13530 13676 13942
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14108 13841 14136 13874
rect 14200 13870 14228 14826
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 13864 14240 13870
rect 14094 13832 14150 13841
rect 14188 13806 14240 13812
rect 14094 13767 14150 13776
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12728 12374 12756 12718
rect 13280 12434 13308 13262
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13188 12406 13308 12434
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12728 11762 12756 12310
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11898 13124 12174
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12530 11384 12586 11393
rect 12530 11319 12586 11328
rect 12544 11150 12572 11319
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10305 12664 10610
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12544 9081 12572 9114
rect 12530 9072 12586 9081
rect 12530 9007 12586 9016
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12544 7018 12572 8298
rect 12452 6990 12572 7018
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6390 12204 6666
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 6089 12296 6258
rect 12254 6080 12310 6089
rect 12254 6015 12310 6024
rect 12268 5574 12296 6015
rect 12452 5710 12480 6990
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12544 6730 12572 6870
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12636 6458 12664 10134
rect 12728 9178 12756 11494
rect 12820 10742 12848 11834
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12716 6656 12768 6662
rect 12820 6644 12848 10678
rect 12912 8634 12940 11698
rect 13188 11354 13216 12406
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13004 10810 13032 11018
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13096 10674 13124 11290
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13280 10130 13308 11154
rect 13556 11150 13584 12854
rect 14108 12442 14136 13262
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13266 9616 13322 9625
rect 13266 9551 13268 9560
rect 13320 9551 13322 9560
rect 13268 9522 13320 9528
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13188 9110 13216 9279
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13372 8974 13400 10610
rect 12992 8968 13044 8974
rect 13360 8968 13412 8974
rect 13044 8916 13308 8922
rect 12992 8910 13308 8916
rect 13360 8910 13412 8916
rect 13004 8906 13308 8910
rect 13004 8900 13320 8906
rect 13004 8894 13268 8900
rect 13268 8842 13320 8848
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12912 7886 12940 8570
rect 13188 8498 13216 8570
rect 13280 8498 13308 8842
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12768 6616 12848 6644
rect 12716 6598 12768 6604
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 12084 3534 12112 4082
rect 12176 3942 12204 5034
rect 12268 4214 12296 5510
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12348 4072 12400 4078
rect 12254 4040 12310 4049
rect 12348 4014 12400 4020
rect 12254 3975 12310 3984
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12268 3670 12296 3975
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11112 3352 11192 3380
rect 11060 3334 11112 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 8760 3120 8812 3126
rect 8758 3088 8760 3097
rect 9312 3120 9364 3126
rect 8812 3088 8814 3097
rect 8116 3052 8168 3058
rect 9312 3062 9364 3068
rect 10980 3058 11008 3334
rect 11532 3194 11560 3470
rect 12176 3448 12204 3606
rect 12360 3602 12388 4014
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12452 3534 12480 5646
rect 12636 5234 12664 6054
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12728 4622 12756 6598
rect 12912 5914 12940 7278
rect 13096 6662 13124 7754
rect 13188 7274 13216 8434
rect 13280 8090 13308 8434
rect 13372 8294 13400 8910
rect 13464 8294 13492 11086
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13372 7546 13400 8230
rect 13464 8090 13492 8230
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13556 7818 13584 11086
rect 13648 9489 13676 11630
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13634 9480 13690 9489
rect 13740 9466 13768 9590
rect 13832 9586 13860 12310
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14016 11608 14044 12242
rect 14094 12200 14150 12209
rect 14094 12135 14096 12144
rect 14148 12135 14150 12144
rect 14096 12106 14148 12112
rect 14096 11620 14148 11626
rect 14016 11580 14096 11608
rect 14096 11562 14148 11568
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13924 10985 13952 11018
rect 13910 10976 13966 10985
rect 13910 10911 13966 10920
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13740 9438 13860 9466
rect 13634 9415 13690 9424
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13648 8974 13676 9114
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8362 13676 8910
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13544 7812 13596 7818
rect 13464 7772 13544 7800
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5794 13032 6190
rect 12912 5766 13032 5794
rect 12912 5642 12940 5766
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12912 5370 12940 5578
rect 12992 5568 13044 5574
rect 13096 5556 13124 6598
rect 13358 6216 13414 6225
rect 13358 6151 13414 6160
rect 13372 6118 13400 6151
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5914 13400 6054
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13044 5528 13124 5556
rect 12992 5510 13044 5516
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12544 3534 12572 4558
rect 12716 4072 12768 4078
rect 12900 4072 12952 4078
rect 12716 4014 12768 4020
rect 12898 4040 12900 4049
rect 12952 4040 12954 4049
rect 12728 3738 12756 4014
rect 12898 3975 12954 3984
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12440 3528 12492 3534
rect 12254 3496 12310 3505
rect 12440 3470 12492 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12176 3440 12254 3448
rect 12176 3420 12256 3440
rect 12308 3431 12310 3440
rect 12716 3460 12768 3466
rect 12256 3402 12308 3408
rect 12716 3402 12768 3408
rect 12728 3194 12756 3402
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 13004 3126 13032 5510
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13096 4010 13124 4762
rect 13084 4004 13136 4010
rect 13084 3946 13136 3952
rect 13188 3890 13216 5578
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13280 4622 13308 5170
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13266 3904 13322 3913
rect 13188 3862 13266 3890
rect 13266 3839 13322 3848
rect 13372 3670 13400 4762
rect 13464 4690 13492 7772
rect 13544 7754 13596 7760
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13648 6390 13676 7210
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13740 6202 13768 8434
rect 13832 7002 13860 9438
rect 13924 8945 13952 10911
rect 14108 10470 14136 11562
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10742 14228 11018
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 9648 14056 9654
rect 14188 9648 14240 9654
rect 14004 9590 14056 9596
rect 14108 9608 14188 9636
rect 14016 9178 14044 9590
rect 14108 9450 14136 9608
rect 14188 9590 14240 9596
rect 14186 9480 14242 9489
rect 14096 9444 14148 9450
rect 14186 9415 14242 9424
rect 14096 9386 14148 9392
rect 14108 9178 14136 9386
rect 14200 9382 14228 9415
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14188 8968 14240 8974
rect 13910 8936 13966 8945
rect 14188 8910 14240 8916
rect 13910 8871 13966 8880
rect 13924 8498 13952 8871
rect 14004 8832 14056 8838
rect 14200 8809 14228 8910
rect 14004 8774 14056 8780
rect 14186 8800 14242 8809
rect 14016 8566 14044 8774
rect 14186 8735 14242 8744
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14016 6730 14044 8502
rect 14200 7410 14228 8735
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13648 6186 13768 6202
rect 13636 6180 13768 6186
rect 13688 6174 13768 6180
rect 13636 6122 13688 6128
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5953 13584 6054
rect 13542 5944 13598 5953
rect 13648 5914 13676 6122
rect 13728 6112 13780 6118
rect 13726 6080 13728 6089
rect 13780 6080 13782 6089
rect 13726 6015 13782 6024
rect 13542 5879 13598 5888
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13544 5704 13596 5710
rect 13542 5672 13544 5681
rect 13596 5672 13598 5681
rect 13542 5607 13598 5616
rect 13740 5302 13768 6015
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 8758 3023 8814 3032
rect 10968 3052 11020 3058
rect 8116 2994 8168 3000
rect 10968 2994 11020 3000
rect 13188 2922 13216 3402
rect 13372 3194 13400 3470
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13464 2990 13492 4014
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3534 13584 3878
rect 13740 3738 13768 5238
rect 13832 4826 13860 5646
rect 13924 5545 13952 5646
rect 13910 5536 13966 5545
rect 13910 5471 13966 5480
rect 13912 5296 13964 5302
rect 14016 5284 14044 6326
rect 14108 5710 14136 6598
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14200 5574 14228 6326
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 13964 5256 14044 5284
rect 13912 5238 13964 5244
rect 13924 5098 13952 5238
rect 14200 5234 14228 5510
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13818 3904 13874 3913
rect 13818 3839 13874 3848
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13728 3528 13780 3534
rect 13832 3516 13860 3839
rect 13780 3488 13860 3516
rect 13728 3470 13780 3476
rect 13924 3466 13952 4626
rect 14200 3534 14228 4626
rect 14292 4146 14320 14350
rect 14476 14074 14504 19790
rect 14568 19718 14596 20538
rect 14660 20534 14688 22918
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14752 20398 14780 20946
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14752 19514 14780 20334
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14660 18834 14688 19314
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14660 17678 14688 18770
rect 14936 17814 14964 22646
rect 15120 22094 15148 23122
rect 15396 23118 15424 23462
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15856 22574 15884 24550
rect 16224 23526 16252 24686
rect 16592 24274 16620 24754
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15028 22066 15148 22094
rect 15028 19922 15056 22066
rect 15660 21956 15712 21962
rect 15660 21898 15712 21904
rect 15672 21690 15700 21898
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 20942 15148 21422
rect 16040 21146 16068 21490
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 16224 20602 16252 23462
rect 16776 23118 16804 25910
rect 17420 25770 17448 26454
rect 17408 25764 17460 25770
rect 17408 25706 17460 25712
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16960 24410 16988 24686
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17144 24206 17172 25094
rect 17684 24608 17736 24614
rect 17788 24596 17816 25298
rect 17736 24568 17816 24596
rect 17684 24550 17736 24556
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17604 23866 17632 24074
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 20058 15516 20198
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19514 15240 19858
rect 15752 19780 15804 19786
rect 15856 19768 15884 19994
rect 15804 19740 15884 19768
rect 15752 19722 15804 19728
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15028 18970 15056 19246
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15764 18834 15792 19722
rect 16040 19514 16068 20334
rect 16224 19718 16252 20538
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 16040 18766 16068 19450
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14568 16794 14596 17614
rect 14936 17134 14964 17750
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14936 16590 14964 17070
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 15910 15148 16390
rect 15488 16182 15516 17138
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15120 15502 15148 15846
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 14618 14596 15302
rect 16040 14618 16068 18566
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17610 16344 18022
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16408 17270 16436 23054
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 22710 17080 22918
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 22030 16712 22510
rect 17236 22094 17264 23054
rect 17420 22710 17448 23258
rect 17512 23050 17540 23258
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17788 22982 17816 24568
rect 17972 24018 18000 26794
rect 18064 25974 18092 26930
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18064 24138 18092 25910
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 17972 23990 18092 24018
rect 18064 23050 18092 23990
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17408 22704 17460 22710
rect 17460 22652 17724 22658
rect 17408 22646 17724 22652
rect 17420 22630 17724 22646
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17604 22234 17632 22374
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17236 22066 17448 22094
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16684 21690 16712 21966
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16776 19786 16804 21966
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19514 16804 19722
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 17144 19174 17172 20742
rect 17328 20058 17356 20946
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17328 19378 17356 19790
rect 17420 19786 17448 22066
rect 17696 22030 17724 22630
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17788 21962 17816 22918
rect 17972 22438 18000 22918
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22030 18000 22374
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17880 20466 17908 21626
rect 17972 20942 18000 21830
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17880 19378 17908 20402
rect 18156 20058 18184 38762
rect 18984 38758 19012 41670
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19444 41206 19472 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19432 41200 19484 41206
rect 19432 41142 19484 41148
rect 19156 40928 19208 40934
rect 19156 40870 19208 40876
rect 20076 40928 20128 40934
rect 20076 40870 20128 40876
rect 19168 40730 19196 40870
rect 19156 40724 19208 40730
rect 19156 40666 19208 40672
rect 19064 40384 19116 40390
rect 19064 40326 19116 40332
rect 19076 40118 19104 40326
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19156 40180 19208 40186
rect 19156 40122 19208 40128
rect 19064 40112 19116 40118
rect 19064 40054 19116 40060
rect 18972 38752 19024 38758
rect 18972 38694 19024 38700
rect 18880 38344 18932 38350
rect 18880 38286 18932 38292
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18524 37330 18552 37810
rect 18892 37670 18920 38286
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18512 37324 18564 37330
rect 18432 37284 18512 37312
rect 18432 35086 18460 37284
rect 18512 37266 18564 37272
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 18800 36922 18828 37062
rect 18892 36922 18920 37606
rect 19168 37262 19196 40122
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 20088 39098 20116 40870
rect 20168 40452 20220 40458
rect 20168 40394 20220 40400
rect 20180 40118 20208 40394
rect 20168 40112 20220 40118
rect 20168 40054 20220 40060
rect 20272 39846 20300 43200
rect 20536 43182 20588 43188
rect 20352 42356 20404 42362
rect 20352 42298 20404 42304
rect 20364 40594 20392 42298
rect 20640 42226 20668 43250
rect 24032 43240 24084 43246
rect 24032 43182 24084 43188
rect 21456 43104 21508 43110
rect 21456 43046 21508 43052
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 20352 40588 20404 40594
rect 20352 40530 20404 40536
rect 20456 40118 20484 41006
rect 20640 40594 20668 42162
rect 20904 42016 20956 42022
rect 20904 41958 20956 41964
rect 20916 41818 20944 41958
rect 20904 41812 20956 41818
rect 20904 41754 20956 41760
rect 20812 41608 20864 41614
rect 20812 41550 20864 41556
rect 20824 41274 20852 41550
rect 20812 41268 20864 41274
rect 20812 41210 20864 41216
rect 20628 40588 20680 40594
rect 20628 40530 20680 40536
rect 21008 40118 21036 42570
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 21100 40186 21128 40666
rect 21088 40180 21140 40186
rect 21088 40122 21140 40128
rect 20444 40112 20496 40118
rect 20444 40054 20496 40060
rect 20996 40112 21048 40118
rect 20996 40054 21048 40060
rect 20720 39976 20772 39982
rect 20720 39918 20772 39924
rect 20260 39840 20312 39846
rect 20260 39782 20312 39788
rect 20076 39092 20128 39098
rect 20076 39034 20128 39040
rect 20272 38894 20300 39782
rect 20732 39642 20760 39918
rect 20720 39636 20772 39642
rect 20720 39578 20772 39584
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20812 39432 20864 39438
rect 20812 39374 20864 39380
rect 20352 39296 20404 39302
rect 20352 39238 20404 39244
rect 20364 38962 20392 39238
rect 20352 38956 20404 38962
rect 20352 38898 20404 38904
rect 20260 38888 20312 38894
rect 20260 38830 20312 38836
rect 20640 38758 20668 39374
rect 20824 39098 20852 39374
rect 21272 39296 21324 39302
rect 21272 39238 21324 39244
rect 20812 39092 20864 39098
rect 20812 39034 20864 39040
rect 20628 38752 20680 38758
rect 20628 38694 20680 38700
rect 20260 38276 20312 38282
rect 20260 38218 20312 38224
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 20272 38010 20300 38218
rect 20640 38214 20668 38694
rect 20720 38412 20772 38418
rect 20720 38354 20772 38360
rect 20628 38208 20680 38214
rect 20628 38150 20680 38156
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 19156 37256 19208 37262
rect 19156 37198 19208 37204
rect 19064 37188 19116 37194
rect 19064 37130 19116 37136
rect 18972 37120 19024 37126
rect 18972 37062 19024 37068
rect 18788 36916 18840 36922
rect 18788 36858 18840 36864
rect 18880 36916 18932 36922
rect 18880 36858 18932 36864
rect 18984 36786 19012 37062
rect 19076 36786 19104 37130
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 18972 36780 19024 36786
rect 18972 36722 19024 36728
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18616 35290 18644 35566
rect 18604 35284 18656 35290
rect 18604 35226 18656 35232
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 18800 34746 18828 36722
rect 18972 35488 19024 35494
rect 18972 35430 19024 35436
rect 18880 35080 18932 35086
rect 18880 35022 18932 35028
rect 18892 34746 18920 35022
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 18880 34740 18932 34746
rect 18880 34682 18932 34688
rect 18984 34626 19012 35430
rect 18800 34598 19012 34626
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18432 32842 18460 33458
rect 18512 33448 18564 33454
rect 18512 33390 18564 33396
rect 18524 33114 18552 33390
rect 18512 33108 18564 33114
rect 18512 33050 18564 33056
rect 18420 32836 18472 32842
rect 18420 32778 18472 32784
rect 18696 32292 18748 32298
rect 18696 32234 18748 32240
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18524 31822 18552 32166
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18432 30734 18460 31078
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18340 30258 18368 30670
rect 18432 30326 18460 30670
rect 18420 30320 18472 30326
rect 18420 30262 18472 30268
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 18248 29186 18276 29650
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18340 29306 18368 29446
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 18248 29158 18368 29186
rect 18340 28014 18368 29158
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18340 26926 18368 27950
rect 18328 26920 18380 26926
rect 18328 26862 18380 26868
rect 18432 26858 18460 30262
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18616 29850 18644 29990
rect 18604 29844 18656 29850
rect 18604 29786 18656 29792
rect 18708 29170 18736 32234
rect 18800 30734 18828 34598
rect 19064 34468 19116 34474
rect 19064 34410 19116 34416
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 18800 30394 18828 30670
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18696 29164 18748 29170
rect 18696 29106 18748 29112
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18524 27130 18552 28494
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18420 26852 18472 26858
rect 18420 26794 18472 26800
rect 18892 25498 18920 32846
rect 18972 30728 19024 30734
rect 18972 30670 19024 30676
rect 18984 30258 19012 30670
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18432 24954 18460 25230
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18984 24818 19012 30194
rect 19076 29714 19104 34410
rect 19168 33930 19196 37198
rect 19260 36786 19288 37946
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19340 36712 19392 36718
rect 19340 36654 19392 36660
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 19352 35850 19380 36654
rect 20548 36038 20576 36654
rect 20640 36106 20668 38150
rect 20732 37874 20760 38354
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20732 37466 20760 37810
rect 20996 37800 21048 37806
rect 20996 37742 21048 37748
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20732 36242 20760 37402
rect 21008 36922 21036 37742
rect 20996 36916 21048 36922
rect 20996 36858 21048 36864
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 21192 36378 21220 36518
rect 21180 36372 21232 36378
rect 21180 36314 21232 36320
rect 20720 36236 20772 36242
rect 20720 36178 20772 36184
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 20536 36032 20588 36038
rect 20536 35974 20588 35980
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19260 35822 19380 35850
rect 20548 35834 20576 35974
rect 20536 35828 20588 35834
rect 19260 35630 19288 35822
rect 20536 35770 20588 35776
rect 20260 35760 20312 35766
rect 20260 35702 20312 35708
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19260 34746 19288 35430
rect 20272 35154 20300 35702
rect 20640 35494 20668 36042
rect 20444 35488 20496 35494
rect 20444 35430 20496 35436
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20260 35148 20312 35154
rect 20260 35090 20312 35096
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 19352 34626 19380 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19260 34610 19380 34626
rect 19248 34604 19380 34610
rect 19300 34598 19380 34604
rect 19248 34546 19300 34552
rect 19156 33924 19208 33930
rect 19156 33866 19208 33872
rect 19260 31346 19288 34546
rect 19340 34128 19392 34134
rect 19340 34070 19392 34076
rect 19352 33522 19380 34070
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 20168 33516 20220 33522
rect 20168 33458 20220 33464
rect 19444 33114 19472 33458
rect 19524 33312 19576 33318
rect 19524 33254 19576 33260
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 19536 32858 19564 33254
rect 20180 33114 20208 33458
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 19444 32830 19564 32858
rect 19996 32966 20116 32994
rect 19444 31958 19472 32830
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 31952 19484 31958
rect 19432 31894 19484 31900
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19352 31482 19380 31690
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19444 31362 19472 31894
rect 19996 31754 20024 32966
rect 20088 32910 20116 32966
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 20272 32774 20300 33594
rect 20364 32978 20392 33798
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20272 31754 20300 31962
rect 20456 31822 20484 35430
rect 20640 35086 20668 35430
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20812 34128 20864 34134
rect 20812 34070 20864 34076
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 20628 33448 20680 33454
rect 20732 33402 20760 33594
rect 20680 33396 20760 33402
rect 20628 33390 20760 33396
rect 20640 33374 20760 33390
rect 20628 33312 20680 33318
rect 20824 33300 20852 34070
rect 20904 34060 20956 34066
rect 20904 34002 20956 34008
rect 20916 33454 20944 34002
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 20680 33272 20852 33300
rect 20628 33254 20680 33260
rect 20824 32910 20852 33272
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20824 32230 20852 32846
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20812 31952 20864 31958
rect 20812 31894 20864 31900
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20444 31816 20496 31822
rect 20496 31776 20668 31804
rect 20444 31758 20496 31764
rect 19996 31726 20116 31754
rect 20088 31686 20116 31726
rect 20168 31748 20220 31754
rect 20272 31726 20392 31754
rect 20168 31690 20220 31696
rect 19984 31680 20036 31686
rect 20076 31680 20128 31686
rect 19984 31622 20036 31628
rect 20074 31648 20076 31657
rect 20128 31648 20130 31657
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19248 31340 19300 31346
rect 19444 31334 19564 31362
rect 19248 31282 19300 31288
rect 19432 31204 19484 31210
rect 19432 31146 19484 31152
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19260 30705 19288 30874
rect 19246 30696 19302 30705
rect 19246 30631 19302 30640
rect 19352 30297 19380 31078
rect 19444 30394 19472 31146
rect 19536 30938 19564 31334
rect 19524 30932 19576 30938
rect 19524 30874 19576 30880
rect 19628 30870 19656 31418
rect 19800 31204 19852 31210
rect 19800 31146 19852 31152
rect 19708 30932 19760 30938
rect 19708 30874 19760 30880
rect 19616 30864 19668 30870
rect 19616 30806 19668 30812
rect 19720 30734 19748 30874
rect 19812 30841 19840 31146
rect 19890 30968 19946 30977
rect 19890 30903 19946 30912
rect 19904 30870 19932 30903
rect 19892 30864 19944 30870
rect 19798 30832 19854 30841
rect 19892 30806 19944 30812
rect 19798 30767 19854 30776
rect 19708 30728 19760 30734
rect 19996 30716 20024 31622
rect 20074 31583 20130 31592
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 20088 30870 20116 31146
rect 20076 30864 20128 30870
rect 20180 30841 20208 31690
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20076 30806 20128 30812
rect 20166 30832 20222 30841
rect 20166 30767 20222 30776
rect 20272 30734 20300 31622
rect 19708 30670 19760 30676
rect 19812 30688 20024 30716
rect 20076 30728 20128 30734
rect 19812 30580 19840 30688
rect 20260 30728 20312 30734
rect 20128 30688 20208 30716
rect 20076 30670 20128 30676
rect 19812 30552 20024 30580
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19338 30288 19394 30297
rect 19338 30223 19340 30232
rect 19392 30223 19394 30232
rect 19800 30252 19852 30258
rect 19340 30194 19392 30200
rect 19800 30194 19852 30200
rect 19432 30184 19484 30190
rect 19812 30161 19840 30194
rect 19432 30126 19484 30132
rect 19798 30152 19854 30161
rect 19444 30054 19472 30126
rect 19996 30122 20024 30552
rect 20180 30410 20208 30688
rect 20260 30670 20312 30676
rect 20260 30592 20312 30598
rect 20258 30560 20260 30569
rect 20312 30560 20314 30569
rect 20258 30495 20314 30504
rect 20088 30382 20208 30410
rect 19798 30087 19854 30096
rect 19984 30116 20036 30122
rect 19984 30058 20036 30064
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19352 28490 19380 29106
rect 19996 28762 20024 29106
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 20088 28626 20116 30382
rect 20168 30320 20220 30326
rect 20168 30262 20220 30268
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28014 20024 28358
rect 20088 28218 20116 28562
rect 20180 28558 20208 30262
rect 20364 30258 20392 31726
rect 20444 31680 20496 31686
rect 20444 31622 20496 31628
rect 20536 31680 20588 31686
rect 20536 31622 20588 31628
rect 20456 30394 20484 31622
rect 20548 30938 20576 31622
rect 20640 31414 20668 31776
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 20732 30954 20760 31826
rect 20824 31414 20852 31894
rect 20812 31408 20864 31414
rect 20812 31350 20864 31356
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20536 30932 20588 30938
rect 20536 30874 20588 30880
rect 20640 30926 20760 30954
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20260 29708 20312 29714
rect 20260 29650 20312 29656
rect 20272 29238 20300 29650
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20364 28694 20392 29446
rect 20548 29306 20576 30670
rect 20640 30190 20668 30926
rect 20824 30734 20852 31214
rect 20916 31142 20944 33390
rect 21008 33046 21036 33390
rect 20996 33040 21048 33046
rect 20996 32982 21048 32988
rect 20996 31680 21048 31686
rect 20994 31648 20996 31657
rect 21048 31648 21050 31657
rect 20994 31583 21050 31592
rect 21100 31346 21128 33594
rect 21284 33522 21312 39238
rect 21468 33998 21496 43046
rect 24044 42906 24072 43182
rect 24320 43178 24348 45222
rect 32324 45082 32352 45222
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 41340 45082 41368 45222
rect 32312 45076 32364 45082
rect 32312 45018 32364 45024
rect 41328 45076 41380 45082
rect 41328 45018 41380 45024
rect 37004 44804 37056 44810
rect 37004 44746 37056 44752
rect 32036 44736 32088 44742
rect 32036 44678 32088 44684
rect 36912 44736 36964 44742
rect 36912 44678 36964 44684
rect 32048 44538 32076 44678
rect 36924 44538 36952 44678
rect 32036 44532 32088 44538
rect 32036 44474 32088 44480
rect 36912 44532 36964 44538
rect 36912 44474 36964 44480
rect 27344 44328 27396 44334
rect 27344 44270 27396 44276
rect 25412 44192 25464 44198
rect 25412 44134 25464 44140
rect 25424 43858 25452 44134
rect 25412 43852 25464 43858
rect 25412 43794 25464 43800
rect 27160 43240 27212 43246
rect 27160 43182 27212 43188
rect 24308 43172 24360 43178
rect 24308 43114 24360 43120
rect 24860 43104 24912 43110
rect 24860 43046 24912 43052
rect 24032 42900 24084 42906
rect 24032 42842 24084 42848
rect 24872 42702 24900 43046
rect 24860 42696 24912 42702
rect 24860 42638 24912 42644
rect 25136 42560 25188 42566
rect 25136 42502 25188 42508
rect 25148 42362 25176 42502
rect 27172 42362 27200 43182
rect 25136 42356 25188 42362
rect 25136 42298 25188 42304
rect 27160 42356 27212 42362
rect 27160 42298 27212 42304
rect 22376 42288 22428 42294
rect 22376 42230 22428 42236
rect 22100 42152 22152 42158
rect 22100 42094 22152 42100
rect 22112 41818 22140 42094
rect 22100 41812 22152 41818
rect 22100 41754 22152 41760
rect 22284 41472 22336 41478
rect 22284 41414 22336 41420
rect 22192 41200 22244 41206
rect 22192 41142 22244 41148
rect 22008 41132 22060 41138
rect 22008 41074 22060 41080
rect 22020 39982 22048 41074
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 22112 40066 22140 40326
rect 22204 40186 22232 41142
rect 22192 40180 22244 40186
rect 22192 40122 22244 40128
rect 22296 40066 22324 41414
rect 22388 40526 22416 42230
rect 27356 42226 27384 44270
rect 31668 44192 31720 44198
rect 31668 44134 31720 44140
rect 36360 44192 36412 44198
rect 36360 44134 36412 44140
rect 31680 43858 31708 44134
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 36372 43858 36400 44134
rect 31668 43852 31720 43858
rect 31668 43794 31720 43800
rect 36360 43852 36412 43858
rect 36360 43794 36412 43800
rect 31208 43784 31260 43790
rect 31208 43726 31260 43732
rect 36084 43784 36136 43790
rect 36084 43726 36136 43732
rect 29184 43648 29236 43654
rect 29184 43590 29236 43596
rect 29196 43382 29224 43590
rect 31220 43450 31248 43726
rect 32588 43716 32640 43722
rect 32588 43658 32640 43664
rect 31208 43444 31260 43450
rect 31208 43386 31260 43392
rect 29184 43376 29236 43382
rect 29184 43318 29236 43324
rect 27436 42288 27488 42294
rect 27436 42230 27488 42236
rect 27344 42220 27396 42226
rect 27344 42162 27396 42168
rect 24400 42152 24452 42158
rect 24400 42094 24452 42100
rect 26884 42152 26936 42158
rect 26884 42094 26936 42100
rect 23572 42016 23624 42022
rect 23572 41958 23624 41964
rect 23584 41818 23612 41958
rect 23572 41812 23624 41818
rect 23572 41754 23624 41760
rect 24216 41608 24268 41614
rect 24216 41550 24268 41556
rect 23572 41540 23624 41546
rect 23572 41482 23624 41488
rect 22560 41064 22612 41070
rect 22560 41006 22612 41012
rect 22928 41064 22980 41070
rect 22928 41006 22980 41012
rect 22376 40520 22428 40526
rect 22376 40462 22428 40468
rect 22112 40050 22232 40066
rect 22112 40044 22244 40050
rect 22112 40038 22192 40044
rect 22296 40038 22508 40066
rect 22192 39986 22244 39992
rect 22008 39976 22060 39982
rect 22008 39918 22060 39924
rect 22100 39296 22152 39302
rect 22100 39238 22152 39244
rect 21640 38888 21692 38894
rect 21640 38830 21692 38836
rect 21652 38214 21680 38830
rect 22112 38418 22140 39238
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 21640 38208 21692 38214
rect 21640 38150 21692 38156
rect 21548 34196 21600 34202
rect 21548 34138 21600 34144
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 21468 33522 21496 33934
rect 21560 33522 21588 34138
rect 21272 33516 21324 33522
rect 21456 33516 21508 33522
rect 21324 33476 21404 33504
rect 21272 33458 21324 33464
rect 21180 33312 21232 33318
rect 21180 33254 21232 33260
rect 21192 32774 21220 33254
rect 21272 33040 21324 33046
rect 21272 32982 21324 32988
rect 21180 32768 21232 32774
rect 21180 32710 21232 32716
rect 21192 32314 21220 32710
rect 21284 32450 21312 32982
rect 21376 32842 21404 33476
rect 21456 33458 21508 33464
rect 21548 33516 21600 33522
rect 21548 33458 21600 33464
rect 21652 32910 21680 38150
rect 22204 37754 22232 39986
rect 22376 39840 22428 39846
rect 22376 39782 22428 39788
rect 22284 39296 22336 39302
rect 22284 39238 22336 39244
rect 22296 38894 22324 39238
rect 22284 38888 22336 38894
rect 22284 38830 22336 38836
rect 22296 37942 22324 38830
rect 22284 37936 22336 37942
rect 22284 37878 22336 37884
rect 22388 37806 22416 39782
rect 22376 37800 22428 37806
rect 22204 37726 22324 37754
rect 22376 37742 22428 37748
rect 21732 37256 21784 37262
rect 21732 37198 21784 37204
rect 21744 36378 21772 37198
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22204 36378 22232 36518
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 22100 36304 22152 36310
rect 22100 36246 22152 36252
rect 22112 35630 22140 36246
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 22020 33658 22048 34478
rect 22296 34134 22324 37726
rect 22480 37466 22508 40038
rect 22572 39438 22600 41006
rect 22940 40730 22968 41006
rect 22928 40724 22980 40730
rect 22928 40666 22980 40672
rect 23584 40050 23612 41482
rect 23940 40928 23992 40934
rect 23940 40870 23992 40876
rect 23952 40730 23980 40870
rect 23940 40724 23992 40730
rect 23940 40666 23992 40672
rect 24124 40520 24176 40526
rect 24124 40462 24176 40468
rect 24136 40186 24164 40462
rect 24032 40180 24084 40186
rect 24032 40122 24084 40128
rect 24124 40180 24176 40186
rect 24124 40122 24176 40128
rect 23572 40044 23624 40050
rect 23572 39986 23624 39992
rect 22560 39432 22612 39438
rect 22560 39374 22612 39380
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22652 38752 22704 38758
rect 22652 38694 22704 38700
rect 22560 38276 22612 38282
rect 22560 38218 22612 38224
rect 22572 37670 22600 38218
rect 22664 38010 22692 38694
rect 22652 38004 22704 38010
rect 22652 37946 22704 37952
rect 22560 37664 22612 37670
rect 22560 37606 22612 37612
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 22572 37074 22600 37606
rect 22480 37046 22600 37074
rect 22480 36106 22508 37046
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 22468 36100 22520 36106
rect 22468 36042 22520 36048
rect 22572 35834 22600 36722
rect 22744 36712 22796 36718
rect 22744 36654 22796 36660
rect 22560 35828 22612 35834
rect 22560 35770 22612 35776
rect 22756 35018 22784 36654
rect 22744 35012 22796 35018
rect 22744 34954 22796 34960
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22572 34474 22600 34886
rect 22560 34468 22612 34474
rect 22560 34410 22612 34416
rect 22284 34128 22336 34134
rect 22284 34070 22336 34076
rect 22572 34066 22600 34410
rect 22560 34060 22612 34066
rect 22560 34002 22612 34008
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 21640 32904 21692 32910
rect 21640 32846 21692 32852
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 22296 32570 22324 33050
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 21284 32422 21404 32450
rect 21192 32286 21312 32314
rect 21180 32224 21232 32230
rect 21180 32166 21232 32172
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 21086 30968 21142 30977
rect 21192 30938 21220 32166
rect 21284 31482 21312 32286
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 21086 30903 21088 30912
rect 21140 30903 21142 30912
rect 21180 30932 21232 30938
rect 21088 30874 21140 30880
rect 21180 30874 21232 30880
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20902 30696 20958 30705
rect 20902 30631 20958 30640
rect 20916 30598 20944 30631
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20824 30274 20852 30534
rect 20732 30246 20852 30274
rect 21100 30258 21128 30874
rect 21284 30734 21312 31418
rect 21376 31346 21404 32422
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 21548 31748 21600 31754
rect 21548 31690 21600 31696
rect 21560 31414 21588 31690
rect 21548 31408 21600 31414
rect 21600 31356 21680 31362
rect 21548 31350 21680 31356
rect 21364 31340 21416 31346
rect 21560 31334 21680 31350
rect 21364 31282 21416 31288
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 20904 30252 20956 30258
rect 20628 30184 20680 30190
rect 20628 30126 20680 30132
rect 20732 30002 20760 30246
rect 20904 30194 20956 30200
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 20640 29974 20760 30002
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19168 27606 19196 27950
rect 19720 27674 19748 27950
rect 20088 27674 20116 28018
rect 19708 27668 19760 27674
rect 19708 27610 19760 27616
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 19156 27600 19208 27606
rect 19156 27542 19208 27548
rect 19156 27396 19208 27402
rect 19156 27338 19208 27344
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19168 24698 19196 27338
rect 20456 27282 20484 29174
rect 20640 28082 20668 29974
rect 20824 29850 20852 30126
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 20916 29306 20944 30194
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 21008 29714 21036 30126
rect 21192 29850 21220 30670
rect 21560 30433 21588 31214
rect 21546 30424 21602 30433
rect 21546 30359 21602 30368
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 20996 29708 21048 29714
rect 20996 29650 21048 29656
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 20824 28558 20852 29106
rect 21008 28626 21036 29106
rect 21192 28762 21220 29786
rect 21652 28994 21680 31334
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22020 30394 22048 30670
rect 22008 30388 22060 30394
rect 22008 30330 22060 30336
rect 22204 29238 22232 32166
rect 22572 31754 22600 34002
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22756 33114 22784 33798
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22572 31726 22784 31754
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22468 30592 22520 30598
rect 22468 30534 22520 30540
rect 22480 30190 22508 30534
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22572 30054 22600 31214
rect 22560 30048 22612 30054
rect 22560 29990 22612 29996
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 21468 28966 21680 28994
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20824 28218 20852 28494
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20456 27254 20576 27282
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19444 26586 19472 26930
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19628 25498 19656 25774
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 20272 25294 20300 26862
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19076 24670 19196 24698
rect 19076 22094 19104 24670
rect 19260 24614 19288 25094
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19168 24342 19196 24550
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23866 19288 24006
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19248 23112 19300 23118
rect 19352 23100 19380 23598
rect 19444 23594 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19300 23072 19380 23100
rect 19248 23054 19300 23060
rect 19352 22953 19380 23072
rect 19522 23080 19578 23089
rect 19522 23015 19524 23024
rect 19576 23015 19578 23024
rect 19524 22986 19576 22992
rect 19338 22944 19394 22953
rect 19338 22879 19394 22888
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22772 19484 22778
rect 19616 22772 19668 22778
rect 19484 22732 19616 22760
rect 19432 22714 19484 22720
rect 19996 22760 20024 24210
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19616 22714 19668 22720
rect 19720 22732 20024 22760
rect 19720 22642 19748 22732
rect 19890 22672 19946 22681
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19800 22636 19852 22642
rect 19890 22607 19946 22616
rect 19800 22578 19852 22584
rect 19706 22536 19762 22545
rect 19294 22500 19346 22506
rect 19706 22471 19708 22480
rect 19294 22442 19346 22448
rect 19760 22471 19762 22480
rect 19708 22442 19760 22448
rect 19306 22386 19334 22442
rect 19524 22432 19576 22438
rect 19430 22400 19486 22409
rect 19306 22358 19430 22386
rect 19524 22374 19576 22380
rect 19430 22335 19486 22344
rect 19536 22250 19564 22374
rect 19812 22250 19840 22578
rect 19536 22222 19840 22250
rect 19076 22066 19196 22094
rect 19168 21894 19196 22066
rect 19904 22012 19932 22607
rect 19996 22166 20024 22732
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19984 22024 20036 22030
rect 19904 21984 19984 22012
rect 19984 21966 20036 21972
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 21966
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18340 20534 18368 20742
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18524 20058 18552 20878
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17328 18834 17356 19314
rect 17868 19168 17920 19174
rect 18156 19122 18184 19994
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 19446 18460 19654
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 17868 19110 17920 19116
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16592 17338 16620 18226
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 17236 17134 17264 18634
rect 17328 17814 17356 18770
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 18426 17632 18634
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17880 17746 17908 19110
rect 17972 19094 18184 19122
rect 17972 18630 18000 19094
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17236 16794 17264 17070
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16250 16620 16390
rect 17512 16250 17540 17138
rect 17604 16998 17632 17546
rect 17880 17338 17908 17682
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17604 16590 17632 16934
rect 18064 16794 18092 17070
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18340 16658 18368 17070
rect 18524 16998 18552 19722
rect 18616 18970 18644 19790
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18708 16794 18736 17070
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 18340 16250 18368 16594
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17960 16176 18012 16182
rect 16302 16144 16358 16153
rect 17960 16118 18012 16124
rect 16302 16079 16358 16088
rect 16316 16046 16344 16079
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17696 15570 17724 15982
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16500 14521 16528 14826
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14618 17172 14758
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16486 14512 16542 14521
rect 16486 14447 16488 14456
rect 16540 14447 16542 14456
rect 16488 14418 16540 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16212 14408 16264 14414
rect 16764 14408 16816 14414
rect 16592 14368 16764 14396
rect 16592 14362 16620 14368
rect 16264 14356 16620 14362
rect 16212 14350 16620 14356
rect 16764 14350 16816 14356
rect 15856 14074 15884 14350
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15948 14006 15976 14350
rect 16132 14074 16160 14350
rect 16224 14334 16620 14350
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14384 13530 14412 13806
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14476 13326 14504 13670
rect 14568 13462 14596 13806
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 12434 14596 13194
rect 14738 12880 14794 12889
rect 14738 12815 14740 12824
rect 14792 12815 14794 12824
rect 14740 12786 14792 12792
rect 14844 12442 14872 13262
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14476 12406 14596 12434
rect 14832 12436 14884 12442
rect 14476 11150 14504 12406
rect 14832 12378 14884 12384
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14660 11694 14688 12038
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14568 11354 14596 11630
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11354 14688 11494
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14752 11286 14780 12038
rect 14936 11937 14964 12650
rect 15028 12646 15056 13262
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 12306 15056 12582
rect 15120 12374 15148 13330
rect 15396 12986 15424 13874
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16960 13394 16988 13806
rect 17052 13734 17080 13806
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13530 17080 13670
rect 17144 13530 17172 13942
rect 17236 13802 17264 14010
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 13530 17264 13738
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17328 13462 17356 13806
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16672 13320 16724 13326
rect 16724 13280 16896 13308
rect 16672 13262 16724 13268
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 15396 12617 15424 12786
rect 15488 12646 15516 12786
rect 15476 12640 15528 12646
rect 15382 12608 15438 12617
rect 15476 12582 15528 12588
rect 15382 12543 15438 12552
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15396 12238 15424 12378
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 14922 11928 14978 11937
rect 14922 11863 14978 11872
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 14740 11280 14792 11286
rect 15212 11257 15240 11630
rect 15304 11354 15332 12174
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14740 11222 14792 11228
rect 15198 11248 15254 11257
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14554 11112 14610 11121
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14384 9178 14412 9522
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14384 6118 14412 8910
rect 14476 8634 14504 11086
rect 14554 11047 14610 11056
rect 14568 8974 14596 11047
rect 14752 10742 14780 11222
rect 15198 11183 15254 11192
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14844 10742 14872 11086
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 10062 14780 10542
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14648 9648 14700 9654
rect 14646 9616 14648 9625
rect 14700 9616 14702 9625
rect 14646 9551 14702 9560
rect 14752 8974 14780 9998
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14568 8634 14596 8910
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14464 6792 14516 6798
rect 14516 6740 14596 6746
rect 14464 6734 14596 6740
rect 14476 6718 14596 6734
rect 14568 6458 14596 6718
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14568 5914 14596 6394
rect 14660 6322 14688 7210
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 4214 14412 5306
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14476 3466 14504 3674
rect 14568 3534 14596 5238
rect 14660 5166 14688 6258
rect 14752 6066 14780 8910
rect 14844 6882 14872 10678
rect 15304 9353 15332 11290
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15396 10810 15424 11154
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 9994 15516 12582
rect 15856 12442 15884 12786
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15568 12232 15620 12238
rect 15752 12232 15804 12238
rect 15568 12174 15620 12180
rect 15658 12200 15714 12209
rect 15580 11694 15608 12174
rect 15714 12180 15752 12186
rect 15714 12174 15804 12180
rect 15714 12158 15792 12174
rect 15658 12135 15714 12144
rect 15948 11694 15976 12650
rect 16040 12102 16068 12650
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15672 9994 15700 11562
rect 16040 11354 16068 11562
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16132 11234 16160 12582
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11694 16252 12038
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16040 11206 16160 11234
rect 16040 10062 16068 11206
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16132 10606 16160 11018
rect 16224 10674 16252 11630
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10130 16160 10542
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15844 10056 15896 10062
rect 16028 10056 16080 10062
rect 15896 10016 15976 10044
rect 15844 9998 15896 10004
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15844 9512 15896 9518
rect 15842 9480 15844 9489
rect 15896 9480 15898 9489
rect 15842 9415 15898 9424
rect 15290 9344 15346 9353
rect 15290 9279 15346 9288
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 14924 8968 14976 8974
rect 14922 8936 14924 8945
rect 14976 8936 14978 8945
rect 14922 8871 14978 8880
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14936 7342 14964 7822
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14936 7002 14964 7278
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 15028 6934 15056 7822
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15016 6928 15068 6934
rect 14844 6854 14964 6882
rect 15016 6870 15068 6876
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14844 6186 14872 6734
rect 14936 6458 14964 6854
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14936 6361 14964 6394
rect 14922 6352 14978 6361
rect 14922 6287 14978 6296
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14936 6066 14964 6122
rect 14752 6038 14964 6066
rect 14936 5370 14964 6038
rect 15028 5710 15056 6870
rect 15212 6798 15240 7686
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15106 6488 15162 6497
rect 15106 6423 15162 6432
rect 15120 6322 15148 6423
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15014 5400 15070 5409
rect 14924 5364 14976 5370
rect 15014 5335 15070 5344
rect 14924 5306 14976 5312
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 15028 4690 15056 5335
rect 15120 5302 15148 6054
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 15212 5234 15240 6734
rect 15304 6662 15332 7754
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15396 6458 15424 7482
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15580 6225 15608 9046
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15672 8022 15700 8434
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15566 6216 15622 6225
rect 15566 6151 15622 6160
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 5370 15608 5646
rect 15672 5574 15700 7686
rect 15948 7546 15976 10016
rect 16028 9998 16080 10004
rect 16040 9674 16068 9998
rect 16040 9646 16160 9674
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 8498 16068 8910
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16040 7954 16068 8434
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16040 7342 16068 7890
rect 16132 7886 16160 9646
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16316 9178 16344 9454
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 7970 16344 8910
rect 16408 8090 16436 12786
rect 16592 12102 16620 13194
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12238 16804 12582
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16776 11082 16804 11698
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16868 10810 16896 13280
rect 16960 12986 16988 13330
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17420 12753 17448 13262
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17512 12850 17540 13126
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17406 12744 17462 12753
rect 17406 12679 17462 12688
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17144 12238 17172 12582
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9586 16712 9862
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16488 9512 16540 9518
rect 16486 9480 16488 9489
rect 16540 9480 16542 9489
rect 16486 9415 16542 9424
rect 16592 9160 16620 9522
rect 16592 9132 16712 9160
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16316 7942 16436 7970
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6798 16068 7278
rect 16132 7018 16160 7822
rect 16132 6990 16344 7018
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15948 6662 15976 6734
rect 15844 6656 15896 6662
rect 15750 6624 15806 6633
rect 15844 6598 15896 6604
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15750 6559 15806 6568
rect 15764 6322 15792 6559
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15856 6186 15884 6598
rect 15948 6254 15976 6598
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15764 5710 15792 5850
rect 15948 5760 15976 6190
rect 16040 5914 16068 6258
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15948 5732 16068 5760
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15580 4826 15608 5306
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15580 4622 15608 4762
rect 15764 4758 15792 5102
rect 15752 4752 15804 4758
rect 15672 4712 15752 4740
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15488 4434 15516 4558
rect 15566 4448 15622 4457
rect 15488 4406 15566 4434
rect 15566 4383 15622 4392
rect 14922 4312 14978 4321
rect 14922 4247 14924 4256
rect 14976 4247 14978 4256
rect 14924 4218 14976 4224
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 13924 3194 13952 3402
rect 14752 3194 14780 3878
rect 14936 3670 14964 4082
rect 15672 4010 15700 4712
rect 15752 4694 15804 4700
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14832 3528 14884 3534
rect 14830 3496 14832 3505
rect 14884 3496 14886 3505
rect 14830 3431 14886 3440
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15488 2990 15516 3878
rect 15672 3058 15700 3946
rect 15764 3738 15792 4082
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 3058 15792 3334
rect 15948 3058 15976 3878
rect 16040 3398 16068 5732
rect 16132 4146 16160 6258
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16224 5710 16252 6122
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16224 3534 16252 4150
rect 16316 3584 16344 6990
rect 16408 6798 16436 7942
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16408 4486 16436 6734
rect 16500 5710 16528 7822
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16396 4480 16448 4486
rect 16500 4457 16528 5646
rect 16396 4422 16448 4428
rect 16486 4448 16542 4457
rect 16486 4383 16542 4392
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3738 16436 4082
rect 16592 4026 16620 8978
rect 16684 6458 16712 9132
rect 16960 8906 16988 12038
rect 17328 11898 17356 12582
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17236 10810 17264 11086
rect 17512 10996 17540 12786
rect 17604 12442 17632 13262
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17788 12306 17816 12582
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17880 11150 17908 13670
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17420 10968 17540 10996
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17316 10668 17368 10674
rect 17420 10656 17448 10968
rect 17500 10804 17552 10810
rect 17552 10764 17632 10792
rect 17500 10746 17552 10752
rect 17368 10628 17448 10656
rect 17316 10610 17368 10616
rect 17328 9761 17356 10610
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17314 9752 17370 9761
rect 17314 9687 17370 9696
rect 17420 9586 17448 10406
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17144 9178 17172 9522
rect 17420 9178 17448 9522
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8974 17264 9046
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17052 7886 17080 8570
rect 17236 8362 17264 8910
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17328 8634 17356 8842
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17316 8492 17368 8498
rect 17420 8480 17448 8774
rect 17512 8566 17540 10542
rect 17604 9586 17632 10764
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17592 9104 17644 9110
rect 17590 9072 17592 9081
rect 17644 9072 17646 9081
rect 17590 9007 17646 9016
rect 17604 8974 17632 9007
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17604 8634 17632 8774
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17368 8452 17448 8480
rect 17316 8434 17368 8440
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16856 6316 16908 6322
rect 16908 6276 16988 6304
rect 16856 6258 16908 6264
rect 16960 6118 16988 6276
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16672 5568 16724 5574
rect 16776 5545 16804 5646
rect 16672 5510 16724 5516
rect 16762 5536 16818 5545
rect 16684 5302 16712 5510
rect 16762 5471 16818 5480
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16500 4010 16620 4026
rect 16488 4004 16620 4010
rect 16540 3998 16620 4004
rect 16488 3946 16540 3952
rect 16960 3942 16988 5714
rect 17052 4146 17080 7686
rect 17224 6656 17276 6662
rect 17328 6644 17356 8434
rect 17604 8294 17632 8570
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17604 7886 17632 8230
rect 17696 7954 17724 11018
rect 17880 10674 17908 11086
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17276 6616 17356 6644
rect 17224 6598 17276 6604
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17144 6089 17172 6122
rect 17130 6080 17186 6089
rect 17130 6015 17186 6024
rect 17144 5409 17172 6015
rect 17236 5914 17264 6598
rect 17314 6488 17370 6497
rect 17370 6446 17448 6474
rect 17314 6423 17370 6432
rect 17420 6322 17448 6446
rect 17590 6352 17646 6361
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17408 6316 17460 6322
rect 17590 6287 17592 6296
rect 17408 6258 17460 6264
rect 17644 6287 17646 6296
rect 17592 6258 17644 6264
rect 17328 6118 17356 6258
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17130 5400 17186 5409
rect 17130 5335 17186 5344
rect 17144 4622 17172 5335
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17132 4140 17184 4146
rect 17328 4128 17356 6054
rect 17696 5710 17724 7686
rect 17788 6458 17816 10542
rect 17972 10266 18000 16118
rect 18340 15570 18368 16186
rect 18800 16114 18828 21490
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19904 21146 19932 21422
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19260 19786 19288 20334
rect 19720 19854 19748 20538
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 17542 18920 18634
rect 19260 18290 19288 19722
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19440 19484 19446
rect 19892 19440 19944 19446
rect 19432 19382 19484 19388
rect 19890 19408 19892 19417
rect 20088 19428 20116 23122
rect 20166 23080 20222 23089
rect 20166 23015 20222 23024
rect 20180 22438 20208 23015
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20364 21622 20392 22918
rect 20548 22094 20576 27254
rect 20640 26994 20668 28018
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 21008 25786 21036 28562
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21284 26382 21312 26726
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21008 25758 21220 25786
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21100 25498 21128 25638
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 20824 23866 20852 24006
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20916 22982 20944 23734
rect 21008 23322 21036 24142
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 21008 22778 21036 23122
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 20548 22066 20668 22094
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20364 20534 20392 21558
rect 20640 20602 20668 22066
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20732 20074 20760 20742
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20548 20058 20760 20074
rect 20536 20052 20760 20058
rect 20588 20046 20760 20052
rect 20536 19994 20588 20000
rect 20824 19786 20852 20198
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 19944 19408 20116 19428
rect 19946 19400 20116 19408
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17338 18920 17478
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18340 15162 18368 15506
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18524 14958 18552 15302
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18064 13462 18092 13874
rect 18248 13870 18276 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12850 18092 13126
rect 18156 13002 18184 13262
rect 18234 13016 18290 13025
rect 18156 12974 18234 13002
rect 18234 12951 18290 12960
rect 18248 12850 18276 12951
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18064 12170 18092 12786
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 18156 11762 18184 12582
rect 18248 12434 18276 12786
rect 18340 12646 18368 13874
rect 18616 13784 18644 14447
rect 18708 14074 18736 14894
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 14074 18828 14214
rect 18892 14074 18920 14282
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18972 13875 19024 13881
rect 18972 13817 19024 13823
rect 18880 13796 18932 13802
rect 18616 13756 18880 13784
rect 18880 13738 18932 13744
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12850 18552 13330
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18708 12442 18736 12718
rect 18696 12436 18748 12442
rect 18248 12406 18552 12434
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18064 11121 18092 11154
rect 18050 11112 18106 11121
rect 18050 11047 18106 11056
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 9654 18092 10406
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17972 8634 18000 9046
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 8430 18092 9590
rect 18156 8566 18184 11018
rect 18340 10810 18368 11698
rect 18432 11354 18460 11698
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10130 18276 10678
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18340 9722 18368 10542
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 9104 18288 9110
rect 18234 9072 18236 9081
rect 18288 9072 18290 9081
rect 18234 9007 18290 9016
rect 18236 8968 18288 8974
rect 18432 8956 18460 11086
rect 18288 8928 18460 8956
rect 18236 8910 18288 8916
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18052 8424 18104 8430
rect 18248 8412 18276 8910
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 8566 18368 8774
rect 18328 8560 18380 8566
rect 18380 8508 18460 8514
rect 18328 8502 18460 8508
rect 18340 8486 18460 8502
rect 18052 8366 18104 8372
rect 18156 8384 18276 8412
rect 18328 8424 18380 8430
rect 18156 7970 18184 8384
rect 18328 8366 18380 8372
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18248 8090 18276 8230
rect 18340 8090 18368 8366
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18156 7942 18276 7970
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17972 6730 18000 7346
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17972 6322 18000 6666
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18064 6225 18092 6598
rect 18050 6216 18106 6225
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 17960 6180 18012 6186
rect 18050 6151 18106 6160
rect 17960 6122 18012 6128
rect 17880 6089 17908 6122
rect 17866 6080 17922 6089
rect 17866 6015 17922 6024
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17684 5704 17736 5710
rect 17498 5672 17554 5681
rect 17684 5646 17736 5652
rect 17498 5607 17554 5616
rect 17184 4100 17356 4128
rect 17132 4082 17184 4088
rect 16948 3936 17000 3942
rect 16946 3904 16948 3913
rect 17000 3904 17002 3913
rect 16946 3839 17002 3848
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16488 3596 16540 3602
rect 16316 3556 16488 3584
rect 16488 3538 16540 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16040 3126 16068 3334
rect 16316 3194 16344 3334
rect 16592 3194 16620 3470
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 17236 3058 17264 4100
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3602 17356 3878
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 17132 2984 17184 2990
rect 17420 2938 17448 4014
rect 17512 4010 17540 5607
rect 17880 4554 17908 5850
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17866 4448 17922 4457
rect 17866 4383 17922 4392
rect 17590 4176 17646 4185
rect 17880 4146 17908 4383
rect 17972 4282 18000 6122
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18064 5710 18092 6054
rect 18156 5710 18184 7414
rect 18248 6798 18276 7942
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 18064 4146 18092 5646
rect 18248 5642 18276 6734
rect 18328 6724 18380 6730
rect 18432 6712 18460 8486
rect 18524 7750 18552 12406
rect 18696 12378 18748 12384
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18708 11150 18736 12174
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 8838 18644 9522
rect 18708 9178 18736 11086
rect 18800 10198 18828 12854
rect 18984 11898 19012 13817
rect 19076 12434 19104 18158
rect 19352 16726 19380 18770
rect 19444 18698 19472 19382
rect 19890 19343 19946 19352
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20456 18358 20484 19654
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20456 17270 20484 18294
rect 20640 18086 20668 19654
rect 21008 19514 21036 20402
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16250 20024 16390
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19996 15434 20024 16186
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15162 20116 15982
rect 20364 15570 20392 16594
rect 20456 16590 20484 17206
rect 20640 17202 20668 18022
rect 20732 17882 20760 18158
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20824 17270 20852 18294
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20444 15564 20496 15570
rect 20548 15552 20576 17138
rect 20496 15524 20576 15552
rect 20444 15506 20496 15512
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20088 14618 20116 14894
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19168 12714 19196 14554
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19352 13258 19380 14418
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20088 13938 20116 14554
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19536 12442 19564 12718
rect 19524 12436 19576 12442
rect 19076 12406 19380 12434
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 10674 19104 10950
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19168 10588 19196 12106
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10742 19288 11086
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19168 10560 19288 10588
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18800 9761 18828 9930
rect 18786 9752 18842 9761
rect 18786 9687 18842 9696
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18800 9110 18828 9687
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18878 9072 18934 9081
rect 18984 9058 19012 9522
rect 18934 9030 19012 9058
rect 18878 9007 18934 9016
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18616 7954 18644 8774
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18380 6684 18460 6712
rect 18328 6666 18380 6672
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 18142 5536 18198 5545
rect 18142 5471 18198 5480
rect 18156 4486 18184 5471
rect 18234 4992 18290 5001
rect 18234 4927 18290 4936
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 17590 4111 17646 4120
rect 17868 4140 17920 4146
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17604 3534 17632 4111
rect 17868 4082 17920 4088
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17592 3528 17644 3534
rect 18064 3516 18092 4082
rect 18156 4049 18184 4422
rect 18248 4146 18276 4927
rect 18326 4176 18382 4185
rect 18236 4140 18288 4146
rect 18432 4146 18460 6684
rect 18524 6644 18552 7686
rect 18616 7392 18644 7890
rect 18800 7410 18828 8298
rect 18892 8090 18920 8366
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18696 7404 18748 7410
rect 18616 7364 18696 7392
rect 18696 7346 18748 7352
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18604 6656 18656 6662
rect 18524 6616 18604 6644
rect 18604 6598 18656 6604
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5914 18552 6190
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18616 5778 18644 6598
rect 18708 5846 18736 7346
rect 18800 6118 18828 7346
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4146 18644 4558
rect 18892 4146 18920 6870
rect 19168 4826 19196 9998
rect 19260 7426 19288 10560
rect 19352 9178 19380 12406
rect 19996 12434 20024 12786
rect 19524 12378 19576 12384
rect 19812 12406 20024 12434
rect 19812 12374 19840 12406
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19444 11150 19472 12310
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19522 11520 19578 11529
rect 19522 11455 19578 11464
rect 19536 11150 19564 11455
rect 19996 11354 20024 12106
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10810 19472 10950
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19444 10470 19472 10542
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 7546 19380 8842
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19260 7398 19380 7426
rect 19352 7206 19380 7398
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19260 6322 19288 6802
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19352 6202 19380 7142
rect 19260 6174 19380 6202
rect 19260 5522 19288 6174
rect 19338 5944 19394 5953
rect 19444 5914 19472 10406
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19812 9926 19840 9998
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9178 20024 9998
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19536 8294 19564 8434
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19996 8090 20024 8910
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19338 5879 19340 5888
rect 19392 5879 19394 5888
rect 19432 5908 19484 5914
rect 19340 5850 19392 5856
rect 19432 5850 19484 5856
rect 19432 5704 19484 5710
rect 19338 5672 19394 5681
rect 19394 5652 19432 5658
rect 19394 5646 19484 5652
rect 19394 5630 19472 5646
rect 19338 5607 19394 5616
rect 19260 5494 19472 5522
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18984 4282 19012 4694
rect 19444 4622 19472 5494
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18326 4111 18328 4120
rect 18236 4082 18288 4088
rect 18380 4111 18382 4120
rect 18420 4140 18472 4146
rect 18328 4082 18380 4088
rect 18420 4082 18472 4088
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18142 4040 18198 4049
rect 18142 3975 18198 3984
rect 18432 3942 18460 4082
rect 18892 4026 18920 4082
rect 18800 3998 18920 4026
rect 18984 4010 19012 4218
rect 19062 4176 19118 4185
rect 19118 4146 19196 4162
rect 19118 4140 19208 4146
rect 19118 4134 19156 4140
rect 19062 4111 19118 4120
rect 19156 4082 19208 4088
rect 19352 4078 19380 4490
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4146 20024 7890
rect 20088 6934 20116 12174
rect 20180 10810 20208 15302
rect 20364 15162 20392 15370
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20456 15094 20484 15506
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 21100 14482 21128 24006
rect 21192 21622 21220 25758
rect 21468 23322 21496 28966
rect 22756 28626 22784 31726
rect 22836 31272 22888 31278
rect 22836 31214 22888 31220
rect 22848 30938 22876 31214
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 21732 28484 21784 28490
rect 21732 28426 21784 28432
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21560 28082 21588 28358
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21560 23526 21588 28018
rect 21744 28014 21772 28426
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21652 26450 21680 27406
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21928 27130 21956 27338
rect 22112 27130 22140 28358
rect 22572 28014 22600 28358
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 27674 22600 27950
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 22100 27124 22152 27130
rect 22100 27066 22152 27072
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21652 26246 21680 26386
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21652 25362 21680 26182
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22020 25362 22048 25638
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 21652 24886 21680 25298
rect 21640 24880 21692 24886
rect 21640 24822 21692 24828
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22020 24206 22048 24550
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22112 24070 22140 25842
rect 22480 25498 22508 25842
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22204 24410 22232 24754
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21284 21486 21312 23122
rect 21560 23118 21588 23462
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21836 22234 21864 22374
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21284 21010 21312 21422
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21652 20942 21680 21558
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21192 19718 21220 20742
rect 21928 19990 21956 22918
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22020 21690 22048 22578
rect 22204 21894 22232 24074
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23526 22324 24006
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22296 21690 22324 23462
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21192 19514 21220 19654
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21376 17660 21404 19314
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 18834 21496 19178
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21928 18766 21956 19926
rect 22388 19786 22416 21966
rect 22480 21010 22508 23054
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22480 19922 22508 20946
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22388 19446 22416 19722
rect 22480 19514 22508 19858
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22480 19378 22508 19450
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22204 18970 22232 19314
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17746 21680 18022
rect 21928 17882 21956 18566
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21456 17672 21508 17678
rect 21284 17632 21456 17660
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20732 13462 20760 13942
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20732 12850 20760 13398
rect 21100 13326 21128 14282
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20916 12986 20944 13262
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20180 9178 20208 9658
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8294 20208 8774
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20180 6254 20208 8230
rect 20272 7954 20300 11154
rect 20364 11150 20392 12038
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20364 9586 20392 11086
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20364 8634 20392 8910
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20180 4146 20208 5646
rect 20456 5642 20484 11290
rect 20732 11082 20760 12786
rect 21100 11694 21128 13262
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 9518 20576 10542
rect 20640 9926 20668 11018
rect 20720 10668 20772 10674
rect 20824 10656 20852 11630
rect 20772 10628 20852 10656
rect 20720 10610 20772 10616
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20548 5642 20576 9114
rect 20640 8974 20668 9862
rect 20732 9518 20760 10610
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8090 20668 8910
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 18972 4004 19024 4010
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18800 3738 18828 3998
rect 18972 3946 19024 3952
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18892 3738 18920 3878
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18236 3528 18288 3534
rect 18064 3488 18236 3516
rect 17592 3470 17644 3476
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19444 3482 19472 4082
rect 20180 3602 20208 4082
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 19248 3470 19300 3476
rect 19260 3194 19288 3470
rect 19352 3454 19472 3482
rect 19352 3194 19380 3454
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3194 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20180 3194 20208 3538
rect 20824 3534 20852 7346
rect 21192 6186 21220 15098
rect 21284 15026 21312 17632
rect 21456 17614 21508 17620
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 15042 21496 17478
rect 21744 16658 21772 17614
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 22112 16574 22140 18634
rect 22572 17270 22600 20470
rect 22664 20058 22692 24210
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22756 22778 22784 22986
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22204 16794 22232 17070
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22664 16726 22692 16934
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 21836 16546 22140 16574
rect 21836 16114 21864 16546
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21560 15473 21588 15506
rect 21546 15464 21602 15473
rect 21546 15399 21602 15408
rect 21272 15020 21324 15026
rect 21468 15014 21680 15042
rect 21272 14962 21324 14968
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21272 11144 21324 11150
rect 21270 11112 21272 11121
rect 21324 11112 21326 11121
rect 21270 11047 21326 11056
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21284 9722 21312 10542
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21376 8634 21404 14894
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21468 10810 21496 13194
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21560 10606 21588 12174
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 9654 21588 10542
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21376 7546 21404 8366
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21468 7342 21496 9454
rect 21652 8344 21680 15014
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11354 21772 12038
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21744 8974 21772 9318
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21560 8316 21680 8344
rect 21560 8090 21588 8316
rect 21836 8276 21864 16050
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14890 21956 14962
rect 22204 14890 22232 15438
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22020 14482 22048 14826
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22296 14056 22324 16390
rect 22388 15026 22416 16594
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15706 22508 15846
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22664 15162 22692 15914
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22204 14028 22324 14056
rect 22560 14068 22612 14074
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22112 13734 22140 13874
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12850 21956 13330
rect 22006 13288 22062 13297
rect 22006 13223 22062 13232
rect 22020 13190 22048 13223
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22204 13138 22232 14028
rect 22560 14010 22612 14016
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22296 13530 22324 13806
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22006 13016 22062 13025
rect 22006 12951 22062 12960
rect 22020 12850 22048 12951
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21928 12306 21956 12786
rect 22112 12442 22140 13126
rect 22204 13110 22324 13138
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12646 22232 12786
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22098 12336 22154 12345
rect 21916 12300 21968 12306
rect 22098 12271 22154 12280
rect 21916 12242 21968 12248
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 10266 21956 12038
rect 22020 11694 22048 12174
rect 22112 11898 22140 12271
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22008 11688 22060 11694
rect 22060 11636 22140 11642
rect 22008 11630 22140 11636
rect 22020 11614 22140 11630
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11150 22048 11494
rect 22112 11150 22140 11614
rect 22296 11354 22324 13110
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22098 10976 22154 10985
rect 22098 10911 22154 10920
rect 22112 10810 22140 10911
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 22098 10704 22154 10713
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21928 9722 21956 9930
rect 22020 9926 22048 10678
rect 22098 10639 22100 10648
rect 22152 10639 22154 10648
rect 22100 10610 22152 10616
rect 22204 10198 22232 11018
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22296 10266 22324 10610
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22192 10192 22244 10198
rect 22388 10146 22416 13942
rect 22572 13734 22600 14010
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22480 13025 22508 13670
rect 22572 13394 22600 13670
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22466 13016 22522 13025
rect 22466 12951 22522 12960
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22480 11898 22508 12310
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22572 11778 22600 13330
rect 22664 12102 22692 14894
rect 22756 14074 22784 21490
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22848 16998 22876 18158
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22848 16590 22876 16934
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22940 15978 22968 39374
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23768 38962 23796 39238
rect 24044 38962 24072 40122
rect 24228 39914 24256 41550
rect 24412 40662 24440 42094
rect 24400 40656 24452 40662
rect 24400 40598 24452 40604
rect 24216 39908 24268 39914
rect 24216 39850 24268 39856
rect 24228 38962 24256 39850
rect 24412 39506 24440 40598
rect 24952 40384 25004 40390
rect 24952 40326 25004 40332
rect 24584 39976 24636 39982
rect 24584 39918 24636 39924
rect 24400 39500 24452 39506
rect 24400 39442 24452 39448
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24320 39098 24348 39238
rect 24308 39092 24360 39098
rect 24308 39034 24360 39040
rect 24412 38962 24440 39442
rect 24596 39098 24624 39918
rect 24964 39370 24992 40326
rect 25872 40044 25924 40050
rect 25872 39986 25924 39992
rect 25228 39840 25280 39846
rect 25228 39782 25280 39788
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 24952 39364 25004 39370
rect 24952 39306 25004 39312
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 25044 39024 25096 39030
rect 25044 38966 25096 38972
rect 23756 38956 23808 38962
rect 23756 38898 23808 38904
rect 24032 38956 24084 38962
rect 24032 38898 24084 38904
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 23572 38888 23624 38894
rect 23572 38830 23624 38836
rect 23584 38554 23612 38830
rect 24492 38820 24544 38826
rect 24492 38762 24544 38768
rect 24504 38706 24532 38762
rect 24504 38678 24900 38706
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 24872 38010 24900 38678
rect 25056 38486 25084 38966
rect 25240 38894 25268 39782
rect 25228 38888 25280 38894
rect 25228 38830 25280 38836
rect 25332 38758 25360 39782
rect 25884 39642 25912 39986
rect 26700 39840 26752 39846
rect 26700 39782 26752 39788
rect 26792 39840 26844 39846
rect 26792 39782 26844 39788
rect 25872 39636 25924 39642
rect 25872 39578 25924 39584
rect 26148 39500 26200 39506
rect 26148 39442 26200 39448
rect 26160 38894 26188 39442
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 26344 38758 26372 39238
rect 26712 38894 26740 39782
rect 26804 39506 26832 39782
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 26896 39030 26924 42094
rect 27068 42016 27120 42022
rect 27068 41958 27120 41964
rect 27080 41414 27108 41958
rect 27080 41386 27384 41414
rect 26976 40044 27028 40050
rect 26976 39986 27028 39992
rect 26884 39024 26936 39030
rect 26884 38966 26936 38972
rect 26792 38956 26844 38962
rect 26792 38898 26844 38904
rect 26700 38888 26752 38894
rect 26700 38830 26752 38836
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 26332 38752 26384 38758
rect 26332 38694 26384 38700
rect 25044 38480 25096 38486
rect 25044 38422 25096 38428
rect 25412 38412 25464 38418
rect 25412 38354 25464 38360
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 24768 37732 24820 37738
rect 24768 37674 24820 37680
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 23768 36802 23796 37062
rect 23860 36922 23888 37198
rect 23940 37120 23992 37126
rect 23940 37062 23992 37068
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23952 36854 23980 37062
rect 23940 36848 23992 36854
rect 23768 36774 23888 36802
rect 23940 36790 23992 36796
rect 23664 36712 23716 36718
rect 23664 36654 23716 36660
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 23124 36242 23152 36518
rect 23676 36378 23704 36654
rect 23664 36372 23716 36378
rect 23664 36314 23716 36320
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 23584 35698 23612 36178
rect 23756 36168 23808 36174
rect 23756 36110 23808 36116
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23584 34610 23612 35634
rect 23768 35290 23796 36110
rect 23860 36106 23888 36774
rect 23952 36174 23980 36790
rect 24412 36378 24440 37198
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 23940 36168 23992 36174
rect 23940 36110 23992 36116
rect 24032 36168 24084 36174
rect 24032 36110 24084 36116
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23756 35284 23808 35290
rect 23756 35226 23808 35232
rect 24044 34950 24072 36110
rect 24780 36106 24808 37674
rect 25332 37262 25360 37810
rect 25424 37330 25452 38354
rect 25412 37324 25464 37330
rect 25412 37266 25464 37272
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 25056 36922 25084 37062
rect 25424 36922 25452 37266
rect 25688 37256 25740 37262
rect 25688 37198 25740 37204
rect 25044 36916 25096 36922
rect 25044 36858 25096 36864
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24872 36310 24900 36518
rect 24860 36304 24912 36310
rect 24860 36246 24912 36252
rect 24872 36174 24900 36246
rect 25240 36174 25268 36654
rect 25424 36242 25452 36858
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24952 36168 25004 36174
rect 24952 36110 25004 36116
rect 25228 36168 25280 36174
rect 25228 36110 25280 36116
rect 24768 36100 24820 36106
rect 24596 36060 24768 36088
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 24492 34944 24544 34950
rect 24492 34886 24544 34892
rect 24044 34610 24072 34886
rect 24504 34678 24532 34886
rect 24492 34672 24544 34678
rect 24492 34614 24544 34620
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 23480 34400 23532 34406
rect 23480 34342 23532 34348
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23492 34066 23520 34342
rect 23584 34066 23612 34342
rect 23480 34060 23532 34066
rect 23480 34002 23532 34008
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 23032 29238 23060 33866
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23400 33590 23428 33798
rect 23584 33590 23612 33866
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23676 32910 23704 34546
rect 24044 34354 24072 34546
rect 23952 34326 24072 34354
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23860 33114 23888 33254
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23584 31754 23612 32846
rect 23676 32366 23704 32846
rect 23664 32360 23716 32366
rect 23664 32302 23716 32308
rect 23492 31726 23612 31754
rect 23388 30592 23440 30598
rect 23388 30534 23440 30540
rect 23204 30048 23256 30054
rect 23400 30002 23428 30534
rect 23492 30138 23520 31726
rect 23572 31408 23624 31414
rect 23572 31350 23624 31356
rect 23584 30274 23612 31350
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23860 30920 23888 31078
rect 23768 30892 23888 30920
rect 23768 30802 23796 30892
rect 23952 30818 23980 34326
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 32298 24440 33934
rect 24596 33862 24624 36060
rect 24768 36042 24820 36048
rect 24676 34060 24728 34066
rect 24676 34002 24728 34008
rect 24768 34060 24820 34066
rect 24768 34002 24820 34008
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24596 32824 24624 33798
rect 24688 33114 24716 34002
rect 24780 33386 24808 34002
rect 24872 33998 24900 36110
rect 24964 35834 24992 36110
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 25056 34202 25084 35022
rect 25240 34678 25268 36110
rect 25700 35086 25728 37198
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 25976 36174 26004 36722
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25976 35766 26004 36110
rect 25964 35760 26016 35766
rect 25964 35702 26016 35708
rect 25976 35290 26004 35702
rect 26056 35624 26108 35630
rect 26056 35566 26108 35572
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 25688 35080 25740 35086
rect 25688 35022 25740 35028
rect 25228 34672 25280 34678
rect 25228 34614 25280 34620
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24768 33380 24820 33386
rect 24768 33322 24820 33328
rect 24676 33108 24728 33114
rect 24676 33050 24728 33056
rect 24872 32910 24900 33934
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24676 32836 24728 32842
rect 24596 32796 24676 32824
rect 24400 32292 24452 32298
rect 24400 32234 24452 32240
rect 24032 31816 24084 31822
rect 24032 31758 24084 31764
rect 23756 30796 23808 30802
rect 23756 30738 23808 30744
rect 23860 30790 23980 30818
rect 23584 30258 23704 30274
rect 23572 30252 23704 30258
rect 23624 30246 23704 30252
rect 23572 30194 23624 30200
rect 23492 30122 23612 30138
rect 23492 30116 23624 30122
rect 23492 30110 23572 30116
rect 23572 30058 23624 30064
rect 23256 29996 23336 30002
rect 23204 29990 23336 29996
rect 23216 29974 23336 29990
rect 23400 29974 23612 30002
rect 23020 29232 23072 29238
rect 23020 29174 23072 29180
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23032 28218 23060 28494
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23124 27606 23152 28154
rect 23308 27878 23336 29974
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23124 26518 23152 27542
rect 23112 26512 23164 26518
rect 23112 26454 23164 26460
rect 23308 26246 23336 27814
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23492 26926 23520 27474
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23492 26450 23520 26862
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 23308 25906 23336 26182
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23492 25786 23520 26386
rect 23584 26382 23612 29974
rect 23676 28218 23704 30246
rect 23860 28626 23888 30790
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23952 30394 23980 30670
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 23848 28620 23900 28626
rect 23848 28562 23900 28568
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28218 23796 28358
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23584 26042 23612 26182
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23664 25832 23716 25838
rect 23216 25498 23244 25774
rect 23492 25758 23612 25786
rect 23664 25774 23716 25780
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23204 25492 23256 25498
rect 23204 25434 23256 25440
rect 23492 25226 23520 25638
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23492 24886 23520 25162
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 23584 24274 23612 25758
rect 23676 25498 23704 25774
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23664 25152 23716 25158
rect 23768 25140 23796 27270
rect 23860 26042 23888 28562
rect 24044 28558 24072 31758
rect 24596 31754 24624 32796
rect 24676 32778 24728 32784
rect 24872 32026 24900 32846
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24964 31890 24992 32710
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24124 30796 24176 30802
rect 24124 30738 24176 30744
rect 24136 29714 24164 30738
rect 24504 30190 24532 31622
rect 24872 31482 24900 31758
rect 25056 31482 25084 33594
rect 25700 32842 25728 35022
rect 26068 34746 26096 35566
rect 26056 34740 26108 34746
rect 26056 34682 26108 34688
rect 26068 33998 26096 34682
rect 26056 33992 26108 33998
rect 26056 33934 26108 33940
rect 26240 33652 26292 33658
rect 26240 33594 26292 33600
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 26252 32434 26280 33594
rect 26344 33046 26372 38694
rect 26712 35986 26740 38830
rect 26804 37194 26832 38898
rect 26792 37188 26844 37194
rect 26792 37130 26844 37136
rect 26804 36106 26832 37130
rect 26792 36100 26844 36106
rect 26792 36042 26844 36048
rect 26712 35958 26832 35986
rect 26424 35760 26476 35766
rect 26424 35702 26476 35708
rect 26436 35154 26464 35702
rect 26804 35494 26832 35958
rect 26792 35488 26844 35494
rect 26792 35430 26844 35436
rect 26424 35148 26476 35154
rect 26424 35090 26476 35096
rect 26804 34542 26832 35430
rect 26792 34536 26844 34542
rect 26792 34478 26844 34484
rect 26896 34406 26924 38966
rect 26988 38758 27016 39986
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 27160 38276 27212 38282
rect 27160 38218 27212 38224
rect 26976 37664 27028 37670
rect 26976 37606 27028 37612
rect 26988 37330 27016 37606
rect 26976 37324 27028 37330
rect 26976 37266 27028 37272
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 26976 36576 27028 36582
rect 26976 36518 27028 36524
rect 26988 36242 27016 36518
rect 26976 36236 27028 36242
rect 26976 36178 27028 36184
rect 27080 35834 27108 36722
rect 27068 35828 27120 35834
rect 27068 35770 27120 35776
rect 26884 34400 26936 34406
rect 26884 34342 26936 34348
rect 27068 34400 27120 34406
rect 27068 34342 27120 34348
rect 26608 33992 26660 33998
rect 26608 33934 26660 33940
rect 26424 33924 26476 33930
rect 26424 33866 26476 33872
rect 26436 33658 26464 33866
rect 26424 33652 26476 33658
rect 26424 33594 26476 33600
rect 26436 33386 26464 33594
rect 26516 33584 26568 33590
rect 26516 33526 26568 33532
rect 26424 33380 26476 33386
rect 26424 33322 26476 33328
rect 26528 33114 26556 33526
rect 26620 33454 26648 33934
rect 26896 33522 26924 34342
rect 27080 34066 27108 34342
rect 27068 34060 27120 34066
rect 27068 34002 27120 34008
rect 26884 33516 26936 33522
rect 26884 33458 26936 33464
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 26516 33108 26568 33114
rect 26516 33050 26568 33056
rect 26332 33040 26384 33046
rect 26332 32982 26384 32988
rect 26424 32904 26476 32910
rect 26424 32846 26476 32852
rect 26436 32502 26464 32846
rect 26620 32570 26648 33390
rect 27172 32910 27200 38218
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 27264 32978 27292 34546
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 26608 32564 26660 32570
rect 26608 32506 26660 32512
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 25148 32026 25176 32302
rect 26884 32292 26936 32298
rect 26884 32234 26936 32240
rect 25136 32020 25188 32026
rect 25136 31962 25188 31968
rect 26896 31754 26924 32234
rect 27172 32026 27200 32846
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 27264 31906 27292 32914
rect 27080 31878 27292 31906
rect 27080 31754 27108 31878
rect 26424 31748 26476 31754
rect 26424 31690 26476 31696
rect 26712 31726 26924 31754
rect 26988 31726 27108 31754
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 24400 30184 24452 30190
rect 24400 30126 24452 30132
rect 24492 30184 24544 30190
rect 24492 30126 24544 30132
rect 24412 29850 24440 30126
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 24504 29646 24532 30126
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24676 28960 24728 28966
rect 24676 28902 24728 28908
rect 24032 28552 24084 28558
rect 24032 28494 24084 28500
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24412 27674 24440 28018
rect 24688 28014 24716 28902
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 24584 27872 24636 27878
rect 24584 27814 24636 27820
rect 24596 27674 24624 27814
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 24688 27538 24716 27950
rect 24676 27532 24728 27538
rect 24676 27474 24728 27480
rect 24964 27470 24992 27950
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24412 27130 24440 27406
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24308 26920 24360 26926
rect 24308 26862 24360 26868
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 24044 25294 24072 26182
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 23716 25112 23796 25140
rect 23664 25094 23716 25100
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 23216 23202 23244 23598
rect 23032 23174 23244 23202
rect 23032 22098 23060 23174
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23400 22409 23428 22578
rect 23386 22400 23442 22409
rect 23386 22335 23442 22344
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21010 23152 21286
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23308 20602 23336 21490
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23124 18426 23152 18702
rect 23400 18426 23428 21966
rect 23492 20602 23520 24006
rect 23676 22778 23704 25094
rect 23756 24676 23808 24682
rect 23756 24618 23808 24624
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23768 22658 23796 24618
rect 24228 23322 24256 25230
rect 24320 24070 24348 26862
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 24032 23044 24084 23050
rect 24032 22986 24084 22992
rect 24124 23044 24176 23050
rect 24124 22986 24176 22992
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 23584 22630 23796 22658
rect 23584 21554 23612 22630
rect 23756 22568 23808 22574
rect 23940 22568 23992 22574
rect 23756 22510 23808 22516
rect 23846 22536 23902 22545
rect 23768 22094 23796 22510
rect 23940 22510 23992 22516
rect 23846 22471 23902 22480
rect 23676 22066 23796 22094
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23492 18222 23520 18770
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 23124 15706 23152 17614
rect 23492 16658 23520 18158
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23492 15570 23520 16050
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23202 15464 23258 15473
rect 23202 15399 23204 15408
rect 23256 15399 23258 15408
rect 23204 15370 23256 15376
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22848 14074 22876 14486
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 23112 13932 23164 13938
rect 23164 13892 23244 13920
rect 23112 13874 23164 13880
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22756 13326 22784 13738
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22480 11750 22600 11778
rect 22480 11558 22508 11750
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 10656 22508 11494
rect 22572 10985 22600 11562
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 11150 22692 11494
rect 22756 11286 22784 13262
rect 22848 12782 22876 13738
rect 23216 13326 23244 13892
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23400 13734 23428 13806
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12782 22968 13126
rect 23032 12986 23060 13262
rect 23216 12986 23244 13262
rect 23400 13161 23428 13262
rect 23386 13152 23442 13161
rect 23386 13087 23442 13096
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 22756 11150 22784 11222
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22848 11014 22876 11494
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22836 11008 22888 11014
rect 22558 10976 22614 10985
rect 22836 10950 22888 10956
rect 22558 10911 22614 10920
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22652 10668 22704 10674
rect 22480 10628 22652 10656
rect 22652 10610 22704 10616
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 10198 22508 10474
rect 22192 10134 22244 10140
rect 22296 10118 22416 10146
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21928 8498 21956 9522
rect 22020 9110 22048 9522
rect 22112 9450 22140 9998
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22296 9178 22324 10118
rect 22376 9988 22428 9994
rect 22376 9930 22428 9936
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22388 9178 22416 9930
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22480 9110 22508 9930
rect 22664 9450 22692 10610
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22756 9194 22784 10134
rect 22940 10062 22968 10746
rect 23032 10713 23060 11086
rect 23124 10810 23152 12378
rect 23216 11558 23244 12922
rect 23400 12850 23428 13087
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23492 12646 23520 13806
rect 23584 13530 23612 20334
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23584 12442 23612 13330
rect 23676 13258 23704 22066
rect 23860 22030 23888 22471
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23952 21486 23980 22510
rect 24044 21690 24072 22986
rect 24136 22710 24164 22986
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23952 20398 23980 21422
rect 24044 20874 24072 21626
rect 24032 20868 24084 20874
rect 24032 20810 24084 20816
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23768 18970 23796 19450
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23768 18426 23796 18906
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23768 16250 23796 18362
rect 24044 18358 24072 20810
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23860 16046 23888 16390
rect 24504 16250 24532 22986
rect 24596 21146 24624 24142
rect 25056 23866 25084 31418
rect 26436 31414 26464 31690
rect 26424 31408 26476 31414
rect 26424 31350 26476 31356
rect 25872 31272 25924 31278
rect 25872 31214 25924 31220
rect 25884 30938 25912 31214
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30938 26096 31078
rect 25872 30932 25924 30938
rect 25872 30874 25924 30880
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26252 29850 26280 30534
rect 26436 30326 26464 31350
rect 26712 30666 26740 31726
rect 26792 31340 26844 31346
rect 26792 31282 26844 31288
rect 26700 30660 26752 30666
rect 26700 30602 26752 30608
rect 26712 30394 26740 30602
rect 26700 30388 26752 30394
rect 26700 30330 26752 30336
rect 26424 30320 26476 30326
rect 26424 30262 26476 30268
rect 26424 30184 26476 30190
rect 26424 30126 26476 30132
rect 26240 29844 26292 29850
rect 26240 29786 26292 29792
rect 26252 28558 26280 29786
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26344 29170 26372 29446
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26252 28218 26280 28494
rect 25320 28212 25372 28218
rect 25320 28154 25372 28160
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 25332 27402 25360 28154
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25332 26926 25360 27338
rect 26252 27130 26280 28154
rect 26344 27538 26372 29106
rect 26332 27532 26384 27538
rect 26332 27474 26384 27480
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25332 25974 25360 26862
rect 25412 26852 25464 26858
rect 25412 26794 25464 26800
rect 25424 26314 25452 26794
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25424 25974 25452 26250
rect 25320 25968 25372 25974
rect 25320 25910 25372 25916
rect 25412 25968 25464 25974
rect 25412 25910 25464 25916
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25148 24614 25176 25230
rect 25700 24954 25728 25298
rect 25884 25158 25912 25774
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25884 24682 25912 25094
rect 26068 24682 26096 25638
rect 26160 24954 26188 25842
rect 26436 25786 26464 30126
rect 26804 28966 26832 31282
rect 26792 28960 26844 28966
rect 26792 28902 26844 28908
rect 26252 25758 26464 25786
rect 26252 25430 26280 25758
rect 26332 25696 26384 25702
rect 26332 25638 26384 25644
rect 26700 25696 26752 25702
rect 26700 25638 26752 25644
rect 26344 25430 26372 25638
rect 26712 25498 26740 25638
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26332 25424 26384 25430
rect 26332 25366 26384 25372
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26148 24948 26200 24954
rect 26148 24890 26200 24896
rect 26160 24818 26188 24890
rect 26252 24818 26280 25230
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 25872 24676 25924 24682
rect 25872 24618 25924 24624
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 25056 22094 25084 23802
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25608 22778 25636 23054
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25884 22710 25912 23054
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25332 22234 25360 22374
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 24964 22066 25084 22094
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24872 20330 24900 21898
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24872 19854 24900 20266
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18358 24716 18566
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24688 15366 24716 16390
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24228 15162 24256 15302
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23860 13326 23888 13670
rect 24688 13326 24716 13942
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24780 13326 24808 13670
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23940 13184 23992 13190
rect 23768 13144 23940 13172
rect 23768 12986 23796 13144
rect 23940 13126 23992 13132
rect 24228 12986 24256 13262
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23308 11762 23336 12242
rect 24320 12170 24348 12786
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23018 10704 23074 10713
rect 23018 10639 23074 10648
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22664 9166 22784 9194
rect 22664 9110 22692 9166
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22020 8634 22048 8910
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22480 8566 22508 9046
rect 22664 8922 22692 9046
rect 22572 8894 22692 8922
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 21652 8248 21864 8276
rect 22100 8288 22152 8294
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20916 3448 20944 5578
rect 21652 4214 21680 8248
rect 22100 8230 22152 8236
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21836 7546 21864 7822
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21928 6458 21956 7890
rect 22112 7818 22140 8230
rect 22204 7954 22232 8366
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 22296 8090 22324 8298
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22204 7274 22232 7890
rect 22468 7472 22520 7478
rect 22572 7460 22600 8894
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 7818 22692 8774
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22756 7546 22784 7686
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22520 7432 22600 7460
rect 22468 7414 22520 7420
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22480 6458 22508 7414
rect 22848 7410 22876 9386
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22112 5778 22140 6190
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22572 5574 22600 6190
rect 22848 5574 22876 7346
rect 22940 6118 22968 9862
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22572 5030 22600 5510
rect 23032 5114 23060 8978
rect 23308 5914 23336 11698
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10674 23520 11222
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 8634 23428 9590
rect 23492 9042 23520 10610
rect 23952 9722 23980 10610
rect 24320 10538 24348 10950
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23492 8498 23520 8774
rect 23676 8634 23704 9454
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24412 9178 24440 9318
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24504 8922 24532 11086
rect 24596 10810 24624 13262
rect 24688 11898 24716 13262
rect 24964 12889 24992 22066
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25056 20942 25084 21966
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25148 18358 25176 22102
rect 25700 22030 25728 22578
rect 25780 22500 25832 22506
rect 25780 22442 25832 22448
rect 25792 22094 25820 22442
rect 25884 22216 25912 22646
rect 25964 22228 26016 22234
rect 25884 22188 25964 22216
rect 25964 22170 26016 22176
rect 26068 22166 26096 24618
rect 26160 22642 26188 24754
rect 26252 23594 26280 24754
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 26148 22636 26200 22642
rect 26200 22596 26280 22624
rect 26148 22578 26200 22584
rect 26252 22234 26280 22596
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26056 22160 26108 22166
rect 26056 22102 26108 22108
rect 25792 22066 25912 22094
rect 25884 22030 25912 22066
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25884 21350 25912 21966
rect 26252 21622 26280 22170
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25502 20632 25558 20641
rect 25502 20567 25558 20576
rect 25516 19417 25544 20567
rect 25778 20088 25834 20097
rect 25778 20023 25834 20032
rect 25792 19990 25820 20023
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25502 19408 25558 19417
rect 25502 19343 25504 19352
rect 25556 19343 25558 19352
rect 25700 19334 25728 19790
rect 25792 19446 25820 19926
rect 25884 19854 25912 21286
rect 25976 21146 26004 21286
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25504 19314 25556 19320
rect 25608 19306 25728 19334
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25608 18290 25636 19306
rect 25884 18970 25912 19790
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25608 17678 25636 18226
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25700 17202 25728 18294
rect 25792 17746 25820 18702
rect 25884 18086 25912 18702
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25884 17882 25912 18022
rect 25872 17876 25924 17882
rect 25872 17818 25924 17824
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25700 16590 25728 17138
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25700 16182 25728 16526
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25240 14618 25268 14894
rect 25332 14618 25360 14894
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25976 14550 26004 20742
rect 26068 19922 26096 20878
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26160 19786 26188 20198
rect 26344 19990 26372 21966
rect 26332 19984 26384 19990
rect 26332 19926 26384 19932
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26160 19514 26188 19722
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26160 18766 26188 19110
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26056 18080 26108 18086
rect 26160 18068 26188 18702
rect 26252 18426 26280 19314
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26240 18080 26292 18086
rect 26160 18040 26240 18068
rect 26056 18022 26108 18028
rect 26240 18022 26292 18028
rect 26068 17134 26096 18022
rect 26252 17814 26280 18022
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26344 17678 26372 18906
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26344 16590 26372 17614
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26344 15502 26372 16526
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26252 14890 26280 15302
rect 26240 14884 26292 14890
rect 26240 14826 26292 14832
rect 25964 14544 26016 14550
rect 25964 14486 26016 14492
rect 26252 14414 26280 14826
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 25424 13530 25452 14350
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25502 13016 25558 13025
rect 25502 12951 25504 12960
rect 25556 12951 25558 12960
rect 25504 12922 25556 12928
rect 24950 12880 25006 12889
rect 24950 12815 25006 12824
rect 25608 12646 25636 13330
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 26160 12889 26188 13126
rect 26240 12912 26292 12918
rect 26146 12880 26202 12889
rect 25872 12844 25924 12850
rect 26240 12854 26292 12860
rect 26146 12815 26202 12824
rect 25872 12786 25924 12792
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24688 11354 24716 11698
rect 24780 11626 24808 12038
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24964 11218 24992 11698
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 24584 10804 24636 10810
rect 24584 10746 24636 10752
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24688 9722 24716 10610
rect 25056 10538 25084 10950
rect 25148 10606 25176 12242
rect 25608 11762 25636 12582
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25884 10810 25912 12786
rect 26056 12776 26108 12782
rect 26056 12718 26108 12724
rect 26068 12306 26096 12718
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 26252 12170 26280 12854
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26344 12374 26372 12650
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26240 12164 26292 12170
rect 26240 12106 26292 12112
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25044 10532 25096 10538
rect 25044 10474 25096 10480
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 25148 9674 25176 10542
rect 24688 9178 24716 9658
rect 25148 9646 25268 9674
rect 25240 9518 25268 9646
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24780 9110 24808 9318
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24504 8894 24624 8922
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23664 8492 23716 8498
rect 24032 8492 24084 8498
rect 23716 8452 24032 8480
rect 23664 8434 23716 8440
rect 24032 8434 24084 8440
rect 23492 8090 23520 8434
rect 24596 8430 24624 8894
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24596 8294 24624 8366
rect 24584 8288 24636 8294
rect 24584 8230 24636 8236
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 24596 7954 24624 8230
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24320 7410 24348 7686
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24596 7342 24624 7890
rect 24688 7410 24716 7890
rect 24872 7818 24900 9318
rect 25240 9042 25268 9454
rect 25516 9382 25544 10610
rect 26344 10606 26372 12310
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24964 8634 24992 8842
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24964 7546 24992 8298
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23492 6866 23520 7142
rect 24596 6866 24624 7278
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 24596 5846 24624 6802
rect 24688 5914 24716 7346
rect 25056 7002 25084 7414
rect 25240 7290 25268 8978
rect 26160 8974 26188 9318
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25332 7546 25360 8366
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25700 7886 25728 8230
rect 25884 8090 25912 8774
rect 26344 8362 26372 8774
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25318 7304 25374 7313
rect 25240 7262 25318 7290
rect 25318 7239 25374 7248
rect 25332 7206 25360 7239
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 25608 6866 25636 7142
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23400 5234 23428 5578
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22940 5086 23060 5114
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 22296 4010 22324 4558
rect 22848 4486 22876 5034
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4214 22876 4422
rect 22836 4208 22888 4214
rect 22940 4185 22968 5086
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 23032 4622 23060 4966
rect 23400 4826 23428 5170
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 23124 4282 23152 4422
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23204 4208 23256 4214
rect 22836 4150 22888 4156
rect 22926 4176 22982 4185
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 20996 3460 21048 3466
rect 20916 3420 20996 3448
rect 20996 3402 21048 3408
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 21008 3126 21036 3402
rect 20996 3120 21048 3126
rect 18694 3088 18750 3097
rect 20996 3062 21048 3068
rect 22204 3058 22232 3674
rect 22296 3466 22324 3946
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3670 22508 3878
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 18694 3023 18696 3032
rect 18748 3023 18750 3032
rect 22192 3052 22244 3058
rect 18696 2994 18748 3000
rect 22192 2994 22244 3000
rect 17184 2932 17448 2938
rect 17132 2926 17448 2932
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 13176 2916 13228 2922
rect 17144 2910 17448 2926
rect 18972 2916 19024 2922
rect 13176 2858 13228 2864
rect 18972 2858 19024 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8680 2650 8708 2858
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 10704 2514 10732 2790
rect 18984 2650 19012 2858
rect 22296 2854 22324 3402
rect 22480 3126 22508 3470
rect 22572 3398 22600 4082
rect 22848 3738 22876 4150
rect 23204 4150 23256 4156
rect 22926 4111 22982 4120
rect 22940 3738 22968 4111
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22940 3058 22968 3674
rect 23216 3534 23244 4150
rect 23492 4010 23520 5646
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23676 4010 23704 4966
rect 23768 4622 23796 5510
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23848 4072 23900 4078
rect 23952 4060 23980 4694
rect 24032 4684 24084 4690
rect 24032 4626 24084 4632
rect 23900 4032 23980 4060
rect 23848 4014 23900 4020
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23308 3210 23336 3878
rect 23584 3670 23612 3946
rect 23952 3738 23980 4032
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23308 3182 23428 3210
rect 23492 3194 23520 3402
rect 23584 3194 23612 3606
rect 24044 3534 24072 4626
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24412 3602 24440 4558
rect 24688 4282 24716 5646
rect 25240 5234 25268 5714
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25608 5030 25636 6802
rect 25700 6662 25728 7346
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 25884 7206 25912 7278
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25700 6458 25728 6598
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26068 5098 26096 5646
rect 26436 5574 26464 23666
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26804 22778 26832 23054
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26528 15706 26556 21830
rect 26988 20806 27016 31726
rect 27080 31686 27108 31726
rect 27068 31680 27120 31686
rect 27068 31622 27120 31628
rect 27356 28082 27384 41386
rect 27448 39506 27476 42230
rect 30932 42016 30984 42022
rect 30932 41958 30984 41964
rect 30944 41414 30972 41958
rect 31220 41818 31248 43386
rect 32600 43314 32628 43658
rect 33048 43648 33100 43654
rect 33048 43590 33100 43596
rect 33060 43450 33088 43590
rect 33048 43444 33100 43450
rect 33048 43386 33100 43392
rect 32588 43308 32640 43314
rect 32588 43250 32640 43256
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31208 41812 31260 41818
rect 31208 41754 31260 41760
rect 30852 41386 30972 41414
rect 27436 39500 27488 39506
rect 27436 39442 27488 39448
rect 27896 39500 27948 39506
rect 27896 39442 27948 39448
rect 28908 39500 28960 39506
rect 28908 39442 28960 39448
rect 27528 38956 27580 38962
rect 27528 38898 27580 38904
rect 27540 38010 27568 38898
rect 27908 38894 27936 39442
rect 28540 39296 28592 39302
rect 28540 39238 28592 39244
rect 28724 39296 28776 39302
rect 28724 39238 28776 39244
rect 27896 38888 27948 38894
rect 27896 38830 27948 38836
rect 28264 38888 28316 38894
rect 28264 38830 28316 38836
rect 28276 38554 28304 38830
rect 28264 38548 28316 38554
rect 28264 38490 28316 38496
rect 28552 38350 28580 39238
rect 28736 39030 28764 39238
rect 28724 39024 28776 39030
rect 28724 38966 28776 38972
rect 28920 38418 28948 39442
rect 29460 39364 29512 39370
rect 29460 39306 29512 39312
rect 30380 39364 30432 39370
rect 30380 39306 30432 39312
rect 29472 38894 29500 39306
rect 29460 38888 29512 38894
rect 29460 38830 29512 38836
rect 29368 38820 29420 38826
rect 29368 38762 29420 38768
rect 29380 38554 29408 38762
rect 29368 38548 29420 38554
rect 29368 38490 29420 38496
rect 28908 38412 28960 38418
rect 28736 38372 28908 38400
rect 28540 38344 28592 38350
rect 28540 38286 28592 38292
rect 28632 38276 28684 38282
rect 28632 38218 28684 38224
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 27448 36582 27476 37810
rect 27540 37330 27568 37946
rect 27712 37936 27764 37942
rect 27712 37878 27764 37884
rect 27528 37324 27580 37330
rect 27528 37266 27580 37272
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 27632 36582 27660 37062
rect 27724 36922 27752 37878
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27816 37466 27844 37742
rect 28644 37738 28672 38218
rect 28736 37942 28764 38372
rect 28908 38354 28960 38360
rect 29472 38350 29500 38830
rect 29552 38752 29604 38758
rect 29552 38694 29604 38700
rect 29564 38418 29592 38694
rect 29552 38412 29604 38418
rect 29552 38354 29604 38360
rect 29460 38344 29512 38350
rect 29460 38286 29512 38292
rect 28724 37936 28776 37942
rect 28724 37878 28776 37884
rect 27896 37732 27948 37738
rect 27896 37674 27948 37680
rect 28632 37732 28684 37738
rect 28632 37674 28684 37680
rect 27804 37460 27856 37466
rect 27804 37402 27856 37408
rect 27712 36916 27764 36922
rect 27712 36858 27764 36864
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27528 36576 27580 36582
rect 27528 36518 27580 36524
rect 27620 36576 27672 36582
rect 27620 36518 27672 36524
rect 27448 34490 27476 36518
rect 27540 35494 27568 36518
rect 27632 35494 27660 36518
rect 27908 35766 27936 37674
rect 28644 37398 28672 37674
rect 29472 37670 29500 38286
rect 30392 38282 30420 39306
rect 29920 38276 29972 38282
rect 29920 38218 29972 38224
rect 30380 38276 30432 38282
rect 30380 38218 30432 38224
rect 29932 38010 29960 38218
rect 30104 38208 30156 38214
rect 30104 38150 30156 38156
rect 29920 38004 29972 38010
rect 29920 37946 29972 37952
rect 30116 37874 30144 38150
rect 30104 37868 30156 37874
rect 30104 37810 30156 37816
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 29460 37664 29512 37670
rect 29460 37606 29512 37612
rect 28632 37392 28684 37398
rect 28632 37334 28684 37340
rect 29012 36854 29040 37606
rect 30012 37392 30064 37398
rect 30012 37334 30064 37340
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 28184 36378 28212 36722
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 28092 35834 28120 35974
rect 28080 35828 28132 35834
rect 28080 35770 28132 35776
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 28184 35698 28212 36314
rect 29012 36174 29040 36790
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 30024 36106 30052 37334
rect 30116 36106 30144 37810
rect 30196 36780 30248 36786
rect 30196 36722 30248 36728
rect 29368 36100 29420 36106
rect 29368 36042 29420 36048
rect 30012 36100 30064 36106
rect 30012 36042 30064 36048
rect 30104 36100 30156 36106
rect 30104 36042 30156 36048
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28552 35698 28580 35974
rect 29380 35766 29408 36042
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29656 35834 29684 35974
rect 29644 35828 29696 35834
rect 30024 35816 30052 36042
rect 29644 35770 29696 35776
rect 29932 35788 30052 35816
rect 29368 35760 29420 35766
rect 29368 35702 29420 35708
rect 28172 35692 28224 35698
rect 28172 35634 28224 35640
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 27896 35624 27948 35630
rect 27896 35566 27948 35572
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27620 35488 27672 35494
rect 27620 35430 27672 35436
rect 27540 34610 27568 35430
rect 27632 34950 27660 35430
rect 27620 34944 27672 34950
rect 27620 34886 27672 34892
rect 27908 34746 27936 35566
rect 27896 34740 27948 34746
rect 27896 34682 27948 34688
rect 28448 34672 28500 34678
rect 28448 34614 28500 34620
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27448 34462 27568 34490
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27448 33572 27476 33866
rect 27540 33674 27568 34462
rect 28460 34202 28488 34614
rect 28448 34196 28500 34202
rect 28448 34138 28500 34144
rect 27540 33646 27660 33674
rect 28552 33658 28580 35634
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 27528 33584 27580 33590
rect 27448 33544 27528 33572
rect 27528 33526 27580 33532
rect 27632 33402 27660 33646
rect 27896 33652 27948 33658
rect 27896 33594 27948 33600
rect 28540 33652 28592 33658
rect 28540 33594 28592 33600
rect 27540 33374 27660 33402
rect 27540 31414 27568 33374
rect 27908 32570 27936 33594
rect 28644 33454 28672 35566
rect 29828 33856 29880 33862
rect 29828 33798 29880 33804
rect 29840 33590 29868 33798
rect 29828 33584 29880 33590
rect 29828 33526 29880 33532
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 28632 33448 28684 33454
rect 28632 33390 28684 33396
rect 28644 33114 28672 33390
rect 28632 33108 28684 33114
rect 28632 33050 28684 33056
rect 27896 32564 27948 32570
rect 27896 32506 27948 32512
rect 28644 31414 28672 33050
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 28632 31408 28684 31414
rect 28632 31350 28684 31356
rect 27436 31272 27488 31278
rect 27436 31214 27488 31220
rect 27448 30394 27476 31214
rect 27436 30388 27488 30394
rect 27436 30330 27488 30336
rect 27540 30326 27568 31350
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28276 30802 28304 31282
rect 29012 30938 29040 33458
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 29748 31822 29776 32302
rect 29932 31822 29960 35788
rect 30116 31822 30144 36042
rect 30208 34746 30236 36722
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30576 35834 30604 36110
rect 30656 36032 30708 36038
rect 30656 35974 30708 35980
rect 30668 35834 30696 35974
rect 30564 35828 30616 35834
rect 30564 35770 30616 35776
rect 30656 35828 30708 35834
rect 30656 35770 30708 35776
rect 30196 34740 30248 34746
rect 30196 34682 30248 34688
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29920 31816 29972 31822
rect 29920 31758 29972 31764
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 29552 31680 29604 31686
rect 29552 31622 29604 31628
rect 29564 31278 29592 31622
rect 30012 31408 30064 31414
rect 30012 31350 30064 31356
rect 29552 31272 29604 31278
rect 29552 31214 29604 31220
rect 29644 31204 29696 31210
rect 29644 31146 29696 31152
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 29288 30870 29316 31078
rect 29276 30864 29328 30870
rect 29276 30806 29328 30812
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 29460 30728 29512 30734
rect 29460 30670 29512 30676
rect 27804 30660 27856 30666
rect 27804 30602 27856 30608
rect 27816 30394 27844 30602
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 28078 30424 28134 30433
rect 27804 30388 27856 30394
rect 28078 30359 28134 30368
rect 27804 30330 27856 30336
rect 27528 30320 27580 30326
rect 27528 30262 27580 30268
rect 27896 30252 27948 30258
rect 27896 30194 27948 30200
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27632 29850 27660 29990
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27436 29640 27488 29646
rect 27436 29582 27488 29588
rect 27448 29170 27476 29582
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27528 29096 27580 29102
rect 27448 29044 27528 29050
rect 27448 29038 27580 29044
rect 27448 29022 27568 29038
rect 27448 28558 27476 29022
rect 27632 28966 27660 29446
rect 27908 29170 27936 30194
rect 27896 29164 27948 29170
rect 27896 29106 27948 29112
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27632 28422 27660 28902
rect 27908 28422 27936 29106
rect 27620 28416 27672 28422
rect 27540 28376 27620 28404
rect 27344 28076 27396 28082
rect 27344 28018 27396 28024
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 27080 24614 27108 24822
rect 27172 24750 27200 25094
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 27540 24682 27568 28376
rect 27896 28416 27948 28422
rect 27620 28358 27672 28364
rect 27816 28376 27896 28404
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27724 24954 27752 25230
rect 27712 24948 27764 24954
rect 27712 24890 27764 24896
rect 27816 24818 27844 28376
rect 27896 28358 27948 28364
rect 28092 28082 28120 30359
rect 29104 30326 29132 30534
rect 29472 30326 29500 30670
rect 29092 30320 29144 30326
rect 29092 30262 29144 30268
rect 29460 30320 29512 30326
rect 29460 30262 29512 30268
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 29012 29306 29040 30126
rect 29104 30036 29132 30262
rect 29656 30258 29684 31146
rect 30024 30938 30052 31350
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29184 30184 29236 30190
rect 29736 30184 29788 30190
rect 29236 30132 29736 30138
rect 29184 30126 29788 30132
rect 29196 30110 29776 30126
rect 29104 30008 29316 30036
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29104 28762 29132 29106
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27528 24676 27580 24682
rect 27528 24618 27580 24624
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27908 22094 27936 27814
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 28368 26926 28396 27406
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28368 26586 28396 26862
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28276 26042 28304 26318
rect 28448 26240 28500 26246
rect 28448 26182 28500 26188
rect 28264 26036 28316 26042
rect 28264 25978 28316 25984
rect 28460 25906 28488 26182
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28552 24614 28580 27950
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28736 26926 28764 27814
rect 29196 26994 29224 28426
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 28724 26920 28776 26926
rect 28724 26862 28776 26868
rect 29104 26518 29132 26930
rect 29092 26512 29144 26518
rect 29092 26454 29144 26460
rect 29196 26432 29224 26930
rect 29288 26790 29316 30008
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29748 28218 29776 28358
rect 29932 28218 29960 28494
rect 29736 28212 29788 28218
rect 29736 28154 29788 28160
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29368 28144 29420 28150
rect 29368 28086 29420 28092
rect 29380 27402 29408 28086
rect 30024 27402 30052 30874
rect 30116 30394 30144 31758
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 30208 30258 30236 34682
rect 30576 34134 30604 35770
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 30760 34202 30788 34546
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30564 34128 30616 34134
rect 30564 34070 30616 34076
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 30564 32224 30616 32230
rect 30564 32166 30616 32172
rect 30576 32026 30604 32166
rect 30668 32026 30696 32302
rect 30564 32020 30616 32026
rect 30564 31962 30616 31968
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30472 31816 30524 31822
rect 30472 31758 30524 31764
rect 30484 31346 30512 31758
rect 30576 31754 30604 31962
rect 30852 31754 30880 41386
rect 31208 37732 31260 37738
rect 31208 37674 31260 37680
rect 31220 36922 31248 37674
rect 31208 36916 31260 36922
rect 31208 36858 31260 36864
rect 31116 36576 31168 36582
rect 31116 36518 31168 36524
rect 31128 36242 31156 36518
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 31116 36032 31168 36038
rect 31116 35974 31168 35980
rect 31128 35766 31156 35974
rect 31220 35766 31248 36858
rect 31312 36530 31340 43046
rect 32600 42226 32628 43250
rect 34060 43104 34112 43110
rect 34060 43046 34112 43052
rect 35532 43104 35584 43110
rect 35532 43046 35584 43052
rect 34072 42362 34100 43046
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34980 42628 35032 42634
rect 34980 42570 35032 42576
rect 34796 42560 34848 42566
rect 34796 42502 34848 42508
rect 34060 42356 34112 42362
rect 34060 42298 34112 42304
rect 34808 42294 34836 42502
rect 34796 42288 34848 42294
rect 34796 42230 34848 42236
rect 32588 42220 32640 42226
rect 32588 42162 32640 42168
rect 34704 42152 34756 42158
rect 34704 42094 34756 42100
rect 34716 41818 34744 42094
rect 34704 41812 34756 41818
rect 34704 41754 34756 41760
rect 32036 41608 32088 41614
rect 32036 41550 32088 41556
rect 33140 41608 33192 41614
rect 33140 41550 33192 41556
rect 34520 41608 34572 41614
rect 34520 41550 34572 41556
rect 32048 39506 32076 41550
rect 33152 41274 33180 41550
rect 33140 41268 33192 41274
rect 33140 41210 33192 41216
rect 34532 40526 34560 41550
rect 34716 41414 34744 41754
rect 34624 41386 34744 41414
rect 34624 41138 34652 41386
rect 34612 41132 34664 41138
rect 34612 41074 34664 41080
rect 34808 41070 34836 42230
rect 34992 42158 35020 42570
rect 35544 42362 35572 43046
rect 35532 42356 35584 42362
rect 35532 42298 35584 42304
rect 35716 42220 35768 42226
rect 35716 42162 35768 42168
rect 34980 42152 35032 42158
rect 34980 42094 35032 42100
rect 35532 42152 35584 42158
rect 35532 42094 35584 42100
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35348 41812 35400 41818
rect 35348 41754 35400 41760
rect 34888 41540 34940 41546
rect 34888 41482 34940 41488
rect 34900 41274 34928 41482
rect 34888 41268 34940 41274
rect 34888 41210 34940 41216
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 34520 40520 34572 40526
rect 34520 40462 34572 40468
rect 34612 40384 34664 40390
rect 34612 40326 34664 40332
rect 32312 39976 32364 39982
rect 32312 39918 32364 39924
rect 34520 39976 34572 39982
rect 34520 39918 34572 39924
rect 31668 39500 31720 39506
rect 31668 39442 31720 39448
rect 31760 39500 31812 39506
rect 31760 39442 31812 39448
rect 32036 39500 32088 39506
rect 32036 39442 32088 39448
rect 31680 39370 31708 39442
rect 31668 39364 31720 39370
rect 31668 39306 31720 39312
rect 31772 39098 31800 39442
rect 32220 39296 32272 39302
rect 32324 39284 32352 39918
rect 32772 39840 32824 39846
rect 32772 39782 32824 39788
rect 32496 39500 32548 39506
rect 32496 39442 32548 39448
rect 32272 39256 32352 39284
rect 32220 39238 32272 39244
rect 31760 39092 31812 39098
rect 31760 39034 31812 39040
rect 31576 38412 31628 38418
rect 31576 38354 31628 38360
rect 31484 38208 31536 38214
rect 31484 38150 31536 38156
rect 31496 37874 31524 38150
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 31312 36502 31524 36530
rect 31392 36236 31444 36242
rect 31392 36178 31444 36184
rect 31116 35760 31168 35766
rect 31116 35702 31168 35708
rect 31208 35760 31260 35766
rect 31208 35702 31260 35708
rect 31404 35698 31432 36178
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31404 35562 31432 35634
rect 31392 35556 31444 35562
rect 31392 35498 31444 35504
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30944 34202 30972 34546
rect 31024 34468 31076 34474
rect 31024 34410 31076 34416
rect 30932 34196 30984 34202
rect 30932 34138 30984 34144
rect 31036 34134 31064 34410
rect 31404 34202 31432 35498
rect 31116 34196 31168 34202
rect 31116 34138 31168 34144
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31024 34128 31076 34134
rect 31024 34070 31076 34076
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30944 32434 30972 32710
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 31024 32224 31076 32230
rect 31024 32166 31076 32172
rect 31036 31822 31064 32166
rect 31128 31822 31156 34138
rect 31392 33992 31444 33998
rect 31392 33934 31444 33940
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 31220 32842 31248 33798
rect 31404 33658 31432 33934
rect 31392 33652 31444 33658
rect 31392 33594 31444 33600
rect 31404 32910 31432 33594
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31208 32836 31260 32842
rect 31208 32778 31260 32784
rect 31392 32768 31444 32774
rect 31392 32710 31444 32716
rect 31404 32502 31432 32710
rect 31208 32496 31260 32502
rect 31208 32438 31260 32444
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 31220 32298 31248 32438
rect 31300 32360 31352 32366
rect 31300 32302 31352 32308
rect 31208 32292 31260 32298
rect 31208 32234 31260 32240
rect 31312 31822 31340 32302
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 30576 31726 30696 31754
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30472 31340 30524 31346
rect 30472 31282 30524 31288
rect 30392 30734 30420 31282
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30196 28484 30248 28490
rect 30196 28426 30248 28432
rect 29368 27396 29420 27402
rect 29368 27338 29420 27344
rect 30012 27396 30064 27402
rect 30012 27338 30064 27344
rect 29460 27328 29512 27334
rect 29460 27270 29512 27276
rect 29472 26994 29500 27270
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29460 26512 29512 26518
rect 29460 26454 29512 26460
rect 29196 26404 29408 26432
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 29012 25974 29040 26318
rect 29184 26308 29236 26314
rect 29184 26250 29236 26256
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 29196 25838 29224 26250
rect 29276 26240 29328 26246
rect 29276 26182 29328 26188
rect 29288 25974 29316 26182
rect 29276 25968 29328 25974
rect 29276 25910 29328 25916
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29012 25430 29040 25638
rect 29196 25498 29224 25774
rect 29184 25492 29236 25498
rect 29184 25434 29236 25440
rect 29000 25424 29052 25430
rect 29000 25366 29052 25372
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29196 23322 29224 24006
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 28092 22642 28120 23054
rect 29000 23044 29052 23050
rect 29000 22986 29052 22992
rect 29012 22778 29040 22986
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 28080 22636 28132 22642
rect 28080 22578 28132 22584
rect 28092 22234 28120 22578
rect 28080 22228 28132 22234
rect 28080 22170 28132 22176
rect 28540 22228 28592 22234
rect 28540 22170 28592 22176
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 27908 22066 28028 22094
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 27816 19718 27844 21898
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27724 19310 27752 19654
rect 27816 19446 27844 19654
rect 27804 19440 27856 19446
rect 27804 19382 27856 19388
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26620 16658 26648 18566
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27080 17202 27108 18158
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27356 17542 27384 17818
rect 27436 17808 27488 17814
rect 27620 17808 27672 17814
rect 27488 17768 27620 17796
rect 27436 17750 27488 17756
rect 27620 17750 27672 17756
rect 27528 17672 27580 17678
rect 27896 17672 27948 17678
rect 27580 17632 27896 17660
rect 27528 17614 27580 17620
rect 27896 17614 27948 17620
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27804 17536 27856 17542
rect 27804 17478 27856 17484
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 27632 16794 27660 17478
rect 27816 17338 27844 17478
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26620 15570 26648 16594
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26528 14550 26556 15438
rect 26712 15094 26740 16050
rect 26700 15088 26752 15094
rect 26700 15030 26752 15036
rect 26516 14544 26568 14550
rect 26516 14486 26568 14492
rect 26896 13734 26924 16186
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26988 15706 27016 16050
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 26988 14346 27016 15030
rect 27172 14618 27200 16594
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27264 14346 27292 15846
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 15094 27568 15302
rect 27816 15094 27844 15370
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27816 14482 27844 15030
rect 27436 14476 27488 14482
rect 27436 14418 27488 14424
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26988 13530 27016 14282
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27448 13394 27476 14418
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 28000 13258 28028 22066
rect 28092 21554 28120 22170
rect 28552 22030 28580 22170
rect 28816 22160 28868 22166
rect 28816 22102 28868 22108
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28828 21962 28856 22102
rect 28920 22094 28948 22170
rect 29104 22098 29132 22918
rect 28920 22066 28994 22094
rect 28966 22032 28994 22066
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 28954 22026 29006 22032
rect 28954 21968 29006 21974
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28632 21956 28684 21962
rect 28632 21898 28684 21904
rect 28816 21956 28868 21962
rect 28816 21898 28868 21904
rect 28276 21690 28304 21898
rect 28644 21690 28672 21898
rect 29196 21894 29224 22918
rect 29276 22636 29328 22642
rect 29380 22624 29408 26404
rect 29472 26042 29500 26454
rect 29564 26450 29592 26930
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29460 26036 29512 26042
rect 29460 25978 29512 25984
rect 29564 25974 29592 26386
rect 29552 25968 29604 25974
rect 29552 25910 29604 25916
rect 29564 25498 29592 25910
rect 29656 25702 29684 27066
rect 30208 27062 30236 28426
rect 30472 28416 30524 28422
rect 30472 28358 30524 28364
rect 30484 28218 30512 28358
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 30576 28014 30604 28494
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30668 27470 30696 31726
rect 30748 31748 30800 31754
rect 30852 31726 30972 31754
rect 30748 31690 30800 31696
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30196 27056 30248 27062
rect 30196 26998 30248 27004
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29748 26518 29776 26930
rect 29736 26512 29788 26518
rect 29736 26454 29788 26460
rect 29748 25906 29776 26454
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 30484 26042 30512 26386
rect 30472 26036 30524 26042
rect 30472 25978 30524 25984
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 29748 25702 29776 25842
rect 29644 25696 29696 25702
rect 29644 25638 29696 25644
rect 29736 25696 29788 25702
rect 29736 25638 29788 25644
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 29552 24336 29604 24342
rect 29552 24278 29604 24284
rect 29564 23866 29592 24278
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29748 23798 29776 25638
rect 30024 24262 30420 24290
rect 30024 24206 30052 24262
rect 30392 24206 30420 24262
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 29736 23792 29788 23798
rect 29736 23734 29788 23740
rect 29932 23730 29960 24142
rect 30116 24070 30144 24142
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29328 22596 29408 22624
rect 29276 22578 29328 22584
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28080 21548 28132 21554
rect 28356 21548 28408 21554
rect 28080 21490 28132 21496
rect 28276 21508 28356 21536
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28184 20466 28212 20946
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 28276 19922 28304 21508
rect 28356 21490 28408 21496
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28644 20942 28672 21286
rect 28736 21146 28764 21490
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28920 21078 28948 21490
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29196 21146 29224 21286
rect 29184 21140 29236 21146
rect 29184 21082 29236 21088
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28552 20602 28580 20878
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 28368 20058 28396 20402
rect 28644 20058 28672 20878
rect 28828 20618 28856 20878
rect 28828 20590 29224 20618
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28908 20324 28960 20330
rect 28908 20266 28960 20272
rect 28920 20058 28948 20266
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28276 19825 28304 19858
rect 28262 19816 28318 19825
rect 28262 19751 28318 19760
rect 28264 19508 28316 19514
rect 28368 19496 28396 19994
rect 29012 19854 29040 20402
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28816 19780 28868 19786
rect 28816 19722 28868 19728
rect 28828 19514 28856 19722
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 28316 19468 28396 19496
rect 28816 19508 28868 19514
rect 28264 19450 28316 19456
rect 28816 19450 28868 19456
rect 29012 18698 29040 19654
rect 29104 19514 29132 20334
rect 29196 19718 29224 20590
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 29000 18692 29052 18698
rect 29000 18634 29052 18640
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29196 17678 29224 18226
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29196 17202 29224 17614
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29288 16182 29316 22578
rect 29564 22030 29592 23054
rect 29656 22642 29684 23462
rect 29828 23044 29880 23050
rect 29828 22986 29880 22992
rect 29840 22778 29868 22986
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29826 22672 29882 22681
rect 29644 22636 29696 22642
rect 29826 22607 29828 22616
rect 29644 22578 29696 22584
rect 29880 22607 29882 22616
rect 29828 22578 29880 22584
rect 29828 22500 29880 22506
rect 29828 22442 29880 22448
rect 29840 22030 29868 22442
rect 29932 22234 29960 23666
rect 30012 23316 30064 23322
rect 30116 23304 30144 23666
rect 30300 23526 30328 24142
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30484 23866 30512 24006
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23322 30328 23462
rect 30064 23276 30144 23304
rect 30012 23258 30064 23264
rect 30116 22574 30144 23276
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30484 23186 30512 23666
rect 30472 23180 30524 23186
rect 30472 23122 30524 23128
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30208 22624 30236 22918
rect 30484 22642 30512 23122
rect 30668 22642 30696 24006
rect 30380 22636 30432 22642
rect 30208 22596 30380 22624
rect 30104 22568 30156 22574
rect 30104 22510 30156 22516
rect 29920 22228 29972 22234
rect 29920 22170 29972 22176
rect 30300 22030 30328 22596
rect 30380 22578 30432 22584
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 29564 21350 29592 21966
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 30012 21072 30064 21078
rect 30012 21014 30064 21020
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29552 20868 29604 20874
rect 29552 20810 29604 20816
rect 29564 20466 29592 20810
rect 29840 20806 29868 20946
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29840 20602 29868 20742
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29564 20210 29592 20402
rect 29826 20360 29882 20369
rect 29826 20295 29828 20304
rect 29880 20295 29882 20304
rect 29920 20324 29972 20330
rect 29828 20266 29880 20272
rect 29920 20266 29972 20272
rect 29380 20182 29592 20210
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29380 19990 29408 20182
rect 29368 19984 29420 19990
rect 29368 19926 29420 19932
rect 29748 19922 29776 20198
rect 29932 19990 29960 20266
rect 30024 20058 30052 21014
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30392 20482 30420 20878
rect 30300 20466 30420 20482
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30288 20460 30420 20466
rect 30340 20454 30420 20460
rect 30288 20402 30340 20408
rect 30116 20058 30144 20402
rect 30208 20346 30236 20402
rect 30484 20346 30512 22578
rect 30576 22506 30604 22578
rect 30564 22500 30616 22506
rect 30564 22442 30616 22448
rect 30760 22030 30788 31690
rect 30840 28144 30892 28150
rect 30840 28086 30892 28092
rect 30852 27878 30880 28086
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30852 23866 30880 24142
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 30748 22024 30800 22030
rect 30748 21966 30800 21972
rect 30760 21010 30788 21966
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 30576 20641 30604 20742
rect 30562 20632 30618 20641
rect 30562 20567 30618 20576
rect 30208 20318 30512 20346
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 29920 19984 29972 19990
rect 29920 19926 29972 19932
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29932 19514 29960 19926
rect 30378 19816 30434 19825
rect 30012 19780 30064 19786
rect 30378 19751 30434 19760
rect 30012 19722 30064 19728
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29276 16176 29328 16182
rect 29276 16118 29328 16124
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 29104 13938 29132 15914
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 29288 15706 29316 15846
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29380 15502 29408 18634
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 29564 17338 29592 17614
rect 29656 17542 29684 18226
rect 30024 17814 30052 19722
rect 30392 19378 30420 19751
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30852 18834 30880 21286
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 30116 17882 30144 18226
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30104 17876 30156 17882
rect 30104 17818 30156 17824
rect 30012 17808 30064 17814
rect 30012 17750 30064 17756
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 30024 17082 30052 17478
rect 30116 17218 30144 17614
rect 30208 17338 30236 18158
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 30392 17814 30420 18022
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30300 17626 30328 17682
rect 30300 17598 30420 17626
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30116 17190 30236 17218
rect 30208 17134 30236 17190
rect 30104 17128 30156 17134
rect 30024 17076 30104 17082
rect 30024 17070 30156 17076
rect 30196 17128 30248 17134
rect 30196 17070 30248 17076
rect 30024 17054 30144 17070
rect 30116 16794 30144 17054
rect 30392 16998 30420 17598
rect 30472 17196 30524 17202
rect 30472 17138 30524 17144
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 29552 16584 29604 16590
rect 30392 16538 30420 16934
rect 30484 16590 30512 17138
rect 30564 17128 30616 17134
rect 30564 17070 30616 17076
rect 29552 16526 29604 16532
rect 29564 16114 29592 16526
rect 30208 16522 30420 16538
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30196 16516 30420 16522
rect 30248 16510 30420 16516
rect 30196 16458 30248 16464
rect 30576 16454 30604 17070
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 29644 16448 29696 16454
rect 29644 16390 29696 16396
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30564 16448 30616 16454
rect 30564 16390 30616 16396
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29656 16046 29684 16390
rect 30116 16046 30144 16390
rect 30286 16144 30342 16153
rect 30286 16079 30288 16088
rect 30340 16079 30342 16088
rect 30288 16050 30340 16056
rect 30668 16046 30696 16526
rect 30840 16516 30892 16522
rect 30840 16458 30892 16464
rect 30852 16182 30880 16458
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 29644 16040 29696 16046
rect 29644 15982 29696 15988
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30656 16040 30708 16046
rect 30840 16040 30892 16046
rect 30656 15982 30708 15988
rect 30838 16008 30840 16017
rect 30892 16008 30894 16017
rect 30116 15706 30144 15982
rect 30838 15943 30894 15952
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30024 14028 30236 14056
rect 30024 13938 30052 14028
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 29184 13864 29236 13870
rect 29184 13806 29236 13812
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 29196 13190 29224 13806
rect 29736 13796 29788 13802
rect 29736 13738 29788 13744
rect 29748 13326 29776 13738
rect 30116 13326 30144 13874
rect 30208 13462 30236 14028
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30196 13456 30248 13462
rect 30196 13398 30248 13404
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30300 13274 30328 13806
rect 30484 13802 30512 14418
rect 30944 14074 30972 31726
rect 31128 31414 31156 31758
rect 31116 31408 31168 31414
rect 31116 31350 31168 31356
rect 31404 31346 31432 32438
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31024 29028 31076 29034
rect 31024 28970 31076 28976
rect 31036 28558 31064 28970
rect 31220 28626 31248 29106
rect 31208 28620 31260 28626
rect 31208 28562 31260 28568
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 31206 28248 31262 28257
rect 31206 28183 31262 28192
rect 31220 28150 31248 28183
rect 31208 28144 31260 28150
rect 31208 28086 31260 28092
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31128 27878 31156 28018
rect 31116 27872 31168 27878
rect 31116 27814 31168 27820
rect 31128 26586 31156 27814
rect 31312 26858 31340 30670
rect 31390 28520 31446 28529
rect 31390 28455 31392 28464
rect 31444 28455 31446 28464
rect 31392 28426 31444 28432
rect 31300 26852 31352 26858
rect 31300 26794 31352 26800
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31404 24410 31432 24754
rect 31392 24404 31444 24410
rect 31392 24346 31444 24352
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 31404 22778 31432 22918
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 31128 20942 31156 22034
rect 31220 20942 31248 22374
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31036 20058 31064 20878
rect 31220 20097 31248 20878
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31312 20369 31340 20402
rect 31298 20360 31354 20369
rect 31298 20295 31354 20304
rect 31206 20088 31262 20097
rect 31024 20052 31076 20058
rect 31206 20023 31262 20032
rect 31024 19994 31076 20000
rect 31116 19168 31168 19174
rect 31116 19110 31168 19116
rect 31128 18834 31156 19110
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 31024 15972 31076 15978
rect 31024 15914 31076 15920
rect 31036 15706 31064 15914
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30944 13938 30972 14010
rect 31128 14006 31156 17546
rect 31392 16992 31444 16998
rect 31392 16934 31444 16940
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31312 16017 31340 16050
rect 31298 16008 31354 16017
rect 31404 15994 31432 16934
rect 31496 16538 31524 36502
rect 31588 36174 31616 38354
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 31680 36378 31708 36858
rect 31668 36372 31720 36378
rect 31668 36314 31720 36320
rect 31576 36168 31628 36174
rect 31576 36110 31628 36116
rect 31588 35714 31616 36110
rect 32128 36032 32180 36038
rect 32128 35974 32180 35980
rect 32140 35834 32168 35974
rect 31760 35828 31812 35834
rect 31760 35770 31812 35776
rect 32128 35828 32180 35834
rect 32128 35770 32180 35776
rect 31668 35760 31720 35766
rect 31588 35708 31668 35714
rect 31588 35702 31720 35708
rect 31588 35686 31708 35702
rect 31772 35086 31800 35770
rect 32324 35698 32352 39256
rect 32404 38956 32456 38962
rect 32404 38898 32456 38904
rect 32416 38554 32444 38898
rect 32508 38826 32536 39442
rect 32784 38894 32812 39782
rect 34532 39642 34560 39918
rect 34520 39636 34572 39642
rect 34520 39578 34572 39584
rect 34624 39438 34652 40326
rect 34704 39840 34756 39846
rect 34808 39794 34836 41006
rect 34900 40934 34928 41210
rect 35360 41070 35388 41754
rect 35440 41472 35492 41478
rect 35440 41414 35492 41420
rect 35348 41064 35400 41070
rect 35348 41006 35400 41012
rect 34888 40928 34940 40934
rect 34888 40870 34940 40876
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35256 40452 35308 40458
rect 35452 40440 35480 41414
rect 35544 40730 35572 42094
rect 35624 42084 35676 42090
rect 35624 42026 35676 42032
rect 35636 41614 35664 42026
rect 35624 41608 35676 41614
rect 35624 41550 35676 41556
rect 35728 41274 35756 42162
rect 36096 41818 36124 43726
rect 36820 43716 36872 43722
rect 36820 43658 36872 43664
rect 36452 43240 36504 43246
rect 36452 43182 36504 43188
rect 36464 42566 36492 43182
rect 36832 42702 36860 43658
rect 36820 42696 36872 42702
rect 36820 42638 36872 42644
rect 36452 42560 36504 42566
rect 36452 42502 36504 42508
rect 36912 42560 36964 42566
rect 36912 42502 36964 42508
rect 36924 42294 36952 42502
rect 36176 42288 36228 42294
rect 36176 42230 36228 42236
rect 36912 42288 36964 42294
rect 36912 42230 36964 42236
rect 36084 41812 36136 41818
rect 36084 41754 36136 41760
rect 36084 41608 36136 41614
rect 36188 41562 36216 42230
rect 36452 42016 36504 42022
rect 36452 41958 36504 41964
rect 36544 42016 36596 42022
rect 36544 41958 36596 41964
rect 36728 42016 36780 42022
rect 36728 41958 36780 41964
rect 36464 41614 36492 41958
rect 36556 41614 36584 41958
rect 36136 41556 36216 41562
rect 36084 41550 36216 41556
rect 36452 41608 36504 41614
rect 36452 41550 36504 41556
rect 36544 41608 36596 41614
rect 36544 41550 36596 41556
rect 35900 41540 35952 41546
rect 36096 41534 36216 41550
rect 35900 41482 35952 41488
rect 35716 41268 35768 41274
rect 35716 41210 35768 41216
rect 35532 40724 35584 40730
rect 35532 40666 35584 40672
rect 35308 40412 35480 40440
rect 35256 40394 35308 40400
rect 35532 40384 35584 40390
rect 35532 40326 35584 40332
rect 34756 39788 34836 39794
rect 34704 39782 34836 39788
rect 34716 39766 34836 39782
rect 34612 39432 34664 39438
rect 34612 39374 34664 39380
rect 33876 39296 33928 39302
rect 32876 39222 33180 39250
rect 33876 39238 33928 39244
rect 32876 39030 32904 39222
rect 32956 39092 33008 39098
rect 32956 39034 33008 39040
rect 32864 39024 32916 39030
rect 32864 38966 32916 38972
rect 32772 38888 32824 38894
rect 32772 38830 32824 38836
rect 32496 38820 32548 38826
rect 32496 38762 32548 38768
rect 32404 38548 32456 38554
rect 32404 38490 32456 38496
rect 32876 37806 32904 38966
rect 32968 37942 32996 39034
rect 33152 39012 33180 39222
rect 33232 39024 33284 39030
rect 33152 38984 33232 39012
rect 33232 38966 33284 38972
rect 33888 38962 33916 39238
rect 33876 38956 33928 38962
rect 33876 38898 33928 38904
rect 34152 38956 34204 38962
rect 34152 38898 34204 38904
rect 33140 38888 33192 38894
rect 33140 38830 33192 38836
rect 33152 38486 33180 38830
rect 33600 38820 33652 38826
rect 33600 38762 33652 38768
rect 33232 38752 33284 38758
rect 33232 38694 33284 38700
rect 33244 38554 33272 38694
rect 33612 38554 33640 38762
rect 33232 38548 33284 38554
rect 33232 38490 33284 38496
rect 33600 38548 33652 38554
rect 33600 38490 33652 38496
rect 33140 38480 33192 38486
rect 33140 38422 33192 38428
rect 33152 38010 33180 38422
rect 33508 38412 33560 38418
rect 33508 38354 33560 38360
rect 33232 38344 33284 38350
rect 33232 38286 33284 38292
rect 33416 38344 33468 38350
rect 33416 38286 33468 38292
rect 33244 38214 33272 38286
rect 33232 38208 33284 38214
rect 33232 38150 33284 38156
rect 33140 38004 33192 38010
rect 33140 37946 33192 37952
rect 32956 37936 33008 37942
rect 32956 37878 33008 37884
rect 32864 37800 32916 37806
rect 32864 37742 32916 37748
rect 32772 37324 32824 37330
rect 32772 37266 32824 37272
rect 32680 36712 32732 36718
rect 32680 36654 32732 36660
rect 32692 36378 32720 36654
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32680 36372 32732 36378
rect 32680 36314 32732 36320
rect 32312 35692 32364 35698
rect 32312 35634 32364 35640
rect 31852 35488 31904 35494
rect 31852 35430 31904 35436
rect 31944 35488 31996 35494
rect 31944 35430 31996 35436
rect 31864 35170 31892 35430
rect 31956 35290 31984 35430
rect 31944 35284 31996 35290
rect 31944 35226 31996 35232
rect 31864 35142 32076 35170
rect 32048 35086 32076 35142
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 32416 35018 32444 36314
rect 32496 36032 32548 36038
rect 32496 35974 32548 35980
rect 32404 35012 32456 35018
rect 32404 34954 32456 34960
rect 32312 34536 32364 34542
rect 32312 34478 32364 34484
rect 32324 33998 32352 34478
rect 32508 33998 32536 35974
rect 32588 35760 32640 35766
rect 32588 35702 32640 35708
rect 32600 33998 32628 35702
rect 32312 33992 32364 33998
rect 32312 33934 32364 33940
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 32588 33992 32640 33998
rect 32588 33934 32640 33940
rect 32036 33856 32088 33862
rect 32036 33798 32088 33804
rect 32128 33856 32180 33862
rect 32128 33798 32180 33804
rect 32048 33658 32076 33798
rect 32036 33652 32088 33658
rect 32036 33594 32088 33600
rect 32140 33590 32168 33798
rect 32324 33658 32352 33934
rect 32312 33652 32364 33658
rect 32312 33594 32364 33600
rect 32508 33590 32536 33934
rect 32128 33584 32180 33590
rect 32128 33526 32180 33532
rect 32496 33584 32548 33590
rect 32496 33526 32548 33532
rect 31576 33448 31628 33454
rect 31576 33390 31628 33396
rect 31588 32298 31616 33390
rect 32140 32366 32168 33526
rect 32600 33318 32628 33934
rect 32784 33930 32812 37266
rect 32876 34202 32904 37742
rect 32956 37664 33008 37670
rect 32956 37606 33008 37612
rect 32968 36650 32996 37606
rect 33140 36916 33192 36922
rect 33140 36858 33192 36864
rect 32956 36644 33008 36650
rect 32956 36586 33008 36592
rect 33152 36378 33180 36858
rect 33244 36718 33272 38150
rect 33428 37874 33456 38286
rect 33520 37874 33548 38354
rect 33876 38276 33928 38282
rect 33876 38218 33928 38224
rect 33416 37868 33468 37874
rect 33416 37810 33468 37816
rect 33508 37868 33560 37874
rect 33508 37810 33560 37816
rect 33324 37120 33376 37126
rect 33324 37062 33376 37068
rect 33232 36712 33284 36718
rect 33232 36654 33284 36660
rect 33244 36582 33272 36654
rect 33336 36650 33364 37062
rect 33428 36786 33456 37810
rect 33520 37262 33548 37810
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33888 37194 33916 38218
rect 33876 37188 33928 37194
rect 33876 37130 33928 37136
rect 34060 37188 34112 37194
rect 34060 37130 34112 37136
rect 33888 36922 33916 37130
rect 34072 36922 34100 37130
rect 33876 36916 33928 36922
rect 33876 36858 33928 36864
rect 34060 36916 34112 36922
rect 34060 36858 34112 36864
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 33876 36780 33928 36786
rect 33876 36722 33928 36728
rect 33968 36780 34020 36786
rect 33968 36722 34020 36728
rect 33324 36644 33376 36650
rect 33324 36586 33376 36592
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 33152 35494 33180 35974
rect 33244 35766 33272 36518
rect 33336 36310 33364 36586
rect 33324 36304 33376 36310
rect 33324 36246 33376 36252
rect 33888 36242 33916 36722
rect 33980 36378 34008 36722
rect 33968 36372 34020 36378
rect 33968 36314 34020 36320
rect 33876 36236 33928 36242
rect 33876 36178 33928 36184
rect 33324 36168 33376 36174
rect 33324 36110 33376 36116
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33336 35766 33364 36110
rect 33232 35760 33284 35766
rect 33232 35702 33284 35708
rect 33324 35760 33376 35766
rect 33324 35702 33376 35708
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 33336 34202 33364 35702
rect 33520 35698 33548 36110
rect 33600 36100 33652 36106
rect 33600 36042 33652 36048
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 33520 34746 33548 35634
rect 33612 35630 33640 36042
rect 33600 35624 33652 35630
rect 33600 35566 33652 35572
rect 33508 34740 33560 34746
rect 33508 34682 33560 34688
rect 32864 34196 32916 34202
rect 32864 34138 32916 34144
rect 33324 34196 33376 34202
rect 33324 34138 33376 34144
rect 32772 33924 32824 33930
rect 32772 33866 32824 33872
rect 32784 33522 32812 33866
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32588 33312 32640 33318
rect 32588 33254 32640 33260
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 31576 32292 31628 32298
rect 31576 32234 31628 32240
rect 32140 32026 32168 32302
rect 32128 32020 32180 32026
rect 32128 31962 32180 31968
rect 31760 31952 31812 31958
rect 31760 31894 31812 31900
rect 31576 31816 31628 31822
rect 31576 31758 31628 31764
rect 31588 31414 31616 31758
rect 31772 31754 31800 31894
rect 31944 31884 31996 31890
rect 31944 31826 31996 31832
rect 31760 31748 31812 31754
rect 31760 31690 31812 31696
rect 31576 31408 31628 31414
rect 31576 31350 31628 31356
rect 31956 31210 31984 31826
rect 32876 31754 32904 34138
rect 33520 34066 33548 34682
rect 33784 34196 33836 34202
rect 33784 34138 33836 34144
rect 33508 34060 33560 34066
rect 33508 34002 33560 34008
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 33060 33522 33088 33798
rect 33244 33522 33272 33798
rect 33416 33652 33468 33658
rect 33416 33594 33468 33600
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33048 33312 33100 33318
rect 33048 33254 33100 33260
rect 32600 31726 32904 31754
rect 31944 31204 31996 31210
rect 31944 31146 31996 31152
rect 32036 30932 32088 30938
rect 32036 30874 32088 30880
rect 32048 30666 32076 30874
rect 31852 30660 31904 30666
rect 31852 30602 31904 30608
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 31864 30394 31892 30602
rect 31852 30388 31904 30394
rect 31852 30330 31904 30336
rect 32600 30258 32628 31726
rect 32864 31476 32916 31482
rect 32864 31418 32916 31424
rect 32680 31204 32732 31210
rect 32680 31146 32732 31152
rect 32692 30394 32720 31146
rect 32876 31142 32904 31418
rect 32772 31136 32824 31142
rect 32772 31078 32824 31084
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32784 30394 32812 31078
rect 32680 30388 32732 30394
rect 32680 30330 32732 30336
rect 32772 30388 32824 30394
rect 32772 30330 32824 30336
rect 32588 30252 32640 30258
rect 32588 30194 32640 30200
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31588 28694 31616 29106
rect 32128 29028 32180 29034
rect 32128 28970 32180 28976
rect 31944 28960 31996 28966
rect 31944 28902 31996 28908
rect 31576 28688 31628 28694
rect 31576 28630 31628 28636
rect 31588 28200 31616 28630
rect 31760 28484 31812 28490
rect 31760 28426 31812 28432
rect 31668 28212 31720 28218
rect 31588 28172 31668 28200
rect 31668 28154 31720 28160
rect 31772 27878 31800 28426
rect 31956 28082 31984 28902
rect 32140 28694 32168 28970
rect 32600 28762 32628 30194
rect 32864 30048 32916 30054
rect 32864 29990 32916 29996
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32128 28688 32180 28694
rect 32128 28630 32180 28636
rect 32312 28552 32364 28558
rect 32312 28494 32364 28500
rect 32036 28416 32088 28422
rect 32036 28358 32088 28364
rect 32048 28082 32076 28358
rect 32324 28257 32352 28494
rect 32680 28416 32732 28422
rect 32680 28358 32732 28364
rect 32310 28248 32366 28257
rect 32310 28183 32312 28192
rect 32364 28183 32366 28192
rect 32312 28154 32364 28160
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 32036 28076 32088 28082
rect 32036 28018 32088 28024
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 31944 27328 31996 27334
rect 31944 27270 31996 27276
rect 31956 26858 31984 27270
rect 32048 27130 32076 28018
rect 32324 27130 32352 28018
rect 32692 27470 32720 28358
rect 32680 27464 32732 27470
rect 32680 27406 32732 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32404 27328 32456 27334
rect 32404 27270 32456 27276
rect 32036 27124 32088 27130
rect 32036 27066 32088 27072
rect 32312 27124 32364 27130
rect 32312 27066 32364 27072
rect 31944 26852 31996 26858
rect 31944 26794 31996 26800
rect 31956 26042 31984 26794
rect 32128 26512 32180 26518
rect 32128 26454 32180 26460
rect 32036 26240 32088 26246
rect 32036 26182 32088 26188
rect 31944 26036 31996 26042
rect 31944 25978 31996 25984
rect 32048 25974 32076 26182
rect 32036 25968 32088 25974
rect 32036 25910 32088 25916
rect 32140 25906 32168 26454
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 31588 24818 31616 25842
rect 32416 25838 32444 27270
rect 32600 26314 32628 27338
rect 32876 27334 32904 29990
rect 33060 28994 33088 33254
rect 33336 32570 33364 33458
rect 33428 32774 33456 33594
rect 33520 32994 33548 34002
rect 33692 33992 33744 33998
rect 33692 33934 33744 33940
rect 33704 33658 33732 33934
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 33796 33522 33824 34138
rect 33784 33516 33836 33522
rect 33784 33458 33836 33464
rect 33888 33386 33916 36178
rect 34164 36106 34192 38898
rect 34808 38350 34836 39766
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35544 39438 35572 40326
rect 35728 40202 35756 41210
rect 35912 40526 35940 41482
rect 36188 41070 36216 41534
rect 36268 41472 36320 41478
rect 36268 41414 36320 41420
rect 36280 41274 36308 41414
rect 36268 41268 36320 41274
rect 36268 41210 36320 41216
rect 36176 41064 36228 41070
rect 36176 41006 36228 41012
rect 36084 40928 36136 40934
rect 36084 40870 36136 40876
rect 35900 40520 35952 40526
rect 35900 40462 35952 40468
rect 35992 40452 36044 40458
rect 35992 40394 36044 40400
rect 35728 40174 35940 40202
rect 36004 40186 36032 40394
rect 35532 39432 35584 39438
rect 35532 39374 35584 39380
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 34808 37330 34836 38286
rect 35256 38276 35308 38282
rect 35256 38218 35308 38224
rect 35268 37806 35296 38218
rect 35544 38010 35572 39374
rect 35912 39030 35940 40174
rect 35992 40180 36044 40186
rect 35992 40122 36044 40128
rect 36096 40118 36124 40870
rect 36188 40458 36216 41006
rect 36740 40730 36768 41958
rect 36728 40724 36780 40730
rect 36728 40666 36780 40672
rect 36924 40526 36952 42230
rect 36912 40520 36964 40526
rect 36912 40462 36964 40468
rect 36176 40452 36228 40458
rect 36176 40394 36228 40400
rect 36084 40112 36136 40118
rect 36084 40054 36136 40060
rect 35900 39024 35952 39030
rect 35900 38966 35952 38972
rect 36728 38888 36780 38894
rect 36728 38830 36780 38836
rect 35900 38752 35952 38758
rect 35900 38694 35952 38700
rect 35532 38004 35584 38010
rect 35532 37946 35584 37952
rect 35912 37806 35940 38694
rect 36740 38214 36768 38830
rect 36912 38820 36964 38826
rect 36912 38762 36964 38768
rect 36924 38350 36952 38762
rect 36912 38344 36964 38350
rect 36912 38286 36964 38292
rect 36728 38208 36780 38214
rect 36728 38150 36780 38156
rect 36740 37942 36768 38150
rect 36728 37936 36780 37942
rect 36728 37878 36780 37884
rect 36820 37868 36872 37874
rect 36820 37810 36872 37816
rect 35256 37800 35308 37806
rect 35256 37742 35308 37748
rect 35900 37800 35952 37806
rect 35900 37742 35952 37748
rect 35808 37664 35860 37670
rect 35808 37606 35860 37612
rect 35992 37664 36044 37670
rect 35992 37606 36044 37612
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 35348 37188 35400 37194
rect 35348 37130 35400 37136
rect 35360 36922 35388 37130
rect 35348 36916 35400 36922
rect 35348 36858 35400 36864
rect 35820 36854 35848 37606
rect 36004 37330 36032 37606
rect 36832 37466 36860 37810
rect 36820 37460 36872 37466
rect 36820 37402 36872 37408
rect 35992 37324 36044 37330
rect 35992 37266 36044 37272
rect 35808 36848 35860 36854
rect 35808 36790 35860 36796
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 34256 36378 34284 36722
rect 36004 36582 36032 37266
rect 36924 37262 36952 38286
rect 36912 37256 36964 37262
rect 36912 37198 36964 37204
rect 35992 36576 36044 36582
rect 35992 36518 36044 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34244 36372 34296 36378
rect 34244 36314 34296 36320
rect 36924 36174 36952 37198
rect 36912 36168 36964 36174
rect 36912 36110 36964 36116
rect 34152 36100 34204 36106
rect 34152 36042 34204 36048
rect 36924 35766 36952 36110
rect 36912 35760 36964 35766
rect 36912 35702 36964 35708
rect 36084 35624 36136 35630
rect 36084 35566 36136 35572
rect 36360 35624 36412 35630
rect 36360 35566 36412 35572
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 34440 35154 34468 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34428 35148 34480 35154
rect 34428 35090 34480 35096
rect 35808 35080 35860 35086
rect 35808 35022 35860 35028
rect 35348 34944 35400 34950
rect 35348 34886 35400 34892
rect 35360 34678 35388 34886
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 35348 34672 35400 34678
rect 35348 34614 35400 34620
rect 34060 34196 34112 34202
rect 34060 34138 34112 34144
rect 33876 33380 33928 33386
rect 33876 33322 33928 33328
rect 33876 33040 33928 33046
rect 33520 32966 33640 32994
rect 33876 32982 33928 32988
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33416 32768 33468 32774
rect 33416 32710 33468 32716
rect 33324 32564 33376 32570
rect 33324 32506 33376 32512
rect 33232 31748 33284 31754
rect 33232 31690 33284 31696
rect 33244 31346 33272 31690
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 33232 30660 33284 30666
rect 33232 30602 33284 30608
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33152 30394 33180 30534
rect 33140 30388 33192 30394
rect 33140 30330 33192 30336
rect 33244 30274 33272 30602
rect 33324 30388 33376 30394
rect 33428 30376 33456 32710
rect 33520 31278 33548 32846
rect 33612 32502 33640 32966
rect 33600 32496 33652 32502
rect 33600 32438 33652 32444
rect 33784 32292 33836 32298
rect 33784 32234 33836 32240
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33376 30348 33456 30376
rect 33324 30330 33376 30336
rect 33152 30258 33272 30274
rect 33140 30252 33272 30258
rect 33192 30246 33272 30252
rect 33140 30194 33192 30200
rect 33520 30054 33548 31214
rect 33692 30796 33744 30802
rect 33692 30738 33744 30744
rect 33704 30258 33732 30738
rect 33692 30252 33744 30258
rect 33692 30194 33744 30200
rect 33508 30048 33560 30054
rect 33508 29990 33560 29996
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33428 29170 33456 29446
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33060 28966 33180 28994
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 32968 28218 32996 28562
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32312 25764 32364 25770
rect 32312 25706 32364 25712
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 31944 25152 31996 25158
rect 31944 25094 31996 25100
rect 31956 24886 31984 25094
rect 32140 24954 32168 25230
rect 32128 24948 32180 24954
rect 32128 24890 32180 24896
rect 31944 24880 31996 24886
rect 31944 24822 31996 24828
rect 32324 24818 32352 25706
rect 32600 24886 32628 26250
rect 32772 26240 32824 26246
rect 32772 26182 32824 26188
rect 32784 25906 32812 26182
rect 32876 25974 32904 26930
rect 32864 25968 32916 25974
rect 32864 25910 32916 25916
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32588 24880 32640 24886
rect 32588 24822 32640 24828
rect 31576 24812 31628 24818
rect 31576 24754 31628 24760
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 31588 22030 31616 24754
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31680 22778 31708 23122
rect 31668 22772 31720 22778
rect 31668 22714 31720 22720
rect 31760 22568 31812 22574
rect 31760 22510 31812 22516
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31772 21962 31800 22510
rect 31760 21956 31812 21962
rect 31760 21898 31812 21904
rect 32048 21894 32076 24754
rect 32692 24274 32720 25774
rect 32680 24268 32732 24274
rect 32680 24210 32732 24216
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 33060 23866 33088 24074
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 32496 23588 32548 23594
rect 32496 23530 32548 23536
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32232 22438 32260 22578
rect 32416 22506 32444 22578
rect 32404 22500 32456 22506
rect 32404 22442 32456 22448
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32232 22098 32260 22374
rect 32220 22092 32272 22098
rect 32220 22034 32272 22040
rect 32220 21956 32272 21962
rect 32220 21898 32272 21904
rect 32312 21956 32364 21962
rect 32312 21898 32364 21904
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31576 19916 31628 19922
rect 31576 19858 31628 19864
rect 31588 19378 31616 19858
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31772 19378 31800 19790
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31680 18222 31708 19314
rect 31864 19242 31892 20878
rect 31852 19236 31904 19242
rect 31852 19178 31904 19184
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31576 17740 31628 17746
rect 31576 17682 31628 17688
rect 31588 17270 31616 17682
rect 31956 17678 31984 21490
rect 32048 19514 32076 21830
rect 32232 20942 32260 21898
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32324 19922 32352 21898
rect 32312 19916 32364 19922
rect 32312 19858 32364 19864
rect 32036 19508 32088 19514
rect 32036 19450 32088 19456
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 32220 17672 32272 17678
rect 32220 17614 32272 17620
rect 32312 17672 32364 17678
rect 32312 17614 32364 17620
rect 31576 17264 31628 17270
rect 31576 17206 31628 17212
rect 32232 17202 32260 17614
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32128 17060 32180 17066
rect 32128 17002 32180 17008
rect 32140 16658 32168 17002
rect 32128 16652 32180 16658
rect 32128 16594 32180 16600
rect 32232 16590 32260 17138
rect 32324 17134 32352 17614
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32416 17202 32444 17478
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 31852 16584 31904 16590
rect 31496 16510 31800 16538
rect 31852 16526 31904 16532
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31496 16114 31524 16390
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31576 16040 31628 16046
rect 31404 15988 31576 15994
rect 31772 15994 31800 16510
rect 31864 16250 31892 16526
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 32218 16144 32274 16153
rect 32218 16079 32220 16088
rect 32272 16079 32274 16088
rect 32220 16050 32272 16056
rect 31404 15982 31628 15988
rect 31404 15966 31616 15982
rect 31680 15966 31800 15994
rect 31850 16008 31906 16017
rect 31298 15943 31354 15952
rect 31300 15700 31352 15706
rect 31300 15642 31352 15648
rect 31312 14414 31340 15642
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31300 14408 31352 14414
rect 31352 14356 31432 14362
rect 31300 14350 31432 14356
rect 31312 14334 31432 14350
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 31116 14000 31168 14006
rect 31116 13942 31168 13948
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30656 13864 30708 13870
rect 30656 13806 30708 13812
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 30472 13796 30524 13802
rect 30472 13738 30524 13744
rect 30668 13410 30696 13806
rect 30760 13530 30788 13806
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30748 13524 30800 13530
rect 30748 13466 30800 13472
rect 30668 13382 30788 13410
rect 30380 13320 30432 13326
rect 30300 13268 30380 13274
rect 30300 13262 30432 13268
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 29184 13184 29236 13190
rect 26974 13152 27030 13161
rect 29184 13126 29236 13132
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 26974 13087 27030 13096
rect 26988 12986 27016 13087
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 29196 12850 29224 13126
rect 29564 12986 29592 13126
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26528 12442 26556 12582
rect 26620 12442 26648 12786
rect 27160 12640 27212 12646
rect 27528 12640 27580 12646
rect 27160 12582 27212 12588
rect 27264 12600 27528 12628
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26608 12436 26660 12442
rect 27172 12434 27200 12582
rect 26608 12378 26660 12384
rect 26988 12406 27200 12434
rect 26988 12306 27016 12406
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 27068 12300 27120 12306
rect 27068 12242 27120 12248
rect 27080 12186 27108 12242
rect 27264 12186 27292 12600
rect 27528 12582 27580 12588
rect 27632 12442 27660 12786
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27632 12306 27660 12378
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27080 12158 27292 12186
rect 27632 12170 27660 12242
rect 27264 11354 27292 12158
rect 27436 12164 27488 12170
rect 27436 12106 27488 12112
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27448 11694 27476 12106
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27528 11688 27580 11694
rect 27632 11676 27660 12106
rect 28828 11830 28856 12786
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 28816 11824 28868 11830
rect 28816 11766 28868 11772
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27580 11648 27660 11676
rect 27528 11630 27580 11636
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 26976 9920 27028 9926
rect 26976 9862 27028 9868
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26620 9042 26648 9454
rect 26988 9042 27016 9862
rect 27264 9042 27292 10542
rect 27356 9722 27384 10610
rect 27436 10600 27488 10606
rect 27540 10588 27568 11630
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27632 11121 27660 11222
rect 27618 11112 27674 11121
rect 27618 11047 27674 11056
rect 27724 10674 27752 11698
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27488 10560 27568 10588
rect 27436 10542 27488 10548
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27356 9450 27384 9658
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 26620 8430 26648 8978
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26896 8634 26924 8774
rect 26884 8628 26936 8634
rect 26884 8570 26936 8576
rect 26608 8424 26660 8430
rect 26608 8366 26660 8372
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7410 26556 7890
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26516 6316 26568 6322
rect 26620 6304 26648 8366
rect 26988 7546 27016 8978
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 26712 7002 26740 7482
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 26804 7313 26832 7346
rect 26790 7304 26846 7313
rect 26790 7239 26846 7248
rect 27080 7206 27108 8366
rect 27160 8356 27212 8362
rect 27160 8298 27212 8304
rect 27172 7478 27200 8298
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 27068 7200 27120 7206
rect 27068 7142 27120 7148
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 26712 6866 26740 6938
rect 27172 6866 27200 7414
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 26568 6276 26648 6304
rect 27080 6746 27108 6802
rect 27264 6746 27292 8978
rect 27448 7954 27476 10542
rect 27724 8974 27752 10610
rect 27816 10266 27844 10746
rect 27804 10260 27856 10266
rect 27804 10202 27856 10208
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 27724 8090 27752 8910
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 27448 7342 27476 7890
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27080 6718 27292 6746
rect 26516 6258 26568 6264
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26528 5302 26556 6258
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26056 5092 26108 5098
rect 26056 5034 26108 5040
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 25412 4548 25464 4554
rect 25412 4490 25464 4496
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24490 4176 24546 4185
rect 24584 4140 24636 4146
rect 24546 4120 24584 4128
rect 24490 4111 24584 4120
rect 24504 4100 24584 4111
rect 24584 4082 24636 4088
rect 25424 4010 25452 4490
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 24504 3738 24532 3946
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24872 3738 24900 3878
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23400 3074 23428 3182
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 22928 3052 22980 3058
rect 23400 3046 23520 3074
rect 24412 3058 24440 3538
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 22928 2994 22980 3000
rect 23492 2990 23520 3046
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 24872 2854 24900 3130
rect 25424 3126 25452 3946
rect 26068 3942 26096 5034
rect 26252 4622 26280 5170
rect 27080 5030 27108 6718
rect 27448 6390 27476 7278
rect 27540 6866 27568 7686
rect 27724 7410 27752 7686
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27724 7002 27752 7346
rect 27712 6996 27764 7002
rect 27712 6938 27764 6944
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27816 6798 27844 9114
rect 27908 8974 27936 11086
rect 28644 10674 28672 11086
rect 29012 10742 29040 12582
rect 29748 12306 29776 13262
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28264 10464 28316 10470
rect 28264 10406 28316 10412
rect 28276 10266 28304 10406
rect 28264 10260 28316 10266
rect 28264 10202 28316 10208
rect 28552 10130 28580 10542
rect 28644 10266 28672 10610
rect 28632 10260 28684 10266
rect 28632 10202 28684 10208
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29288 10130 29316 10202
rect 28540 10124 28592 10130
rect 28540 10066 28592 10072
rect 29276 10124 29328 10130
rect 29276 10066 29328 10072
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28632 10056 28684 10062
rect 28632 9998 28684 10004
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28460 9382 28488 9998
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27908 7546 27936 8910
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28184 8430 28212 8842
rect 28552 8634 28580 9454
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28644 8566 28672 9998
rect 28920 9722 28948 9998
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28920 9586 28948 9658
rect 29288 9586 29316 10066
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28632 8560 28684 8566
rect 28632 8502 28684 8508
rect 28172 8424 28224 8430
rect 28172 8366 28224 8372
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28276 7546 28304 8026
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 27908 6798 27936 7482
rect 28460 6798 28488 7754
rect 28644 7750 28672 8502
rect 28828 8362 28856 9318
rect 29288 8974 29316 9522
rect 29276 8968 29328 8974
rect 29276 8910 29328 8916
rect 29184 8900 29236 8906
rect 29184 8842 29236 8848
rect 29196 8430 29224 8842
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 28828 8090 28856 8298
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 29196 7954 29224 8366
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 28632 7744 28684 7750
rect 28632 7686 28684 7692
rect 28920 7546 28948 7890
rect 29276 7880 29328 7886
rect 29276 7822 29328 7828
rect 29288 7546 29316 7822
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 28724 7472 28776 7478
rect 28722 7440 28724 7449
rect 28776 7440 28778 7449
rect 28722 7375 28778 7384
rect 28920 6882 28948 7482
rect 29012 7274 29224 7290
rect 29000 7268 29236 7274
rect 29052 7262 29184 7268
rect 29000 7210 29052 7216
rect 29184 7210 29236 7216
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 28828 6866 28948 6882
rect 28816 6860 28948 6866
rect 28868 6854 28948 6860
rect 28816 6802 28868 6808
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 27816 6458 27844 6734
rect 28828 6458 28856 6802
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 28920 6322 28948 6734
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 29012 6186 29040 6734
rect 29104 6322 29132 7142
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29000 6180 29052 6186
rect 29000 6122 29052 6128
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28368 4690 28396 4966
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 26068 3126 26096 3878
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 24872 2446 24900 2790
rect 26712 2650 26740 3470
rect 27540 3466 27568 3946
rect 27632 3942 27660 4558
rect 28920 4146 28948 4694
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3602 27660 3878
rect 29012 3738 29040 5102
rect 29380 4826 29408 12174
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 29564 11354 29592 11494
rect 29932 11354 29960 12786
rect 30116 12238 30144 13262
rect 30300 13246 30420 13262
rect 30300 12850 30328 13246
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29472 10742 29500 11018
rect 29748 10810 29776 11086
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29564 9586 29592 10678
rect 29840 10266 29868 11086
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29736 10192 29788 10198
rect 29736 10134 29788 10140
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29564 8498 29592 9522
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29656 8838 29684 9318
rect 29748 9042 29776 10134
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29460 7472 29512 7478
rect 29458 7440 29460 7449
rect 29512 7440 29514 7449
rect 29656 7410 29684 8774
rect 29748 8634 29776 8978
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29840 7886 29868 10202
rect 30024 9518 30052 10542
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30116 7886 30144 11018
rect 30300 10810 30328 12174
rect 30484 10810 30512 13126
rect 30576 12442 30604 13262
rect 30668 12986 30696 13262
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30760 11762 30788 13382
rect 30944 13190 30972 13738
rect 31036 13530 31064 13806
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30932 13184 30984 13190
rect 30932 13126 30984 13132
rect 31128 12238 31156 13942
rect 31208 13524 31260 13530
rect 31208 13466 31260 13472
rect 31220 12850 31248 13466
rect 31312 12986 31340 14214
rect 31404 13734 31432 14334
rect 31496 13870 31524 14758
rect 31680 14414 31708 15966
rect 31850 15943 31852 15952
rect 31904 15943 31906 15952
rect 31852 15914 31904 15920
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 31392 13728 31444 13734
rect 31392 13670 31444 13676
rect 31404 13326 31432 13670
rect 31496 13530 31524 13806
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 31392 13320 31444 13326
rect 31392 13262 31444 13268
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31496 12889 31524 13262
rect 31588 12986 31616 13942
rect 31680 13938 31708 14350
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31680 13326 31708 13874
rect 32508 13394 32536 23530
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32600 22778 32628 22918
rect 32968 22778 32996 22918
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 33152 22080 33180 28966
rect 33520 28490 33548 29990
rect 33692 29572 33744 29578
rect 33692 29514 33744 29520
rect 33704 29170 33732 29514
rect 33692 29164 33744 29170
rect 33692 29106 33744 29112
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33612 27674 33640 27950
rect 33600 27668 33652 27674
rect 33600 27610 33652 27616
rect 33796 27470 33824 32234
rect 33888 28642 33916 32982
rect 34072 32910 34100 34138
rect 34428 33856 34480 33862
rect 34428 33798 34480 33804
rect 34440 33658 34468 33798
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 34520 33652 34572 33658
rect 34520 33594 34572 33600
rect 34532 32978 34560 33594
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 34060 32904 34112 32910
rect 34060 32846 34112 32852
rect 34072 32026 34100 32846
rect 34520 32768 34572 32774
rect 34520 32710 34572 32716
rect 34532 32502 34560 32710
rect 34520 32496 34572 32502
rect 34520 32438 34572 32444
rect 34624 32450 34652 34614
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 35348 34536 35400 34542
rect 35348 34478 35400 34484
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34202 35388 34478
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 34796 34060 34848 34066
rect 34796 34002 34848 34008
rect 34704 33380 34756 33386
rect 34704 33322 34756 33328
rect 34716 33114 34744 33322
rect 34808 33114 34836 34002
rect 35452 33522 35480 34546
rect 35820 34542 35848 35022
rect 36096 34746 36124 35566
rect 36372 35290 36400 35566
rect 36360 35284 36412 35290
rect 36360 35226 36412 35232
rect 36924 35018 36952 35702
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 36912 35012 36964 35018
rect 36912 34954 36964 34960
rect 36084 34740 36136 34746
rect 36084 34682 36136 34688
rect 36188 34678 36216 34954
rect 36544 34944 36596 34950
rect 36544 34886 36596 34892
rect 36556 34678 36584 34886
rect 36176 34672 36228 34678
rect 36176 34614 36228 34620
rect 36544 34672 36596 34678
rect 36544 34614 36596 34620
rect 35808 34536 35860 34542
rect 35808 34478 35860 34484
rect 36268 34536 36320 34542
rect 36268 34478 36320 34484
rect 36544 34536 36596 34542
rect 36544 34478 36596 34484
rect 36280 34406 36308 34478
rect 36268 34400 36320 34406
rect 36268 34342 36320 34348
rect 35348 33516 35400 33522
rect 35348 33458 35400 33464
rect 35440 33516 35492 33522
rect 35440 33458 35492 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 33114 35388 33458
rect 34704 33108 34756 33114
rect 34704 33050 34756 33056
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 35348 33108 35400 33114
rect 35348 33050 35400 33056
rect 35256 32904 35308 32910
rect 35256 32846 35308 32852
rect 35268 32570 35296 32846
rect 35256 32564 35308 32570
rect 35256 32506 35308 32512
rect 34624 32434 34744 32450
rect 34624 32428 34756 32434
rect 34624 32422 34704 32428
rect 34704 32370 34756 32376
rect 34060 32020 34112 32026
rect 34060 31962 34112 31968
rect 34336 31748 34388 31754
rect 34336 31690 34388 31696
rect 34428 31748 34480 31754
rect 34428 31690 34480 31696
rect 34244 30796 34296 30802
rect 34244 30738 34296 30744
rect 34152 30728 34204 30734
rect 34152 30670 34204 30676
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 34072 29850 34100 30194
rect 34164 30190 34192 30670
rect 34256 30258 34284 30738
rect 34244 30252 34296 30258
rect 34348 30240 34376 31690
rect 34440 30938 34468 31690
rect 34428 30932 34480 30938
rect 34428 30874 34480 30880
rect 34428 30252 34480 30258
rect 34348 30212 34428 30240
rect 34244 30194 34296 30200
rect 34428 30194 34480 30200
rect 34152 30184 34204 30190
rect 34152 30126 34204 30132
rect 34060 29844 34112 29850
rect 34060 29786 34112 29792
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33980 29306 34008 29582
rect 34440 29510 34468 30194
rect 34716 29646 34744 32370
rect 36176 32360 36228 32366
rect 36176 32302 36228 32308
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 31482 35388 32166
rect 36188 31754 36216 32302
rect 36004 31726 36216 31754
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 35808 31476 35860 31482
rect 35808 31418 35860 31424
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30796 34848 30802
rect 34796 30738 34848 30744
rect 34808 30394 34836 30738
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 35256 30592 35308 30598
rect 35256 30534 35308 30540
rect 35268 30394 35296 30534
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 35256 30388 35308 30394
rect 35256 30330 35308 30336
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34428 29504 34480 29510
rect 34428 29446 34480 29452
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 34716 29238 34744 29582
rect 34612 29232 34664 29238
rect 34612 29174 34664 29180
rect 34704 29232 34756 29238
rect 34704 29174 34756 29180
rect 33968 29028 34020 29034
rect 33968 28970 34020 28976
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 33980 28762 34008 28970
rect 33968 28756 34020 28762
rect 33968 28698 34020 28704
rect 33888 28614 34008 28642
rect 33876 28144 33928 28150
rect 33876 28086 33928 28092
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 33244 25770 33272 27406
rect 33888 27334 33916 28086
rect 33876 27328 33928 27334
rect 33876 27270 33928 27276
rect 33888 26450 33916 27270
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33980 26382 34008 28614
rect 34532 28529 34560 28970
rect 34518 28520 34574 28529
rect 34518 28455 34574 28464
rect 34336 28416 34388 28422
rect 34336 28358 34388 28364
rect 34348 28014 34376 28358
rect 34336 28008 34388 28014
rect 34336 27950 34388 27956
rect 34348 27538 34376 27950
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34532 27130 34560 28455
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34624 26994 34652 29174
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28558 35388 30670
rect 35716 30660 35768 30666
rect 35716 30602 35768 30608
rect 35728 30394 35756 30602
rect 35716 30388 35768 30394
rect 35716 30330 35768 30336
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 35452 29850 35480 30194
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34072 26314 34100 26794
rect 33600 26308 33652 26314
rect 33600 26250 33652 26256
rect 34060 26308 34112 26314
rect 34060 26250 34112 26256
rect 33612 26042 33640 26250
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33232 25764 33284 25770
rect 33232 25706 33284 25712
rect 34072 23730 34100 26250
rect 34256 26246 34284 26930
rect 34428 26920 34480 26926
rect 34716 26874 34744 27814
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35164 27396 35216 27402
rect 35164 27338 35216 27344
rect 35176 27130 35204 27338
rect 35360 27334 35388 28494
rect 35716 28008 35768 28014
rect 35716 27950 35768 27956
rect 35728 27674 35756 27950
rect 35716 27668 35768 27674
rect 35716 27610 35768 27616
rect 35820 27538 35848 31418
rect 36004 30938 36032 31726
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 36004 30258 36032 30874
rect 36280 30818 36308 34342
rect 36556 33658 36584 34478
rect 36912 33856 36964 33862
rect 36912 33798 36964 33804
rect 36924 33658 36952 33798
rect 36544 33652 36596 33658
rect 36544 33594 36596 33600
rect 36912 33652 36964 33658
rect 36912 33594 36964 33600
rect 36556 31822 36584 33594
rect 36820 33516 36872 33522
rect 36820 33458 36872 33464
rect 36832 31822 36860 33458
rect 36544 31816 36596 31822
rect 36820 31816 36872 31822
rect 36544 31758 36596 31764
rect 36740 31776 36820 31804
rect 36096 30790 36308 30818
rect 35992 30252 36044 30258
rect 35992 30194 36044 30200
rect 35900 29844 35952 29850
rect 35900 29786 35952 29792
rect 35912 28082 35940 29786
rect 35992 28960 36044 28966
rect 35992 28902 36044 28908
rect 36004 28626 36032 28902
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 35900 28076 35952 28082
rect 35900 28018 35952 28024
rect 35808 27532 35860 27538
rect 35808 27474 35860 27480
rect 35348 27328 35400 27334
rect 35348 27270 35400 27276
rect 35164 27124 35216 27130
rect 35164 27066 35216 27072
rect 34480 26868 34744 26874
rect 34428 26862 34744 26868
rect 34440 26846 34744 26862
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34244 26240 34296 26246
rect 34244 26182 34296 26188
rect 34704 26240 34756 26246
rect 34704 26182 34756 26188
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 34152 23724 34204 23730
rect 34256 23712 34284 26182
rect 34716 26042 34744 26182
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 35360 25906 35388 27270
rect 35912 26858 35940 28018
rect 36004 27946 36032 28426
rect 35992 27940 36044 27946
rect 35992 27882 36044 27888
rect 36004 27334 36032 27882
rect 35992 27328 36044 27334
rect 35992 27270 36044 27276
rect 35900 26852 35952 26858
rect 35900 26794 35952 26800
rect 35440 26376 35492 26382
rect 35440 26318 35492 26324
rect 35452 26042 35480 26318
rect 35900 26240 35952 26246
rect 35900 26182 35952 26188
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 35348 25900 35400 25906
rect 35348 25842 35400 25848
rect 34428 24608 34480 24614
rect 34428 24550 34480 24556
rect 34204 23684 34284 23712
rect 34152 23666 34204 23672
rect 34072 23610 34100 23666
rect 33980 23582 34100 23610
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33888 22642 33916 23054
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33980 22094 34008 23582
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 34072 22778 34100 23054
rect 34060 22772 34112 22778
rect 34060 22714 34112 22720
rect 34164 22681 34192 23666
rect 34244 22976 34296 22982
rect 34244 22918 34296 22924
rect 34256 22778 34284 22918
rect 34244 22772 34296 22778
rect 34244 22714 34296 22720
rect 34150 22672 34206 22681
rect 34206 22630 34284 22658
rect 34150 22607 34206 22616
rect 33152 22052 33272 22080
rect 33980 22066 34100 22094
rect 33244 21622 33272 22052
rect 33232 21616 33284 21622
rect 33232 21558 33284 21564
rect 33784 21616 33836 21622
rect 33784 21558 33836 21564
rect 33232 20868 33284 20874
rect 33508 20868 33560 20874
rect 33284 20828 33508 20856
rect 33232 20810 33284 20816
rect 33508 20810 33560 20816
rect 32956 20800 33008 20806
rect 32956 20742 33008 20748
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 32968 20398 32996 20742
rect 33704 20466 33732 20742
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 32956 20392 33008 20398
rect 32956 20334 33008 20340
rect 33416 20324 33468 20330
rect 33416 20266 33468 20272
rect 33428 20058 33456 20266
rect 33600 20256 33652 20262
rect 33600 20198 33652 20204
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 33612 19854 33640 20198
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33796 19718 33824 21558
rect 33968 21548 34020 21554
rect 33968 21490 34020 21496
rect 33980 21146 34008 21490
rect 34072 21418 34100 22066
rect 34152 22092 34204 22098
rect 34152 22034 34204 22040
rect 34060 21412 34112 21418
rect 34060 21354 34112 21360
rect 34164 21146 34192 22034
rect 34256 22030 34284 22630
rect 34440 22234 34468 24550
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 34532 23118 34560 24210
rect 34808 24138 34836 25842
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24132 34848 24138
rect 34796 24074 34848 24080
rect 34704 24064 34756 24070
rect 34704 24006 34756 24012
rect 34716 23866 34744 24006
rect 35452 23866 35480 25978
rect 35912 25974 35940 26182
rect 36004 26042 36032 27270
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 35900 25968 35952 25974
rect 35900 25910 35952 25916
rect 35716 25832 35768 25838
rect 35716 25774 35768 25780
rect 35728 25362 35756 25774
rect 35716 25356 35768 25362
rect 35716 25298 35768 25304
rect 35728 24818 35756 25298
rect 36004 25294 36032 25978
rect 35992 25288 36044 25294
rect 35992 25230 36044 25236
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 35808 24064 35860 24070
rect 35808 24006 35860 24012
rect 34704 23860 34756 23866
rect 34704 23802 34756 23808
rect 35440 23860 35492 23866
rect 35440 23802 35492 23808
rect 35820 23798 35848 24006
rect 35808 23792 35860 23798
rect 35808 23734 35860 23740
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 34244 22024 34296 22030
rect 34244 21966 34296 21972
rect 34532 21622 34560 22374
rect 34624 22166 34652 23666
rect 34704 23588 34756 23594
rect 34704 23530 34756 23536
rect 34716 22642 34744 23530
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34612 22160 34664 22166
rect 34612 22102 34664 22108
rect 34716 22030 34744 22374
rect 34808 22030 34836 22918
rect 35360 22778 35388 23054
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 22094 35388 22714
rect 35360 22066 35572 22094
rect 35544 22030 35572 22066
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 35348 22024 35400 22030
rect 35532 22024 35584 22030
rect 35400 21972 35480 21978
rect 35348 21966 35480 21972
rect 35532 21966 35584 21972
rect 34624 21876 34652 21966
rect 35360 21950 35480 21966
rect 34624 21848 34836 21876
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34428 21344 34480 21350
rect 34428 21286 34480 21292
rect 34348 21146 34376 21286
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 34336 21140 34388 21146
rect 34336 21082 34388 21088
rect 33980 20874 34008 21082
rect 34440 20874 34468 21286
rect 33968 20868 34020 20874
rect 33968 20810 34020 20816
rect 34428 20868 34480 20874
rect 34428 20810 34480 20816
rect 33980 20602 34008 20810
rect 34532 20806 34560 21558
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34520 20800 34572 20806
rect 34520 20742 34572 20748
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 34532 20466 34560 20742
rect 34624 20602 34652 20878
rect 34808 20806 34836 21848
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34716 20534 34744 20742
rect 34704 20528 34756 20534
rect 34704 20470 34756 20476
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34808 20330 34836 20742
rect 34060 20324 34112 20330
rect 34060 20266 34112 20272
rect 34796 20324 34848 20330
rect 34796 20266 34848 20272
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33796 19378 33824 19654
rect 33888 19514 33916 19654
rect 33876 19508 33928 19514
rect 33876 19450 33928 19456
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 32600 18970 32628 19314
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33704 18970 33732 19110
rect 32588 18964 32640 18970
rect 32588 18906 32640 18912
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 32784 15026 32812 15438
rect 32772 15020 32824 15026
rect 32772 14962 32824 14968
rect 32680 13728 32732 13734
rect 32680 13670 32732 13676
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31760 13252 31812 13258
rect 31760 13194 31812 13200
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 31482 12880 31538 12889
rect 31208 12844 31260 12850
rect 31482 12815 31538 12824
rect 31208 12786 31260 12792
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30760 10742 30788 11698
rect 31128 11098 31156 12174
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 31312 11218 31340 11494
rect 31300 11212 31352 11218
rect 31300 11154 31352 11160
rect 31036 11070 31156 11098
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30840 10668 30892 10674
rect 30892 10628 30972 10656
rect 30840 10610 30892 10616
rect 30392 9092 30420 10610
rect 30472 10464 30524 10470
rect 30472 10406 30524 10412
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30484 10062 30512 10406
rect 30472 10056 30524 10062
rect 30472 9998 30524 10004
rect 30484 9450 30512 9998
rect 30760 9926 30788 10406
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30472 9444 30524 9450
rect 30472 9386 30524 9392
rect 30668 9178 30696 9522
rect 30760 9364 30788 9862
rect 30852 9586 30880 10406
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30840 9376 30892 9382
rect 30760 9336 30840 9364
rect 30656 9172 30708 9178
rect 30656 9114 30708 9120
rect 30472 9104 30524 9110
rect 30392 9064 30472 9092
rect 30392 8974 30420 9064
rect 30472 9046 30524 9052
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30656 8900 30708 8906
rect 30656 8842 30708 8848
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30208 8022 30236 8434
rect 30196 8016 30248 8022
rect 30196 7958 30248 7964
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 29920 7812 29972 7818
rect 29920 7754 29972 7760
rect 29828 7744 29880 7750
rect 29828 7686 29880 7692
rect 29458 7375 29514 7384
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29840 7342 29868 7686
rect 29932 7410 29960 7754
rect 30116 7546 30144 7822
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30208 7478 30236 7822
rect 30196 7472 30248 7478
rect 30196 7414 30248 7420
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 29460 7336 29512 7342
rect 29460 7278 29512 7284
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29472 6730 29500 7278
rect 29552 7268 29604 7274
rect 29552 7210 29604 7216
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 29564 6730 29592 7210
rect 30116 6798 30144 7210
rect 30392 7002 30420 8434
rect 30484 7206 30512 8842
rect 30668 8634 30696 8842
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30760 7342 30788 9336
rect 30840 9318 30892 9324
rect 30944 8566 30972 10628
rect 31036 10266 31064 11070
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31128 10742 31156 10950
rect 31116 10736 31168 10742
rect 31116 10678 31168 10684
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 31220 10130 31248 10474
rect 31208 10124 31260 10130
rect 31208 10066 31260 10072
rect 31208 9376 31260 9382
rect 31208 9318 31260 9324
rect 31024 9104 31076 9110
rect 31024 9046 31076 9052
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30840 8424 30892 8430
rect 31036 8412 31064 9046
rect 31220 9042 31248 9318
rect 31208 9036 31260 9042
rect 31208 8978 31260 8984
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 31128 8430 31156 8774
rect 31312 8498 31340 11154
rect 31496 10606 31524 12582
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31588 11150 31616 11562
rect 31680 11150 31708 11698
rect 31576 11144 31628 11150
rect 31576 11086 31628 11092
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31484 10600 31536 10606
rect 31404 10560 31484 10588
rect 31404 9722 31432 10560
rect 31484 10542 31536 10548
rect 31588 9926 31616 11086
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 31576 9920 31628 9926
rect 31576 9862 31628 9868
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 30892 8384 31064 8412
rect 31116 8424 31168 8430
rect 30840 8366 30892 8372
rect 31116 8366 31168 8372
rect 30852 8022 30880 8366
rect 30840 8016 30892 8022
rect 30840 7958 30892 7964
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30472 7200 30524 7206
rect 30472 7142 30524 7148
rect 30564 7200 30616 7206
rect 30840 7200 30892 7206
rect 30564 7142 30616 7148
rect 30760 7148 30840 7154
rect 30760 7142 30892 7148
rect 30576 7002 30604 7142
rect 30760 7126 30880 7142
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30564 6996 30616 7002
rect 30564 6938 30616 6944
rect 30760 6798 30788 7126
rect 31036 7002 31064 7346
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 30840 6928 30892 6934
rect 30840 6870 30892 6876
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29552 6724 29604 6730
rect 29552 6666 29604 6672
rect 30852 6662 30880 6870
rect 31128 6798 31156 7278
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31220 6746 31248 8434
rect 31312 8090 31340 8434
rect 31404 8294 31432 9658
rect 31680 9518 31708 10610
rect 31772 10062 31800 13194
rect 32692 12918 32720 13670
rect 32876 13138 32904 18838
rect 33508 17808 33560 17814
rect 33508 17750 33560 17756
rect 33520 17202 33548 17750
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33612 17202 33640 17614
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33784 17196 33836 17202
rect 33784 17138 33836 17144
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 33060 16794 33088 16934
rect 33048 16788 33100 16794
rect 33048 16730 33100 16736
rect 32956 16516 33008 16522
rect 32956 16458 33008 16464
rect 32968 16250 32996 16458
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33060 15502 33088 16730
rect 33520 16726 33548 17138
rect 33612 16726 33640 17138
rect 33692 16992 33744 16998
rect 33796 16980 33824 17138
rect 33744 16952 33824 16980
rect 33692 16934 33744 16940
rect 33508 16720 33560 16726
rect 33508 16662 33560 16668
rect 33600 16720 33652 16726
rect 33600 16662 33652 16668
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33244 15706 33272 16050
rect 33336 15706 33364 16050
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33600 15904 33652 15910
rect 33600 15846 33652 15852
rect 33232 15700 33284 15706
rect 33232 15642 33284 15648
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33520 15570 33548 15846
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33048 15496 33100 15502
rect 33048 15438 33100 15444
rect 33612 14958 33640 15846
rect 33704 15502 33732 16934
rect 33784 16448 33836 16454
rect 33784 16390 33836 16396
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33796 15706 33824 16390
rect 33888 16114 33916 16390
rect 34072 16114 34100 20266
rect 34336 20256 34388 20262
rect 34336 20198 34388 20204
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34348 17354 34376 20198
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 19378 34468 19654
rect 34532 19514 34560 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34520 19508 34572 19514
rect 34520 19450 34572 19456
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34164 17338 34376 17354
rect 34440 17338 34468 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35452 18766 35480 21950
rect 35636 21010 35664 23462
rect 35820 22710 35848 23734
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35820 22234 35848 22646
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35624 21004 35676 21010
rect 35624 20946 35676 20952
rect 35900 20256 35952 20262
rect 35952 20204 36032 20210
rect 35900 20198 36032 20204
rect 35912 20182 36032 20198
rect 36004 19854 36032 20182
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 35808 19168 35860 19174
rect 35808 19110 35860 19116
rect 35716 18896 35768 18902
rect 35716 18838 35768 18844
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 35440 18760 35492 18766
rect 35440 18702 35492 18708
rect 34716 18086 34744 18702
rect 35728 18222 35756 18838
rect 35820 18766 35848 19110
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 35716 18216 35768 18222
rect 35716 18158 35768 18164
rect 36004 18086 36032 19790
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 35992 18080 36044 18086
rect 35992 18022 36044 18028
rect 34152 17332 34376 17338
rect 34204 17326 34376 17332
rect 34152 17274 34204 17280
rect 34348 17202 34376 17326
rect 34428 17332 34480 17338
rect 34428 17274 34480 17280
rect 34716 17202 34744 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 36004 17542 36032 18022
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 34152 17196 34204 17202
rect 34152 17138 34204 17144
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34164 16794 34192 17138
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34152 16788 34204 16794
rect 34152 16730 34204 16736
rect 34532 16726 34560 16934
rect 34520 16720 34572 16726
rect 34520 16662 34572 16668
rect 34716 16590 34744 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34704 16584 34756 16590
rect 34704 16526 34756 16532
rect 35716 16448 35768 16454
rect 35716 16390 35768 16396
rect 35728 16250 35756 16390
rect 35716 16244 35768 16250
rect 35716 16186 35768 16192
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 34060 16108 34112 16114
rect 34060 16050 34112 16056
rect 33784 15700 33836 15706
rect 33784 15642 33836 15648
rect 33888 15570 33916 16050
rect 34612 16040 34664 16046
rect 34612 15982 34664 15988
rect 34624 15570 34652 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33876 15564 33928 15570
rect 33876 15506 33928 15512
rect 34612 15564 34664 15570
rect 34612 15506 34664 15512
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33600 14952 33652 14958
rect 33600 14894 33652 14900
rect 34624 14890 34652 15506
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 34612 14884 34664 14890
rect 34612 14826 34664 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14618 35388 15438
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35452 15094 35480 15302
rect 36004 15162 36032 17478
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 36096 14822 36124 30790
rect 36452 30592 36504 30598
rect 36452 30534 36504 30540
rect 36464 30258 36492 30534
rect 36556 30258 36584 31758
rect 36740 30394 36768 31776
rect 36820 31758 36872 31764
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36832 30870 36860 31622
rect 36820 30864 36872 30870
rect 36820 30806 36872 30812
rect 36728 30388 36780 30394
rect 36728 30330 36780 30336
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36728 30184 36780 30190
rect 36728 30126 36780 30132
rect 36544 29096 36596 29102
rect 36544 29038 36596 29044
rect 36556 28218 36584 29038
rect 36544 28212 36596 28218
rect 36544 28154 36596 28160
rect 36176 28076 36228 28082
rect 36176 28018 36228 28024
rect 36188 27606 36216 28018
rect 36176 27600 36228 27606
rect 36176 27542 36228 27548
rect 36188 26790 36216 27542
rect 36740 27334 36768 30126
rect 36912 30048 36964 30054
rect 36912 29990 36964 29996
rect 36924 28762 36952 29990
rect 36912 28756 36964 28762
rect 36912 28698 36964 28704
rect 36924 28014 36952 28698
rect 36912 28008 36964 28014
rect 36912 27950 36964 27956
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36740 26994 36768 27270
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 36452 26784 36504 26790
rect 36452 26726 36504 26732
rect 36464 26586 36492 26726
rect 36452 26580 36504 26586
rect 36452 26522 36504 26528
rect 37016 24818 37044 44746
rect 43444 43716 43496 43722
rect 43444 43658 43496 43664
rect 44640 43716 44692 43722
rect 44640 43658 44692 43664
rect 37832 43648 37884 43654
rect 37832 43590 37884 43596
rect 37096 42696 37148 42702
rect 37096 42638 37148 42644
rect 37108 41274 37136 42638
rect 37280 41812 37332 41818
rect 37280 41754 37332 41760
rect 37096 41268 37148 41274
rect 37096 41210 37148 41216
rect 37292 41138 37320 41754
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37556 41064 37608 41070
rect 37556 41006 37608 41012
rect 37568 40730 37596 41006
rect 37556 40724 37608 40730
rect 37556 40666 37608 40672
rect 37372 40384 37424 40390
rect 37372 40326 37424 40332
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 37292 38350 37320 38694
rect 37384 38350 37412 40326
rect 37844 38706 37872 43590
rect 40592 43376 40644 43382
rect 40592 43318 40644 43324
rect 38660 43240 38712 43246
rect 38660 43182 38712 43188
rect 39212 43240 39264 43246
rect 39212 43182 39264 43188
rect 38672 42650 38700 43182
rect 39224 42906 39252 43182
rect 39212 42900 39264 42906
rect 39212 42842 39264 42848
rect 38844 42764 38896 42770
rect 38844 42706 38896 42712
rect 38488 42622 38700 42650
rect 38488 42158 38516 42622
rect 38856 42378 38884 42706
rect 40316 42560 40368 42566
rect 40316 42502 40368 42508
rect 38856 42362 38976 42378
rect 40328 42362 40356 42502
rect 38844 42356 38976 42362
rect 38896 42350 38976 42356
rect 38844 42298 38896 42304
rect 38844 42220 38896 42226
rect 38844 42162 38896 42168
rect 38476 42152 38528 42158
rect 38476 42094 38528 42100
rect 38488 41818 38516 42094
rect 38476 41812 38528 41818
rect 38476 41754 38528 41760
rect 38200 41608 38252 41614
rect 38200 41550 38252 41556
rect 38212 41414 38240 41550
rect 38212 41386 38424 41414
rect 38108 39296 38160 39302
rect 38108 39238 38160 39244
rect 38200 39296 38252 39302
rect 38200 39238 38252 39244
rect 38120 38894 38148 39238
rect 38108 38888 38160 38894
rect 38108 38830 38160 38836
rect 37844 38678 38148 38706
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 37372 38344 37424 38350
rect 37372 38286 37424 38292
rect 37924 38344 37976 38350
rect 37924 38286 37976 38292
rect 37292 37806 37320 38286
rect 37936 38010 37964 38286
rect 37924 38004 37976 38010
rect 37924 37946 37976 37952
rect 37280 37800 37332 37806
rect 37280 37742 37332 37748
rect 38016 37800 38068 37806
rect 38016 37742 38068 37748
rect 37832 37664 37884 37670
rect 37832 37606 37884 37612
rect 37844 37330 37872 37606
rect 37832 37324 37884 37330
rect 37832 37266 37884 37272
rect 38028 37262 38056 37742
rect 38016 37256 38068 37262
rect 38016 37198 38068 37204
rect 38028 36786 38056 37198
rect 38016 36780 38068 36786
rect 38016 36722 38068 36728
rect 37740 36576 37792 36582
rect 37740 36518 37792 36524
rect 37752 36242 37780 36518
rect 37740 36236 37792 36242
rect 37740 36178 37792 36184
rect 37096 36168 37148 36174
rect 37096 36110 37148 36116
rect 37108 35630 37136 36110
rect 37096 35624 37148 35630
rect 37096 35566 37148 35572
rect 37648 34944 37700 34950
rect 37648 34886 37700 34892
rect 37660 34746 37688 34886
rect 37648 34740 37700 34746
rect 37648 34682 37700 34688
rect 37924 34740 37976 34746
rect 37924 34682 37976 34688
rect 37648 34400 37700 34406
rect 37648 34342 37700 34348
rect 37280 34128 37332 34134
rect 37280 34070 37332 34076
rect 37292 33658 37320 34070
rect 37280 33652 37332 33658
rect 37280 33594 37332 33600
rect 37660 32910 37688 34342
rect 37648 32904 37700 32910
rect 37648 32846 37700 32852
rect 37464 32020 37516 32026
rect 37464 31962 37516 31968
rect 37476 31754 37504 31962
rect 37464 31748 37516 31754
rect 37464 31690 37516 31696
rect 37280 28144 37332 28150
rect 37200 28092 37280 28098
rect 37200 28086 37332 28092
rect 37200 28070 37320 28086
rect 37200 27946 37228 28070
rect 37556 28008 37608 28014
rect 37556 27950 37608 27956
rect 37188 27940 37240 27946
rect 37188 27882 37240 27888
rect 37464 27532 37516 27538
rect 37464 27474 37516 27480
rect 37476 27130 37504 27474
rect 37568 27130 37596 27950
rect 37660 27674 37688 32846
rect 37936 31142 37964 34682
rect 38016 34604 38068 34610
rect 38016 34546 38068 34552
rect 38028 32230 38056 34546
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 38016 31884 38068 31890
rect 38016 31826 38068 31832
rect 38028 31346 38056 31826
rect 38120 31770 38148 38678
rect 38212 37670 38240 39238
rect 38396 39098 38424 41386
rect 38488 39982 38516 41754
rect 38856 41274 38884 42162
rect 38948 41818 38976 42350
rect 40316 42356 40368 42362
rect 40316 42298 40368 42304
rect 40604 42294 40632 43318
rect 40684 43104 40736 43110
rect 40684 43046 40736 43052
rect 40696 42770 40724 43046
rect 43456 42906 43484 43658
rect 44652 43625 44680 43658
rect 44638 43616 44694 43625
rect 44638 43551 44694 43560
rect 43444 42900 43496 42906
rect 43444 42842 43496 42848
rect 40684 42764 40736 42770
rect 40684 42706 40736 42712
rect 40592 42288 40644 42294
rect 40592 42230 40644 42236
rect 39396 42220 39448 42226
rect 39396 42162 39448 42168
rect 38936 41812 38988 41818
rect 38936 41754 38988 41760
rect 39408 41478 39436 42162
rect 40604 42158 40632 42230
rect 40592 42152 40644 42158
rect 40592 42094 40644 42100
rect 39948 41608 40000 41614
rect 39948 41550 40000 41556
rect 40314 41576 40370 41585
rect 39488 41540 39540 41546
rect 39488 41482 39540 41488
rect 39120 41472 39172 41478
rect 39120 41414 39172 41420
rect 39304 41472 39356 41478
rect 39304 41414 39356 41420
rect 39396 41472 39448 41478
rect 39396 41414 39448 41420
rect 38844 41268 38896 41274
rect 38844 41210 38896 41216
rect 39132 40526 39160 41414
rect 39316 41274 39344 41414
rect 39304 41268 39356 41274
rect 39304 41210 39356 41216
rect 39408 41206 39436 41414
rect 39396 41200 39448 41206
rect 39396 41142 39448 41148
rect 39120 40520 39172 40526
rect 39120 40462 39172 40468
rect 38476 39976 38528 39982
rect 38476 39918 38528 39924
rect 38752 39976 38804 39982
rect 38752 39918 38804 39924
rect 38764 39642 38792 39918
rect 38752 39636 38804 39642
rect 38752 39578 38804 39584
rect 38752 39432 38804 39438
rect 38752 39374 38804 39380
rect 38384 39092 38436 39098
rect 38384 39034 38436 39040
rect 38292 39024 38344 39030
rect 38292 38966 38344 38972
rect 38304 38758 38332 38966
rect 38292 38752 38344 38758
rect 38292 38694 38344 38700
rect 38304 38418 38332 38694
rect 38292 38412 38344 38418
rect 38292 38354 38344 38360
rect 38200 37664 38252 37670
rect 38200 37606 38252 37612
rect 38396 34610 38424 39034
rect 38660 38208 38712 38214
rect 38660 38150 38712 38156
rect 38672 38010 38700 38150
rect 38764 38010 38792 39374
rect 38660 38004 38712 38010
rect 38660 37946 38712 37952
rect 38752 38004 38804 38010
rect 38752 37946 38804 37952
rect 39500 37806 39528 41482
rect 39960 41478 39988 41550
rect 40696 41546 40724 42706
rect 40776 42696 40828 42702
rect 40776 42638 40828 42644
rect 40314 41511 40316 41520
rect 40368 41511 40370 41520
rect 40408 41540 40460 41546
rect 40316 41482 40368 41488
rect 40408 41482 40460 41488
rect 40684 41540 40736 41546
rect 40684 41482 40736 41488
rect 39948 41472 40000 41478
rect 39948 41414 40000 41420
rect 40040 41472 40092 41478
rect 40040 41414 40092 41420
rect 39960 39642 39988 41414
rect 40052 41138 40080 41414
rect 40420 41206 40448 41482
rect 40408 41200 40460 41206
rect 40408 41142 40460 41148
rect 40040 41132 40092 41138
rect 40040 41074 40092 41080
rect 40420 40730 40448 41142
rect 40696 40730 40724 41482
rect 40788 41274 40816 42638
rect 42248 42220 42300 42226
rect 42248 42162 42300 42168
rect 41144 42152 41196 42158
rect 41144 42094 41196 42100
rect 40868 41812 40920 41818
rect 40868 41754 40920 41760
rect 40880 41614 40908 41754
rect 40960 41744 41012 41750
rect 41012 41692 41092 41698
rect 40960 41686 41092 41692
rect 40972 41670 41092 41686
rect 40868 41608 40920 41614
rect 40868 41550 40920 41556
rect 40960 41608 41012 41614
rect 40960 41550 41012 41556
rect 40776 41268 40828 41274
rect 40776 41210 40828 41216
rect 40972 41206 41000 41550
rect 40960 41200 41012 41206
rect 40960 41142 41012 41148
rect 41064 41002 41092 41670
rect 41156 41070 41184 42094
rect 41236 42016 41288 42022
rect 41236 41958 41288 41964
rect 41604 42016 41656 42022
rect 41604 41958 41656 41964
rect 41248 41818 41276 41958
rect 41236 41812 41288 41818
rect 41236 41754 41288 41760
rect 41616 41682 41644 41958
rect 42260 41818 42288 42162
rect 42432 42152 42484 42158
rect 42432 42094 42484 42100
rect 42340 42016 42392 42022
rect 42340 41958 42392 41964
rect 42248 41812 42300 41818
rect 42248 41754 42300 41760
rect 41604 41676 41656 41682
rect 41604 41618 41656 41624
rect 41616 41585 41644 41618
rect 41602 41576 41658 41585
rect 41328 41540 41380 41546
rect 41602 41511 41658 41520
rect 41788 41540 41840 41546
rect 41328 41482 41380 41488
rect 41788 41482 41840 41488
rect 41340 41138 41368 41482
rect 41328 41132 41380 41138
rect 41328 41074 41380 41080
rect 41800 41070 41828 41482
rect 42064 41472 42116 41478
rect 42064 41414 42116 41420
rect 42076 41274 42104 41414
rect 42064 41268 42116 41274
rect 42064 41210 42116 41216
rect 42352 41138 42380 41958
rect 42444 41682 42472 42094
rect 42432 41676 42484 41682
rect 42432 41618 42484 41624
rect 43352 41676 43404 41682
rect 43352 41618 43404 41624
rect 42340 41132 42392 41138
rect 42340 41074 42392 41080
rect 41144 41064 41196 41070
rect 41144 41006 41196 41012
rect 41788 41064 41840 41070
rect 41788 41006 41840 41012
rect 41052 40996 41104 41002
rect 41052 40938 41104 40944
rect 40408 40724 40460 40730
rect 40408 40666 40460 40672
rect 40684 40724 40736 40730
rect 40684 40666 40736 40672
rect 40592 40520 40644 40526
rect 40592 40462 40644 40468
rect 40132 40384 40184 40390
rect 40132 40326 40184 40332
rect 40144 39642 40172 40326
rect 40604 40050 40632 40462
rect 40776 40384 40828 40390
rect 40776 40326 40828 40332
rect 40788 40050 40816 40326
rect 41156 40118 41184 41006
rect 41880 40928 41932 40934
rect 41880 40870 41932 40876
rect 41144 40112 41196 40118
rect 41144 40054 41196 40060
rect 41892 40050 41920 40870
rect 40592 40044 40644 40050
rect 40592 39986 40644 39992
rect 40776 40044 40828 40050
rect 40776 39986 40828 39992
rect 41880 40044 41932 40050
rect 41880 39986 41932 39992
rect 39948 39636 40000 39642
rect 39948 39578 40000 39584
rect 40132 39636 40184 39642
rect 40132 39578 40184 39584
rect 40144 38894 40172 39578
rect 40224 39432 40276 39438
rect 40224 39374 40276 39380
rect 39856 38888 39908 38894
rect 39856 38830 39908 38836
rect 40132 38888 40184 38894
rect 40132 38830 40184 38836
rect 39868 38350 39896 38830
rect 40236 38758 40264 39374
rect 40604 39370 40632 39986
rect 41144 39840 41196 39846
rect 41144 39782 41196 39788
rect 41236 39840 41288 39846
rect 41236 39782 41288 39788
rect 41156 39438 41184 39782
rect 41144 39432 41196 39438
rect 41144 39374 41196 39380
rect 40592 39364 40644 39370
rect 40592 39306 40644 39312
rect 40316 39296 40368 39302
rect 40316 39238 40368 39244
rect 40328 38962 40356 39238
rect 40316 38956 40368 38962
rect 40316 38898 40368 38904
rect 40868 38956 40920 38962
rect 40868 38898 40920 38904
rect 40316 38820 40368 38826
rect 40316 38762 40368 38768
rect 40224 38752 40276 38758
rect 40224 38694 40276 38700
rect 39856 38344 39908 38350
rect 39856 38286 39908 38292
rect 39488 37800 39540 37806
rect 39488 37742 39540 37748
rect 38660 37664 38712 37670
rect 38660 37606 38712 37612
rect 38844 37664 38896 37670
rect 38844 37606 38896 37612
rect 38672 37262 38700 37606
rect 38856 37262 38884 37606
rect 39500 37466 39528 37742
rect 39488 37460 39540 37466
rect 39488 37402 39540 37408
rect 38660 37256 38712 37262
rect 38660 37198 38712 37204
rect 38844 37256 38896 37262
rect 38844 37198 38896 37204
rect 38672 36786 38700 37198
rect 38660 36780 38712 36786
rect 38660 36722 38712 36728
rect 38856 36718 38884 37198
rect 38844 36712 38896 36718
rect 38844 36654 38896 36660
rect 38856 36378 38884 36654
rect 38844 36372 38896 36378
rect 38844 36314 38896 36320
rect 39580 36168 39632 36174
rect 39580 36110 39632 36116
rect 38844 36032 38896 36038
rect 38844 35974 38896 35980
rect 38856 35562 38884 35974
rect 39396 35624 39448 35630
rect 39396 35566 39448 35572
rect 38844 35556 38896 35562
rect 38844 35498 38896 35504
rect 39408 35494 39436 35566
rect 39396 35488 39448 35494
rect 39396 35430 39448 35436
rect 38752 35148 38804 35154
rect 38752 35090 38804 35096
rect 38384 34604 38436 34610
rect 38384 34546 38436 34552
rect 38476 34400 38528 34406
rect 38476 34342 38528 34348
rect 38488 34066 38516 34342
rect 38476 34060 38528 34066
rect 38476 34002 38528 34008
rect 38488 33946 38516 34002
rect 38396 33918 38516 33946
rect 38292 33584 38344 33590
rect 38292 33526 38344 33532
rect 38304 33114 38332 33526
rect 38396 33318 38424 33918
rect 38764 33862 38792 35090
rect 39120 35080 39172 35086
rect 39120 35022 39172 35028
rect 39132 34746 39160 35022
rect 39120 34740 39172 34746
rect 39120 34682 39172 34688
rect 39408 34406 39436 35430
rect 39592 35290 39620 36110
rect 39764 36032 39816 36038
rect 39764 35974 39816 35980
rect 39776 35834 39804 35974
rect 39764 35828 39816 35834
rect 39764 35770 39816 35776
rect 39868 35494 39896 38286
rect 40040 38276 40092 38282
rect 40040 38218 40092 38224
rect 40132 38276 40184 38282
rect 40132 38218 40184 38224
rect 39948 37800 40000 37806
rect 39948 37742 40000 37748
rect 39960 36650 39988 37742
rect 40052 37262 40080 38218
rect 40144 38010 40172 38218
rect 40132 38004 40184 38010
rect 40132 37946 40184 37952
rect 40236 37874 40264 38694
rect 40328 37874 40356 38762
rect 40880 38554 40908 38898
rect 40868 38548 40920 38554
rect 40868 38490 40920 38496
rect 40224 37868 40276 37874
rect 40224 37810 40276 37816
rect 40316 37868 40368 37874
rect 40316 37810 40368 37816
rect 41248 37330 41276 39782
rect 42444 39506 42472 41618
rect 43076 41540 43128 41546
rect 43076 41482 43128 41488
rect 42708 41200 42760 41206
rect 42708 41142 42760 41148
rect 42524 41064 42576 41070
rect 42524 41006 42576 41012
rect 42536 40526 42564 41006
rect 42720 40730 42748 41142
rect 42800 40928 42852 40934
rect 42800 40870 42852 40876
rect 42708 40724 42760 40730
rect 42708 40666 42760 40672
rect 42524 40520 42576 40526
rect 42524 40462 42576 40468
rect 42812 39982 42840 40870
rect 42800 39976 42852 39982
rect 42800 39918 42852 39924
rect 42812 39642 42840 39918
rect 42892 39840 42944 39846
rect 42892 39782 42944 39788
rect 42904 39642 42932 39782
rect 42800 39636 42852 39642
rect 42800 39578 42852 39584
rect 42892 39636 42944 39642
rect 42892 39578 42944 39584
rect 42432 39500 42484 39506
rect 42432 39442 42484 39448
rect 42156 39432 42208 39438
rect 42156 39374 42208 39380
rect 42524 39432 42576 39438
rect 42524 39374 42576 39380
rect 42168 38214 42196 39374
rect 42536 38554 42564 39374
rect 42524 38548 42576 38554
rect 42524 38490 42576 38496
rect 42812 38418 42840 39578
rect 42708 38412 42760 38418
rect 42708 38354 42760 38360
rect 42800 38412 42852 38418
rect 42800 38354 42852 38360
rect 42616 38344 42668 38350
rect 42616 38286 42668 38292
rect 42156 38208 42208 38214
rect 42156 38150 42208 38156
rect 41236 37324 41288 37330
rect 41236 37266 41288 37272
rect 40040 37256 40092 37262
rect 40040 37198 40092 37204
rect 41248 37126 41276 37266
rect 41144 37120 41196 37126
rect 41144 37062 41196 37068
rect 41236 37120 41288 37126
rect 41236 37062 41288 37068
rect 41420 37120 41472 37126
rect 41420 37062 41472 37068
rect 41604 37120 41656 37126
rect 41604 37062 41656 37068
rect 41788 37120 41840 37126
rect 41788 37062 41840 37068
rect 39948 36644 40000 36650
rect 39948 36586 40000 36592
rect 40132 36644 40184 36650
rect 40132 36586 40184 36592
rect 40144 36242 40172 36586
rect 40132 36236 40184 36242
rect 40132 36178 40184 36184
rect 39948 36168 40000 36174
rect 39948 36110 40000 36116
rect 39856 35488 39908 35494
rect 39856 35430 39908 35436
rect 39960 35290 39988 36110
rect 40144 35894 40172 36178
rect 40052 35866 40172 35894
rect 39580 35284 39632 35290
rect 39580 35226 39632 35232
rect 39948 35284 40000 35290
rect 39948 35226 40000 35232
rect 39856 35216 39908 35222
rect 39856 35158 39908 35164
rect 39764 35080 39816 35086
rect 39764 35022 39816 35028
rect 39488 34944 39540 34950
rect 39776 34932 39804 35022
rect 39540 34904 39804 34932
rect 39488 34886 39540 34892
rect 39500 34610 39528 34886
rect 39488 34604 39540 34610
rect 39488 34546 39540 34552
rect 39396 34400 39448 34406
rect 39396 34342 39448 34348
rect 39500 34202 39528 34546
rect 39488 34196 39540 34202
rect 39488 34138 39540 34144
rect 39868 33998 39896 35158
rect 39856 33992 39908 33998
rect 39856 33934 39908 33940
rect 38752 33856 38804 33862
rect 38752 33798 38804 33804
rect 39764 33856 39816 33862
rect 39764 33798 39816 33804
rect 39776 33658 39804 33798
rect 39764 33652 39816 33658
rect 39764 33594 39816 33600
rect 39776 33318 39804 33594
rect 38384 33312 38436 33318
rect 38384 33254 38436 33260
rect 39764 33312 39816 33318
rect 39764 33254 39816 33260
rect 38292 33108 38344 33114
rect 38292 33050 38344 33056
rect 38396 31890 38424 33254
rect 38568 32904 38620 32910
rect 38568 32846 38620 32852
rect 38580 31890 38608 32846
rect 39396 32836 39448 32842
rect 39396 32778 39448 32784
rect 38384 31884 38436 31890
rect 38384 31826 38436 31832
rect 38568 31884 38620 31890
rect 38568 31826 38620 31832
rect 38120 31742 38700 31770
rect 38108 31680 38160 31686
rect 38108 31622 38160 31628
rect 38016 31340 38068 31346
rect 38016 31282 38068 31288
rect 37924 31136 37976 31142
rect 37924 31078 37976 31084
rect 37936 30734 37964 31078
rect 37924 30728 37976 30734
rect 37924 30670 37976 30676
rect 38016 30660 38068 30666
rect 38016 30602 38068 30608
rect 37832 30252 37884 30258
rect 37832 30194 37884 30200
rect 37844 29306 37872 30194
rect 38028 30122 38056 30602
rect 38016 30116 38068 30122
rect 38016 30058 38068 30064
rect 38028 29578 38056 30058
rect 38120 30054 38148 31622
rect 38476 31340 38528 31346
rect 38476 31282 38528 31288
rect 38384 31272 38436 31278
rect 38384 31214 38436 31220
rect 38396 30938 38424 31214
rect 38384 30932 38436 30938
rect 38384 30874 38436 30880
rect 38200 30728 38252 30734
rect 38200 30670 38252 30676
rect 38212 30394 38240 30670
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 38108 30048 38160 30054
rect 38108 29990 38160 29996
rect 38016 29572 38068 29578
rect 38016 29514 38068 29520
rect 37832 29300 37884 29306
rect 37832 29242 37884 29248
rect 37832 29096 37884 29102
rect 37832 29038 37884 29044
rect 37844 28558 37872 29038
rect 38212 29034 38332 29050
rect 38200 29028 38332 29034
rect 38252 29022 38332 29028
rect 38200 28970 38252 28976
rect 37924 28756 37976 28762
rect 37924 28698 37976 28704
rect 37832 28552 37884 28558
rect 37832 28494 37884 28500
rect 37648 27668 37700 27674
rect 37648 27610 37700 27616
rect 37740 27600 37792 27606
rect 37740 27542 37792 27548
rect 37752 27402 37780 27542
rect 37740 27396 37792 27402
rect 37740 27338 37792 27344
rect 37464 27124 37516 27130
rect 37464 27066 37516 27072
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 37476 26994 37504 27066
rect 37752 27062 37780 27338
rect 37740 27056 37792 27062
rect 37740 26998 37792 27004
rect 37936 26994 37964 28698
rect 38200 28416 38252 28422
rect 38200 28358 38252 28364
rect 38212 28218 38240 28358
rect 38200 28212 38252 28218
rect 38200 28154 38252 28160
rect 38016 28144 38068 28150
rect 38016 28086 38068 28092
rect 38028 28014 38056 28086
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 38108 27872 38160 27878
rect 38108 27814 38160 27820
rect 38120 27334 38148 27814
rect 38108 27328 38160 27334
rect 38108 27270 38160 27276
rect 37372 26988 37424 26994
rect 37372 26930 37424 26936
rect 37464 26988 37516 26994
rect 37464 26930 37516 26936
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37924 26988 37976 26994
rect 37924 26930 37976 26936
rect 37096 26376 37148 26382
rect 37096 26318 37148 26324
rect 37108 26042 37136 26318
rect 37096 26036 37148 26042
rect 37096 25978 37148 25984
rect 37384 25906 37412 26930
rect 37660 26314 37688 26930
rect 37844 26586 37872 26930
rect 37832 26580 37884 26586
rect 37832 26522 37884 26528
rect 38016 26376 38068 26382
rect 38016 26318 38068 26324
rect 37648 26308 37700 26314
rect 37648 26250 37700 26256
rect 37372 25900 37424 25906
rect 37372 25842 37424 25848
rect 37280 25696 37332 25702
rect 37280 25638 37332 25644
rect 37292 25498 37320 25638
rect 37280 25492 37332 25498
rect 37280 25434 37332 25440
rect 37004 24812 37056 24818
rect 37004 24754 37056 24760
rect 36912 24608 36964 24614
rect 36912 24550 36964 24556
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 36280 20466 36308 22170
rect 36372 21690 36400 24142
rect 36924 23866 36952 24550
rect 37556 24200 37608 24206
rect 37556 24142 37608 24148
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 37372 24064 37424 24070
rect 37372 24006 37424 24012
rect 36912 23860 36964 23866
rect 36912 23802 36964 23808
rect 37096 23656 37148 23662
rect 37096 23598 37148 23604
rect 37108 23322 37136 23598
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 37108 22642 37136 23258
rect 37292 23050 37320 24006
rect 37384 23186 37412 24006
rect 37372 23180 37424 23186
rect 37372 23122 37424 23128
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 37568 22778 37596 24142
rect 37556 22772 37608 22778
rect 37556 22714 37608 22720
rect 37096 22636 37148 22642
rect 37096 22578 37148 22584
rect 36820 22568 36872 22574
rect 36820 22510 36872 22516
rect 36832 21894 36860 22510
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36360 21684 36412 21690
rect 36360 21626 36412 21632
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36648 20602 36676 20878
rect 37660 20602 37688 26250
rect 38028 25158 38056 26318
rect 38120 26314 38148 27270
rect 38212 27062 38240 28154
rect 38200 27056 38252 27062
rect 38200 26998 38252 27004
rect 38108 26308 38160 26314
rect 38108 26250 38160 26256
rect 38120 25838 38148 26250
rect 38108 25832 38160 25838
rect 38108 25774 38160 25780
rect 38120 25362 38148 25774
rect 38108 25356 38160 25362
rect 38108 25298 38160 25304
rect 38016 25152 38068 25158
rect 38016 25094 38068 25100
rect 38028 22710 38056 25094
rect 38016 22704 38068 22710
rect 38016 22646 38068 22652
rect 38108 22568 38160 22574
rect 38108 22510 38160 22516
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36556 19922 36584 20266
rect 36648 20058 36676 20538
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 36636 20052 36688 20058
rect 36636 19994 36688 20000
rect 36544 19916 36596 19922
rect 36544 19858 36596 19864
rect 37476 19786 37504 20402
rect 37556 20392 37608 20398
rect 37556 20334 37608 20340
rect 37464 19780 37516 19786
rect 37464 19722 37516 19728
rect 37476 18222 37504 19722
rect 37568 18630 37596 20334
rect 38016 19712 38068 19718
rect 38016 19654 38068 19660
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37844 18698 37872 19110
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37936 18426 37964 18770
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37188 18148 37240 18154
rect 37188 18090 37240 18096
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 37016 17202 37044 17614
rect 37200 17542 37228 18090
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37372 18080 37424 18086
rect 37372 18022 37424 18028
rect 37292 17746 37320 18022
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37004 17196 37056 17202
rect 37004 17138 37056 17144
rect 37200 17134 37228 17478
rect 37384 17338 37412 18022
rect 37372 17332 37424 17338
rect 37372 17274 37424 17280
rect 37188 17128 37240 17134
rect 37188 17070 37240 17076
rect 37200 15434 37228 17070
rect 37476 16522 37504 18158
rect 37464 16516 37516 16522
rect 37464 16458 37516 16464
rect 38028 15706 38056 19654
rect 38016 15700 38068 15706
rect 38016 15642 38068 15648
rect 38016 15564 38068 15570
rect 38016 15506 38068 15512
rect 37188 15428 37240 15434
rect 37188 15370 37240 15376
rect 37200 14958 37228 15370
rect 38028 15162 38056 15506
rect 38120 15366 38148 22510
rect 38304 22094 38332 29022
rect 38396 27606 38424 30874
rect 38488 30394 38516 31282
rect 38568 30660 38620 30666
rect 38568 30602 38620 30608
rect 38476 30388 38528 30394
rect 38476 30330 38528 30336
rect 38580 29850 38608 30602
rect 38568 29844 38620 29850
rect 38568 29786 38620 29792
rect 38476 29572 38528 29578
rect 38476 29514 38528 29520
rect 38384 27600 38436 27606
rect 38384 27542 38436 27548
rect 38488 27402 38516 29514
rect 38672 29170 38700 31742
rect 39212 31680 39264 31686
rect 39212 31622 39264 31628
rect 39224 31414 39252 31622
rect 38752 31408 38804 31414
rect 39212 31408 39264 31414
rect 38752 31350 38804 31356
rect 39132 31368 39212 31396
rect 38764 30938 38792 31350
rect 38752 30932 38804 30938
rect 38752 30874 38804 30880
rect 38752 30728 38804 30734
rect 38752 30670 38804 30676
rect 38764 29646 38792 30670
rect 39132 30598 39160 31368
rect 39212 31350 39264 31356
rect 39304 30660 39356 30666
rect 39304 30602 39356 30608
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 39120 30592 39172 30598
rect 39120 30534 39172 30540
rect 38856 30394 38884 30534
rect 38844 30388 38896 30394
rect 38844 30330 38896 30336
rect 39132 30326 39160 30534
rect 39316 30410 39344 30602
rect 39224 30382 39344 30410
rect 39120 30320 39172 30326
rect 39120 30262 39172 30268
rect 39224 30054 39252 30382
rect 39212 30048 39264 30054
rect 39212 29990 39264 29996
rect 38752 29640 38804 29646
rect 38752 29582 38804 29588
rect 39120 29640 39172 29646
rect 39120 29582 39172 29588
rect 38844 29572 38896 29578
rect 38844 29514 38896 29520
rect 38660 29164 38712 29170
rect 38660 29106 38712 29112
rect 38856 28966 38884 29514
rect 38936 29504 38988 29510
rect 38936 29446 38988 29452
rect 38948 29238 38976 29446
rect 38936 29232 38988 29238
rect 38936 29174 38988 29180
rect 38948 28966 38976 29174
rect 38844 28960 38896 28966
rect 38844 28902 38896 28908
rect 38936 28960 38988 28966
rect 38936 28902 38988 28908
rect 38568 28552 38620 28558
rect 38568 28494 38620 28500
rect 38580 27946 38608 28494
rect 38844 28416 38896 28422
rect 38844 28358 38896 28364
rect 38568 27940 38620 27946
rect 38568 27882 38620 27888
rect 38856 27470 38884 28358
rect 39132 27470 39160 29582
rect 39304 29164 39356 29170
rect 39304 29106 39356 29112
rect 39212 29028 39264 29034
rect 39212 28970 39264 28976
rect 39224 27878 39252 28970
rect 39316 28082 39344 29106
rect 39304 28076 39356 28082
rect 39304 28018 39356 28024
rect 39212 27872 39264 27878
rect 39212 27814 39264 27820
rect 38660 27464 38712 27470
rect 38660 27406 38712 27412
rect 38844 27464 38896 27470
rect 38844 27406 38896 27412
rect 39120 27464 39172 27470
rect 39120 27406 39172 27412
rect 38476 27396 38528 27402
rect 38476 27338 38528 27344
rect 38672 27130 38700 27406
rect 38660 27124 38712 27130
rect 38660 27066 38712 27072
rect 38384 25832 38436 25838
rect 38384 25774 38436 25780
rect 38396 25498 38424 25774
rect 38384 25492 38436 25498
rect 38384 25434 38436 25440
rect 38672 23798 38700 27066
rect 39132 27062 39160 27406
rect 39224 27402 39252 27814
rect 39212 27396 39264 27402
rect 39212 27338 39264 27344
rect 39120 27056 39172 27062
rect 39120 26998 39172 27004
rect 39304 24744 39356 24750
rect 39304 24686 39356 24692
rect 39028 24608 39080 24614
rect 39028 24550 39080 24556
rect 39040 24342 39068 24550
rect 39028 24336 39080 24342
rect 39028 24278 39080 24284
rect 39212 24064 39264 24070
rect 39212 24006 39264 24012
rect 39224 23866 39252 24006
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 38660 23792 38712 23798
rect 38660 23734 38712 23740
rect 39316 23610 39344 24686
rect 39408 24410 39436 32778
rect 39488 32020 39540 32026
rect 39488 31962 39540 31968
rect 39500 30734 39528 31962
rect 39776 31890 39804 33254
rect 40052 32842 40080 35866
rect 40960 35624 41012 35630
rect 40960 35566 41012 35572
rect 40132 35488 40184 35494
rect 40132 35430 40184 35436
rect 40144 35222 40172 35430
rect 40972 35290 41000 35566
rect 41156 35290 41184 37062
rect 41432 36378 41460 37062
rect 41616 36922 41644 37062
rect 41800 36922 41828 37062
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41788 36916 41840 36922
rect 41788 36858 41840 36864
rect 41420 36372 41472 36378
rect 41420 36314 41472 36320
rect 40960 35284 41012 35290
rect 40960 35226 41012 35232
rect 41144 35284 41196 35290
rect 41144 35226 41196 35232
rect 40132 35216 40184 35222
rect 40132 35158 40184 35164
rect 40868 35080 40920 35086
rect 40868 35022 40920 35028
rect 40880 34066 40908 35022
rect 42064 35012 42116 35018
rect 42064 34954 42116 34960
rect 42076 34746 42104 34954
rect 42168 34950 42196 38150
rect 42628 38010 42656 38286
rect 42616 38004 42668 38010
rect 42616 37946 42668 37952
rect 42248 37460 42300 37466
rect 42248 37402 42300 37408
rect 42260 36922 42288 37402
rect 42720 37210 42748 38354
rect 42984 38208 43036 38214
rect 42984 38150 43036 38156
rect 42996 38010 43024 38150
rect 42984 38004 43036 38010
rect 42984 37946 43036 37952
rect 43088 37890 43116 41482
rect 43168 40928 43220 40934
rect 43168 40870 43220 40876
rect 43260 40928 43312 40934
rect 43260 40870 43312 40876
rect 43180 40730 43208 40870
rect 43168 40724 43220 40730
rect 43168 40666 43220 40672
rect 43272 40526 43300 40870
rect 43364 40730 43392 41618
rect 43352 40724 43404 40730
rect 43352 40666 43404 40672
rect 43260 40520 43312 40526
rect 43260 40462 43312 40468
rect 43272 40050 43300 40462
rect 43260 40044 43312 40050
rect 43260 39986 43312 39992
rect 43272 38350 43300 39986
rect 43260 38344 43312 38350
rect 43260 38286 43312 38292
rect 42996 37862 43116 37890
rect 42996 37262 43024 37862
rect 43168 37800 43220 37806
rect 43168 37742 43220 37748
rect 42628 37194 42748 37210
rect 42984 37256 43036 37262
rect 42984 37198 43036 37204
rect 42616 37188 42748 37194
rect 42668 37182 42748 37188
rect 42616 37130 42668 37136
rect 42248 36916 42300 36922
rect 42248 36858 42300 36864
rect 42248 36780 42300 36786
rect 42248 36722 42300 36728
rect 42260 36038 42288 36722
rect 42628 36378 42656 37130
rect 42996 36854 43024 37198
rect 43180 37126 43208 37742
rect 43456 37346 43484 42842
rect 44180 42016 44232 42022
rect 44180 41958 44232 41964
rect 44088 41472 44140 41478
rect 44088 41414 44140 41420
rect 44100 40934 44128 41414
rect 44192 41138 44220 41958
rect 44180 41132 44232 41138
rect 44180 41074 44232 41080
rect 44088 40928 44140 40934
rect 44088 40870 44140 40876
rect 44180 39500 44232 39506
rect 44180 39442 44232 39448
rect 44192 39098 44220 39442
rect 44180 39092 44232 39098
rect 44180 39034 44232 39040
rect 44192 38026 44220 39034
rect 44192 37998 44312 38026
rect 43364 37318 43484 37346
rect 43168 37120 43220 37126
rect 43168 37062 43220 37068
rect 42984 36848 43036 36854
rect 42984 36790 43036 36796
rect 43076 36576 43128 36582
rect 43076 36518 43128 36524
rect 42616 36372 42668 36378
rect 42616 36314 42668 36320
rect 43088 36174 43116 36518
rect 43180 36378 43208 37062
rect 43168 36372 43220 36378
rect 43168 36314 43220 36320
rect 42708 36168 42760 36174
rect 42708 36110 42760 36116
rect 43076 36168 43128 36174
rect 43076 36110 43128 36116
rect 42248 36032 42300 36038
rect 42248 35974 42300 35980
rect 42260 35086 42288 35974
rect 42616 35488 42668 35494
rect 42616 35430 42668 35436
rect 42248 35080 42300 35086
rect 42248 35022 42300 35028
rect 42156 34944 42208 34950
rect 42156 34886 42208 34892
rect 42260 34746 42288 35022
rect 42064 34740 42116 34746
rect 42064 34682 42116 34688
rect 42248 34740 42300 34746
rect 42248 34682 42300 34688
rect 41420 34604 41472 34610
rect 41420 34546 41472 34552
rect 41432 34066 41460 34546
rect 40868 34060 40920 34066
rect 40868 34002 40920 34008
rect 41420 34060 41472 34066
rect 41420 34002 41472 34008
rect 40408 33856 40460 33862
rect 40408 33798 40460 33804
rect 40592 33856 40644 33862
rect 40592 33798 40644 33804
rect 40132 33448 40184 33454
rect 40132 33390 40184 33396
rect 40144 33114 40172 33390
rect 40132 33108 40184 33114
rect 40132 33050 40184 33056
rect 40420 33046 40448 33798
rect 40408 33040 40460 33046
rect 40408 32982 40460 32988
rect 40604 32910 40632 33798
rect 40880 33658 40908 34002
rect 42076 33998 42104 34682
rect 42628 34678 42656 35430
rect 42720 35154 42748 36110
rect 42708 35148 42760 35154
rect 42708 35090 42760 35096
rect 42720 34746 42748 35090
rect 43260 34944 43312 34950
rect 43260 34886 43312 34892
rect 42708 34740 42760 34746
rect 42708 34682 42760 34688
rect 42616 34672 42668 34678
rect 42616 34614 42668 34620
rect 42156 34604 42208 34610
rect 42156 34546 42208 34552
rect 42168 33998 42196 34546
rect 43272 33998 43300 34886
rect 42064 33992 42116 33998
rect 42064 33934 42116 33940
rect 42156 33992 42208 33998
rect 42156 33934 42208 33940
rect 43260 33992 43312 33998
rect 43260 33934 43312 33940
rect 42076 33658 42104 33934
rect 40868 33652 40920 33658
rect 40868 33594 40920 33600
rect 42064 33652 42116 33658
rect 42064 33594 42116 33600
rect 42524 33312 42576 33318
rect 42524 33254 42576 33260
rect 40592 32904 40644 32910
rect 40592 32846 40644 32852
rect 40040 32836 40092 32842
rect 40040 32778 40092 32784
rect 42432 32428 42484 32434
rect 42432 32370 42484 32376
rect 42248 32224 42300 32230
rect 42248 32166 42300 32172
rect 41052 31952 41104 31958
rect 41052 31894 41104 31900
rect 39672 31884 39724 31890
rect 39672 31826 39724 31832
rect 39764 31884 39816 31890
rect 39764 31826 39816 31832
rect 40040 31884 40092 31890
rect 40040 31826 40092 31832
rect 39684 31754 39712 31826
rect 39672 31748 39724 31754
rect 39672 31690 39724 31696
rect 39776 31686 39804 31826
rect 39764 31680 39816 31686
rect 39764 31622 39816 31628
rect 39764 31204 39816 31210
rect 39764 31146 39816 31152
rect 39776 30734 39804 31146
rect 40052 31142 40080 31826
rect 40776 31816 40828 31822
rect 40776 31758 40828 31764
rect 40684 31748 40736 31754
rect 40684 31690 40736 31696
rect 40696 31414 40724 31690
rect 40684 31408 40736 31414
rect 40684 31350 40736 31356
rect 40592 31272 40644 31278
rect 40592 31214 40644 31220
rect 40040 31136 40092 31142
rect 40040 31078 40092 31084
rect 40604 30938 40632 31214
rect 40592 30932 40644 30938
rect 40592 30874 40644 30880
rect 39488 30728 39540 30734
rect 39488 30670 39540 30676
rect 39764 30728 39816 30734
rect 39764 30670 39816 30676
rect 40500 30728 40552 30734
rect 40500 30670 40552 30676
rect 39776 30190 39804 30670
rect 40512 30394 40540 30670
rect 40500 30388 40552 30394
rect 40500 30330 40552 30336
rect 39764 30184 39816 30190
rect 39764 30126 39816 30132
rect 40592 30048 40644 30054
rect 40592 29990 40644 29996
rect 39856 29640 39908 29646
rect 39856 29582 39908 29588
rect 39580 27668 39632 27674
rect 39580 27610 39632 27616
rect 39592 25294 39620 27610
rect 39868 27606 39896 29582
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 39948 28960 40000 28966
rect 39948 28902 40000 28908
rect 39960 28558 39988 28902
rect 39948 28552 40000 28558
rect 39948 28494 40000 28500
rect 39856 27600 39908 27606
rect 39856 27542 39908 27548
rect 39856 27328 39908 27334
rect 39856 27270 39908 27276
rect 39868 27062 39896 27270
rect 39960 27062 39988 28494
rect 40512 28150 40540 29446
rect 40604 29306 40632 29990
rect 40696 29510 40724 31350
rect 40788 31142 40816 31758
rect 40776 31136 40828 31142
rect 40776 31078 40828 31084
rect 40788 30734 40816 31078
rect 41064 30938 41092 31894
rect 42156 31816 42208 31822
rect 42156 31758 42208 31764
rect 41144 31680 41196 31686
rect 41144 31622 41196 31628
rect 41052 30932 41104 30938
rect 41052 30874 41104 30880
rect 41156 30802 41184 31622
rect 42168 31482 42196 31758
rect 42156 31476 42208 31482
rect 42156 31418 42208 31424
rect 41328 30932 41380 30938
rect 41328 30874 41380 30880
rect 42156 30932 42208 30938
rect 42260 30920 42288 32166
rect 42444 31482 42472 32370
rect 42536 31890 42564 33254
rect 43364 32978 43392 37318
rect 44284 37262 44312 37998
rect 44272 37256 44324 37262
rect 44272 37198 44324 37204
rect 44284 36922 44312 37198
rect 44272 36916 44324 36922
rect 44272 36858 44324 36864
rect 43444 35080 43496 35086
rect 43444 35022 43496 35028
rect 43456 34202 43484 35022
rect 43720 34944 43772 34950
rect 43720 34886 43772 34892
rect 43732 34678 43760 34886
rect 43720 34672 43772 34678
rect 43720 34614 43772 34620
rect 44284 34610 44312 36858
rect 44272 34604 44324 34610
rect 44272 34546 44324 34552
rect 43444 34196 43496 34202
rect 43444 34138 43496 34144
rect 44638 34096 44694 34105
rect 44638 34031 44640 34040
rect 44692 34031 44694 34040
rect 44640 34002 44692 34008
rect 43904 33856 43956 33862
rect 43904 33798 43956 33804
rect 44088 33856 44140 33862
rect 44088 33798 44140 33804
rect 43916 33590 43944 33798
rect 43444 33584 43496 33590
rect 43444 33526 43496 33532
rect 43904 33584 43956 33590
rect 43904 33526 43956 33532
rect 43352 32972 43404 32978
rect 43352 32914 43404 32920
rect 43352 32224 43404 32230
rect 43352 32166 43404 32172
rect 42892 32020 42944 32026
rect 42892 31962 42944 31968
rect 42524 31884 42576 31890
rect 42524 31826 42576 31832
rect 42432 31476 42484 31482
rect 42432 31418 42484 31424
rect 42208 30892 42288 30920
rect 42156 30874 42208 30880
rect 41144 30796 41196 30802
rect 41144 30738 41196 30744
rect 40776 30728 40828 30734
rect 40776 30670 40828 30676
rect 41144 30184 41196 30190
rect 41144 30126 41196 30132
rect 41052 30048 41104 30054
rect 41052 29990 41104 29996
rect 40776 29640 40828 29646
rect 40776 29582 40828 29588
rect 40684 29504 40736 29510
rect 40684 29446 40736 29452
rect 40592 29300 40644 29306
rect 40592 29242 40644 29248
rect 40788 28626 40816 29582
rect 41064 29578 41092 29990
rect 41156 29850 41184 30126
rect 41236 30048 41288 30054
rect 41236 29990 41288 29996
rect 41144 29844 41196 29850
rect 41144 29786 41196 29792
rect 41248 29714 41276 29990
rect 41236 29708 41288 29714
rect 41236 29650 41288 29656
rect 41052 29572 41104 29578
rect 41052 29514 41104 29520
rect 40868 29096 40920 29102
rect 40868 29038 40920 29044
rect 40776 28620 40828 28626
rect 40776 28562 40828 28568
rect 40684 28484 40736 28490
rect 40684 28426 40736 28432
rect 40696 28218 40724 28426
rect 40684 28212 40736 28218
rect 40684 28154 40736 28160
rect 40500 28144 40552 28150
rect 40500 28086 40552 28092
rect 40880 28014 40908 29038
rect 40224 28008 40276 28014
rect 40224 27950 40276 27956
rect 40868 28008 40920 28014
rect 40868 27950 40920 27956
rect 40040 27872 40092 27878
rect 40040 27814 40092 27820
rect 39856 27056 39908 27062
rect 39856 26998 39908 27004
rect 39948 27056 40000 27062
rect 39948 26998 40000 27004
rect 40052 26314 40080 27814
rect 40132 26784 40184 26790
rect 40132 26726 40184 26732
rect 40144 26450 40172 26726
rect 40132 26444 40184 26450
rect 40132 26386 40184 26392
rect 40040 26308 40092 26314
rect 40040 26250 40092 26256
rect 39580 25288 39632 25294
rect 39580 25230 39632 25236
rect 39396 24404 39448 24410
rect 39396 24346 39448 24352
rect 40052 24274 40080 26250
rect 40132 25968 40184 25974
rect 40132 25910 40184 25916
rect 40144 25498 40172 25910
rect 40132 25492 40184 25498
rect 40132 25434 40184 25440
rect 40236 25294 40264 27950
rect 41064 27538 41092 29514
rect 41144 28484 41196 28490
rect 41144 28426 41196 28432
rect 41052 27532 41104 27538
rect 41052 27474 41104 27480
rect 40776 27464 40828 27470
rect 40776 27406 40828 27412
rect 40684 26920 40736 26926
rect 40684 26862 40736 26868
rect 40592 25696 40644 25702
rect 40592 25638 40644 25644
rect 40604 25294 40632 25638
rect 40696 25498 40724 26862
rect 40684 25492 40736 25498
rect 40684 25434 40736 25440
rect 40788 25294 40816 27406
rect 40960 26920 41012 26926
rect 40960 26862 41012 26868
rect 40972 26790 41000 26862
rect 40960 26784 41012 26790
rect 40960 26726 41012 26732
rect 40972 25498 41000 26726
rect 41156 26382 41184 28426
rect 41340 27402 41368 30874
rect 42536 30818 42564 31826
rect 42904 31482 42932 31962
rect 43364 31890 43392 32166
rect 43352 31884 43404 31890
rect 43352 31826 43404 31832
rect 43456 31754 43484 33526
rect 44100 33046 44128 33798
rect 44088 33040 44140 33046
rect 44088 32982 44140 32988
rect 43536 32972 43588 32978
rect 43536 32914 43588 32920
rect 43548 31754 43576 32914
rect 43812 32768 43864 32774
rect 43812 32710 43864 32716
rect 43824 32570 43852 32710
rect 43812 32564 43864 32570
rect 43812 32506 43864 32512
rect 44272 31884 44324 31890
rect 44272 31826 44324 31832
rect 44284 31754 44312 31826
rect 43444 31748 43496 31754
rect 43548 31726 43760 31754
rect 44284 31726 44404 31754
rect 43444 31690 43496 31696
rect 42892 31476 42944 31482
rect 42892 31418 42944 31424
rect 42800 31340 42852 31346
rect 42800 31282 42852 31288
rect 41984 30790 42564 30818
rect 42812 30802 42840 31282
rect 43168 31272 43220 31278
rect 43168 31214 43220 31220
rect 42800 30796 42852 30802
rect 41984 30734 42012 30790
rect 42800 30738 42852 30744
rect 41972 30728 42024 30734
rect 41972 30670 42024 30676
rect 41880 30592 41932 30598
rect 41880 30534 41932 30540
rect 41892 30258 41920 30534
rect 41880 30252 41932 30258
rect 41880 30194 41932 30200
rect 41984 28626 42012 30670
rect 43076 30592 43128 30598
rect 43076 30534 43128 30540
rect 43088 30394 43116 30534
rect 43076 30388 43128 30394
rect 43076 30330 43128 30336
rect 42524 30184 42576 30190
rect 42524 30126 42576 30132
rect 42536 29850 42564 30126
rect 42524 29844 42576 29850
rect 42524 29786 42576 29792
rect 43088 29714 43116 30330
rect 43180 30258 43208 31214
rect 43352 30796 43404 30802
rect 43352 30738 43404 30744
rect 43168 30252 43220 30258
rect 43168 30194 43220 30200
rect 43076 29708 43128 29714
rect 43076 29650 43128 29656
rect 42984 29572 43036 29578
rect 42984 29514 43036 29520
rect 42708 29504 42760 29510
rect 42708 29446 42760 29452
rect 42720 29306 42748 29446
rect 42708 29300 42760 29306
rect 42708 29242 42760 29248
rect 42800 29232 42852 29238
rect 42800 29174 42852 29180
rect 42432 28960 42484 28966
rect 42432 28902 42484 28908
rect 41972 28620 42024 28626
rect 41972 28562 42024 28568
rect 42444 28490 42472 28902
rect 42432 28484 42484 28490
rect 42432 28426 42484 28432
rect 42340 28416 42392 28422
rect 42340 28358 42392 28364
rect 41696 28008 41748 28014
rect 41696 27950 41748 27956
rect 41708 27606 41736 27950
rect 41696 27600 41748 27606
rect 41696 27542 41748 27548
rect 41328 27396 41380 27402
rect 41328 27338 41380 27344
rect 41236 27328 41288 27334
rect 41236 27270 41288 27276
rect 41248 26994 41276 27270
rect 41236 26988 41288 26994
rect 41236 26930 41288 26936
rect 41144 26376 41196 26382
rect 41144 26318 41196 26324
rect 41156 25974 41184 26318
rect 41144 25968 41196 25974
rect 41144 25910 41196 25916
rect 41052 25696 41104 25702
rect 41052 25638 41104 25644
rect 40960 25492 41012 25498
rect 40960 25434 41012 25440
rect 41064 25294 41092 25638
rect 40224 25288 40276 25294
rect 40224 25230 40276 25236
rect 40592 25288 40644 25294
rect 40592 25230 40644 25236
rect 40776 25288 40828 25294
rect 40776 25230 40828 25236
rect 41052 25288 41104 25294
rect 41052 25230 41104 25236
rect 40604 24954 40632 25230
rect 40592 24948 40644 24954
rect 40592 24890 40644 24896
rect 40132 24880 40184 24886
rect 40132 24822 40184 24828
rect 40040 24268 40092 24274
rect 40040 24210 40092 24216
rect 39396 23656 39448 23662
rect 39316 23604 39396 23610
rect 39316 23598 39448 23604
rect 39316 23582 39436 23598
rect 38752 22976 38804 22982
rect 38752 22918 38804 22924
rect 38764 22778 38792 22918
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38304 22066 38424 22094
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20466 38332 20878
rect 38292 20460 38344 20466
rect 38292 20402 38344 20408
rect 38304 20058 38332 20402
rect 38292 20052 38344 20058
rect 38292 19994 38344 20000
rect 38200 19168 38252 19174
rect 38200 19110 38252 19116
rect 38212 18902 38240 19110
rect 38200 18896 38252 18902
rect 38200 18838 38252 18844
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 38304 18426 38332 18770
rect 38292 18420 38344 18426
rect 38292 18362 38344 18368
rect 38108 15360 38160 15366
rect 38108 15302 38160 15308
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 38212 15094 38240 15302
rect 38200 15088 38252 15094
rect 38200 15030 38252 15036
rect 37188 14952 37240 14958
rect 37188 14894 37240 14900
rect 36084 14816 36136 14822
rect 36084 14758 36136 14764
rect 36820 14816 36872 14822
rect 36820 14758 36872 14764
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 36096 14414 36124 14758
rect 36832 14482 36860 14758
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 35440 14408 35492 14414
rect 35440 14350 35492 14356
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 35452 14074 35480 14350
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 32956 13796 33008 13802
rect 32956 13738 33008 13744
rect 32968 13530 32996 13738
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 32956 13524 33008 13530
rect 32956 13466 33008 13472
rect 33324 13184 33376 13190
rect 32876 13110 32996 13138
rect 33324 13126 33376 13132
rect 33968 13184 34020 13190
rect 33968 13126 34020 13132
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 32772 12980 32824 12986
rect 32824 12940 32904 12968
rect 32772 12922 32824 12928
rect 32680 12912 32732 12918
rect 32680 12854 32732 12860
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 32036 11348 32088 11354
rect 32036 11290 32088 11296
rect 32048 11150 32076 11290
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 31944 11008 31996 11014
rect 31944 10950 31996 10956
rect 31956 10810 31984 10950
rect 31944 10804 31996 10810
rect 31944 10746 31996 10752
rect 31956 10674 31984 10746
rect 31944 10668 31996 10674
rect 31944 10610 31996 10616
rect 32048 10606 32076 11086
rect 32036 10600 32088 10606
rect 32036 10542 32088 10548
rect 31944 10532 31996 10538
rect 31944 10474 31996 10480
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31772 9518 31800 9862
rect 31668 9512 31720 9518
rect 31668 9454 31720 9460
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31496 8362 31524 9114
rect 31588 9110 31616 9318
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31680 8974 31708 9454
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31484 8356 31536 8362
rect 31484 8298 31536 8304
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 31496 7886 31524 8298
rect 31576 8288 31628 8294
rect 31576 8230 31628 8236
rect 31588 8090 31616 8230
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31588 7342 31616 8026
rect 31772 7818 31800 9318
rect 31760 7812 31812 7818
rect 31760 7754 31812 7760
rect 31772 7478 31800 7754
rect 31864 7478 31892 10202
rect 31956 9382 31984 10474
rect 32048 9586 32076 10542
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 31944 9376 31996 9382
rect 31944 9318 31996 9324
rect 31944 8492 31996 8498
rect 31944 8434 31996 8440
rect 31956 8294 31984 8434
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31496 6798 31524 7142
rect 31484 6792 31536 6798
rect 31220 6718 31340 6746
rect 31484 6734 31536 6740
rect 31312 6662 31340 6718
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 31114 5536 31170 5545
rect 31114 5471 31170 5480
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30668 4826 30696 4966
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 30656 4820 30708 4826
rect 30656 4762 30708 4768
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 29196 4214 29224 4490
rect 29184 4208 29236 4214
rect 29184 4150 29236 4156
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27632 3058 27660 3538
rect 29196 3398 29224 4150
rect 30944 4078 30972 5170
rect 31128 5098 31156 5471
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31116 5092 31168 5098
rect 31116 5034 31168 5040
rect 31220 5080 31248 5170
rect 31576 5092 31628 5098
rect 31220 5052 31576 5080
rect 29460 4072 29512 4078
rect 29460 4014 29512 4020
rect 30932 4072 30984 4078
rect 30932 4014 30984 4020
rect 29472 3738 29500 4014
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 29184 3392 29236 3398
rect 29236 3340 29316 3346
rect 29184 3334 29316 3340
rect 29196 3318 29316 3334
rect 29288 3126 29316 3318
rect 31220 3194 31248 5052
rect 31576 5034 31628 5040
rect 31864 4282 31892 7414
rect 32140 5098 32168 12582
rect 32220 11620 32272 11626
rect 32220 11562 32272 11568
rect 32232 11150 32260 11562
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32220 10804 32272 10810
rect 32220 10746 32272 10752
rect 32232 9586 32260 10746
rect 32220 9580 32272 9586
rect 32220 9522 32272 9528
rect 32232 8634 32260 9522
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32324 5370 32352 12786
rect 32416 12714 32444 12786
rect 32692 12730 32720 12854
rect 32876 12782 32904 12940
rect 32968 12850 32996 13110
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 33232 12844 33284 12850
rect 33232 12786 33284 12792
rect 32864 12776 32916 12782
rect 32404 12708 32456 12714
rect 32692 12702 32812 12730
rect 32864 12718 32916 12724
rect 32404 12650 32456 12656
rect 32496 12640 32548 12646
rect 32496 12582 32548 12588
rect 32508 11082 32536 12582
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32600 11218 32628 11290
rect 32680 11280 32732 11286
rect 32784 11268 32812 12702
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32876 11354 32904 11630
rect 32968 11626 32996 12786
rect 32956 11620 33008 11626
rect 32956 11562 33008 11568
rect 32864 11348 32916 11354
rect 32864 11290 32916 11296
rect 32732 11240 32812 11268
rect 32680 11222 32732 11228
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 32508 10674 32536 11018
rect 32968 10674 32996 11562
rect 33244 11218 33272 12786
rect 33232 11212 33284 11218
rect 33232 11154 33284 11160
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32876 9654 32904 10406
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33152 7546 33180 8978
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 32864 6656 32916 6662
rect 32864 6598 32916 6604
rect 32876 5914 32904 6598
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 33152 5778 33180 7482
rect 32772 5772 32824 5778
rect 32772 5714 32824 5720
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 32312 5364 32364 5370
rect 32312 5306 32364 5312
rect 32784 5234 32812 5714
rect 33048 5568 33100 5574
rect 33048 5510 33100 5516
rect 32772 5228 32824 5234
rect 32772 5170 32824 5176
rect 32128 5092 32180 5098
rect 32128 5034 32180 5040
rect 32036 5024 32088 5030
rect 32036 4966 32088 4972
rect 32048 4690 32076 4966
rect 32784 4690 32812 5170
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 31852 4276 31904 4282
rect 31852 4218 31904 4224
rect 33060 4146 33088 5510
rect 33244 5302 33272 8298
rect 33336 5642 33364 13126
rect 33980 12238 34008 13126
rect 34348 12850 34376 13126
rect 34716 12850 34744 13670
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34704 12844 34756 12850
rect 34704 12786 34756 12792
rect 34808 12782 34836 13874
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35728 12850 35756 14350
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 35820 13530 35848 13874
rect 36084 13864 36136 13870
rect 36084 13806 36136 13812
rect 35900 13728 35952 13734
rect 35900 13670 35952 13676
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35912 12918 35940 13670
rect 36096 13394 36124 13806
rect 36832 13734 36860 14418
rect 36820 13728 36872 13734
rect 36820 13670 36872 13676
rect 37556 13524 37608 13530
rect 37556 13466 37608 13472
rect 36084 13388 36136 13394
rect 36084 13330 36136 13336
rect 36176 13388 36228 13394
rect 36176 13330 36228 13336
rect 35900 12912 35952 12918
rect 35900 12854 35952 12860
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 34796 12776 34848 12782
rect 34796 12718 34848 12724
rect 34808 12238 34836 12718
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35912 12434 35940 12854
rect 36096 12850 36124 13330
rect 36188 12986 36216 13330
rect 37568 13258 37596 13466
rect 38396 13258 38424 22066
rect 38764 21554 38792 22714
rect 39316 22574 39344 23582
rect 40144 23526 40172 24822
rect 40224 24200 40276 24206
rect 40224 24142 40276 24148
rect 40236 23866 40264 24142
rect 41064 23866 41092 25230
rect 41156 24070 41184 25910
rect 41248 25294 41276 26930
rect 41340 26926 41368 27338
rect 41328 26920 41380 26926
rect 41328 26862 41380 26868
rect 42156 26784 42208 26790
rect 42156 26726 42208 26732
rect 42168 26586 42196 26726
rect 42156 26580 42208 26586
rect 42156 26522 42208 26528
rect 42352 26450 42380 28358
rect 42524 28076 42576 28082
rect 42524 28018 42576 28024
rect 42536 27130 42564 28018
rect 42812 27538 42840 29174
rect 42892 29096 42944 29102
rect 42892 29038 42944 29044
rect 42904 28762 42932 29038
rect 42892 28756 42944 28762
rect 42892 28698 42944 28704
rect 42996 28490 43024 29514
rect 43180 29510 43208 30194
rect 43076 29504 43128 29510
rect 43076 29446 43128 29452
rect 43168 29504 43220 29510
rect 43168 29446 43220 29452
rect 43088 28626 43116 29446
rect 43076 28620 43128 28626
rect 43076 28562 43128 28568
rect 42984 28484 43036 28490
rect 42984 28426 43036 28432
rect 42800 27532 42852 27538
rect 42800 27474 42852 27480
rect 42800 27328 42852 27334
rect 42800 27270 42852 27276
rect 42892 27328 42944 27334
rect 42892 27270 42944 27276
rect 42524 27124 42576 27130
rect 42524 27066 42576 27072
rect 42812 26926 42840 27270
rect 42800 26920 42852 26926
rect 42800 26862 42852 26868
rect 42340 26444 42392 26450
rect 42340 26386 42392 26392
rect 41604 26240 41656 26246
rect 41604 26182 41656 26188
rect 41616 25906 41644 26182
rect 41604 25900 41656 25906
rect 41604 25842 41656 25848
rect 41236 25288 41288 25294
rect 41236 25230 41288 25236
rect 41144 24064 41196 24070
rect 41144 24006 41196 24012
rect 42248 24064 42300 24070
rect 42248 24006 42300 24012
rect 40224 23860 40276 23866
rect 40224 23802 40276 23808
rect 41052 23860 41104 23866
rect 41052 23802 41104 23808
rect 41156 23798 41184 24006
rect 42260 23866 42288 24006
rect 42812 23866 42840 26862
rect 42904 26858 42932 27270
rect 42892 26852 42944 26858
rect 42892 26794 42944 26800
rect 42904 26042 42932 26794
rect 43088 26058 43116 28562
rect 43180 27470 43208 29446
rect 43168 27464 43220 27470
rect 43168 27406 43220 27412
rect 42892 26036 42944 26042
rect 42892 25978 42944 25984
rect 42996 26030 43116 26058
rect 42892 25832 42944 25838
rect 42892 25774 42944 25780
rect 42248 23860 42300 23866
rect 42248 23802 42300 23808
rect 42800 23860 42852 23866
rect 42800 23802 42852 23808
rect 41144 23792 41196 23798
rect 41144 23734 41196 23740
rect 41512 23792 41564 23798
rect 41512 23734 41564 23740
rect 40132 23520 40184 23526
rect 40132 23462 40184 23468
rect 40144 22778 40172 23462
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 39304 22568 39356 22574
rect 39304 22510 39356 22516
rect 39856 22568 39908 22574
rect 39856 22510 39908 22516
rect 38844 22160 38896 22166
rect 38844 22102 38896 22108
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38856 21486 38884 22102
rect 39488 21888 39540 21894
rect 39488 21830 39540 21836
rect 39500 21554 39528 21830
rect 39488 21548 39540 21554
rect 39488 21490 39540 21496
rect 39580 21548 39632 21554
rect 39580 21490 39632 21496
rect 38844 21480 38896 21486
rect 38844 21422 38896 21428
rect 39304 21480 39356 21486
rect 39304 21422 39356 21428
rect 38568 21004 38620 21010
rect 38568 20946 38620 20952
rect 38580 19922 38608 20946
rect 38856 20942 38884 21422
rect 39120 21344 39172 21350
rect 39120 21286 39172 21292
rect 39028 21072 39080 21078
rect 39028 21014 39080 21020
rect 38844 20936 38896 20942
rect 38844 20878 38896 20884
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 38844 20256 38896 20262
rect 38844 20198 38896 20204
rect 38568 19916 38620 19922
rect 38568 19858 38620 19864
rect 38752 18692 38804 18698
rect 38752 18634 38804 18640
rect 38660 18624 38712 18630
rect 38660 18566 38712 18572
rect 38672 18426 38700 18566
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38764 17882 38792 18634
rect 38856 18426 38884 20198
rect 38948 20058 38976 20878
rect 39040 20466 39068 21014
rect 39132 20466 39160 21286
rect 39028 20460 39080 20466
rect 39028 20402 39080 20408
rect 39120 20460 39172 20466
rect 39120 20402 39172 20408
rect 38936 20052 38988 20058
rect 38936 19994 38988 20000
rect 38936 18896 38988 18902
rect 38936 18838 38988 18844
rect 38844 18420 38896 18426
rect 38844 18362 38896 18368
rect 38948 18170 38976 18838
rect 39316 18766 39344 21422
rect 39396 21344 39448 21350
rect 39396 21286 39448 21292
rect 39408 21010 39436 21286
rect 39592 21146 39620 21490
rect 39868 21418 39896 22510
rect 39948 22500 40000 22506
rect 39948 22442 40000 22448
rect 39960 21622 39988 22442
rect 40144 22098 40172 22714
rect 40408 22704 40460 22710
rect 40408 22646 40460 22652
rect 40224 22432 40276 22438
rect 40224 22374 40276 22380
rect 40132 22092 40184 22098
rect 40132 22034 40184 22040
rect 40236 22030 40264 22374
rect 40420 22234 40448 22646
rect 40960 22500 41012 22506
rect 40960 22442 41012 22448
rect 40408 22228 40460 22234
rect 40408 22170 40460 22176
rect 40500 22160 40552 22166
rect 40552 22108 40632 22114
rect 40500 22102 40632 22108
rect 40512 22086 40632 22102
rect 40972 22098 41000 22442
rect 41144 22432 41196 22438
rect 41144 22374 41196 22380
rect 41156 22098 41184 22374
rect 41236 22228 41288 22234
rect 41236 22170 41288 22176
rect 41248 22098 41276 22170
rect 40224 22024 40276 22030
rect 40224 21966 40276 21972
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 40224 21888 40276 21894
rect 40224 21830 40276 21836
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 39948 21616 40000 21622
rect 39948 21558 40000 21564
rect 39948 21480 40000 21486
rect 39948 21422 40000 21428
rect 39856 21412 39908 21418
rect 39856 21354 39908 21360
rect 39580 21140 39632 21146
rect 39580 21082 39632 21088
rect 39396 21004 39448 21010
rect 39396 20946 39448 20952
rect 39396 20800 39448 20806
rect 39592 20754 39620 21082
rect 39448 20748 39620 20754
rect 39396 20742 39620 20748
rect 39408 20726 39620 20742
rect 39396 19984 39448 19990
rect 39396 19926 39448 19932
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39304 18760 39356 18766
rect 39304 18702 39356 18708
rect 38856 18142 38976 18170
rect 39120 18148 39172 18154
rect 38752 17876 38804 17882
rect 38752 17818 38804 17824
rect 38764 17134 38792 17818
rect 38856 17338 38884 18142
rect 39120 18090 39172 18096
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 38844 17332 38896 17338
rect 38844 17274 38896 17280
rect 38752 17128 38804 17134
rect 38752 17070 38804 17076
rect 38856 16794 38884 17274
rect 38844 16788 38896 16794
rect 38844 16730 38896 16736
rect 38948 13394 38976 18022
rect 39028 17536 39080 17542
rect 39028 17478 39080 17484
rect 39040 16794 39068 17478
rect 39132 17338 39160 18090
rect 39224 17338 39252 18702
rect 39408 18442 39436 19926
rect 39488 19712 39540 19718
rect 39488 19654 39540 19660
rect 39500 19514 39528 19654
rect 39592 19514 39620 20726
rect 39868 20602 39896 21354
rect 39960 20942 39988 21422
rect 40052 21146 40080 21626
rect 40236 21554 40264 21830
rect 40132 21548 40184 21554
rect 40132 21490 40184 21496
rect 40224 21548 40276 21554
rect 40224 21490 40276 21496
rect 40040 21140 40092 21146
rect 40040 21082 40092 21088
rect 39948 20936 40000 20942
rect 39948 20878 40000 20884
rect 39856 20596 39908 20602
rect 39856 20538 39908 20544
rect 39764 20528 39816 20534
rect 39960 20482 39988 20878
rect 39816 20476 39988 20482
rect 39764 20470 39988 20476
rect 39776 20454 39988 20470
rect 40144 19854 40172 21490
rect 40236 21350 40264 21490
rect 40224 21344 40276 21350
rect 40224 21286 40276 21292
rect 40236 20806 40264 21286
rect 40328 20942 40356 21898
rect 40604 21554 40632 22086
rect 40960 22092 41012 22098
rect 40960 22034 41012 22040
rect 41144 22092 41196 22098
rect 41144 22034 41196 22040
rect 41236 22092 41288 22098
rect 41236 22034 41288 22040
rect 41524 22030 41552 23734
rect 42432 23520 42484 23526
rect 42432 23462 42484 23468
rect 41696 22432 41748 22438
rect 41696 22374 41748 22380
rect 41708 22030 41736 22374
rect 42156 22092 42208 22098
rect 42156 22034 42208 22040
rect 40776 22024 40828 22030
rect 40776 21966 40828 21972
rect 41328 22024 41380 22030
rect 41328 21966 41380 21972
rect 41512 22024 41564 22030
rect 41512 21966 41564 21972
rect 41696 22024 41748 22030
rect 41696 21966 41748 21972
rect 42064 22024 42116 22030
rect 42064 21966 42116 21972
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 40408 21344 40460 21350
rect 40408 21286 40460 21292
rect 40316 20936 40368 20942
rect 40316 20878 40368 20884
rect 40224 20800 40276 20806
rect 40224 20742 40276 20748
rect 40328 20602 40356 20878
rect 40316 20596 40368 20602
rect 40316 20538 40368 20544
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 39764 19780 39816 19786
rect 39764 19722 39816 19728
rect 39488 19508 39540 19514
rect 39488 19450 39540 19456
rect 39580 19508 39632 19514
rect 39580 19450 39632 19456
rect 39672 18624 39724 18630
rect 39672 18566 39724 18572
rect 39316 18414 39436 18442
rect 39684 18426 39712 18566
rect 39580 18420 39632 18426
rect 39120 17332 39172 17338
rect 39120 17274 39172 17280
rect 39212 17332 39264 17338
rect 39212 17274 39264 17280
rect 39028 16788 39080 16794
rect 39028 16730 39080 16736
rect 39120 15564 39172 15570
rect 39120 15506 39172 15512
rect 39028 13932 39080 13938
rect 39028 13874 39080 13880
rect 39040 13530 39068 13874
rect 39132 13530 39160 15506
rect 39316 15502 39344 18414
rect 39580 18362 39632 18368
rect 39672 18420 39724 18426
rect 39672 18362 39724 18368
rect 39592 18306 39620 18362
rect 39592 18290 39712 18306
rect 39396 18284 39448 18290
rect 39592 18284 39724 18290
rect 39592 18278 39672 18284
rect 39396 18226 39448 18232
rect 39672 18226 39724 18232
rect 39408 18154 39436 18226
rect 39776 18170 39804 19722
rect 40420 18834 40448 21286
rect 40788 21078 40816 21966
rect 40868 21888 40920 21894
rect 40868 21830 40920 21836
rect 41144 21888 41196 21894
rect 41144 21830 41196 21836
rect 40880 21690 40908 21830
rect 41156 21690 41184 21830
rect 40868 21684 40920 21690
rect 40868 21626 40920 21632
rect 41144 21684 41196 21690
rect 41144 21626 41196 21632
rect 41236 21412 41288 21418
rect 41236 21354 41288 21360
rect 40776 21072 40828 21078
rect 40776 21014 40828 21020
rect 41248 20874 41276 21354
rect 41340 21350 41368 21966
rect 41524 21690 41552 21966
rect 41512 21684 41564 21690
rect 41512 21626 41564 21632
rect 42076 21486 42104 21966
rect 41420 21480 41472 21486
rect 41420 21422 41472 21428
rect 41696 21480 41748 21486
rect 41696 21422 41748 21428
rect 42064 21480 42116 21486
rect 42064 21422 42116 21428
rect 41328 21344 41380 21350
rect 41328 21286 41380 21292
rect 41340 21146 41368 21286
rect 41328 21140 41380 21146
rect 41328 21082 41380 21088
rect 41432 21078 41460 21422
rect 41420 21072 41472 21078
rect 41420 21014 41472 21020
rect 41708 20942 41736 21422
rect 41972 21412 42024 21418
rect 41972 21354 42024 21360
rect 41696 20936 41748 20942
rect 41696 20878 41748 20884
rect 41236 20868 41288 20874
rect 41236 20810 41288 20816
rect 40408 18828 40460 18834
rect 40408 18770 40460 18776
rect 41984 18766 42012 21354
rect 42168 21146 42196 22034
rect 42340 21888 42392 21894
rect 42340 21830 42392 21836
rect 42156 21140 42208 21146
rect 42156 21082 42208 21088
rect 42168 20942 42196 21082
rect 42156 20936 42208 20942
rect 42156 20878 42208 20884
rect 42168 20602 42196 20878
rect 42248 20800 42300 20806
rect 42248 20742 42300 20748
rect 42156 20596 42208 20602
rect 42156 20538 42208 20544
rect 42260 20534 42288 20742
rect 42248 20528 42300 20534
rect 42248 20470 42300 20476
rect 42352 18970 42380 21830
rect 42444 21554 42472 23462
rect 42812 23118 42840 23802
rect 42904 23798 42932 25774
rect 42996 24410 43024 26030
rect 43076 25900 43128 25906
rect 43076 25842 43128 25848
rect 43088 25158 43116 25842
rect 43180 25838 43208 27406
rect 43260 27056 43312 27062
rect 43260 26998 43312 27004
rect 43272 26314 43300 26998
rect 43260 26308 43312 26314
rect 43260 26250 43312 26256
rect 43168 25832 43220 25838
rect 43168 25774 43220 25780
rect 43272 25226 43300 26250
rect 43260 25220 43312 25226
rect 43260 25162 43312 25168
rect 43076 25152 43128 25158
rect 43076 25094 43128 25100
rect 42984 24404 43036 24410
rect 42984 24346 43036 24352
rect 42892 23792 42944 23798
rect 42892 23734 42944 23740
rect 42996 23730 43024 24346
rect 42984 23724 43036 23730
rect 42984 23666 43036 23672
rect 43088 23526 43116 25094
rect 43364 24206 43392 30738
rect 43456 30734 43484 31690
rect 43444 30728 43496 30734
rect 43444 30670 43496 30676
rect 43444 25696 43496 25702
rect 43444 25638 43496 25644
rect 43456 25362 43484 25638
rect 43444 25356 43496 25362
rect 43444 25298 43496 25304
rect 43536 24268 43588 24274
rect 43536 24210 43588 24216
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 43168 24064 43220 24070
rect 43168 24006 43220 24012
rect 43076 23520 43128 23526
rect 43076 23462 43128 23468
rect 42800 23112 42852 23118
rect 43088 23066 43116 23462
rect 43180 23186 43208 24006
rect 43364 23798 43392 24142
rect 43352 23792 43404 23798
rect 43404 23752 43484 23780
rect 43352 23734 43404 23740
rect 43352 23656 43404 23662
rect 43352 23598 43404 23604
rect 43168 23180 43220 23186
rect 43168 23122 43220 23128
rect 43260 23112 43312 23118
rect 42852 23060 43024 23066
rect 42800 23054 43024 23060
rect 42812 23038 43024 23054
rect 43088 23038 43208 23066
rect 43260 23054 43312 23060
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 42812 22030 42840 22918
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42800 22024 42852 22030
rect 42800 21966 42852 21972
rect 42432 21548 42484 21554
rect 42432 21490 42484 21496
rect 42524 21548 42576 21554
rect 42524 21490 42576 21496
rect 42536 20942 42564 21490
rect 42628 21078 42656 21966
rect 42904 21554 42932 22102
rect 42996 21690 43024 23038
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 42984 21684 43036 21690
rect 42984 21626 43036 21632
rect 43088 21554 43116 22578
rect 43180 22574 43208 23038
rect 43272 22710 43300 23054
rect 43260 22704 43312 22710
rect 43260 22646 43312 22652
rect 43168 22568 43220 22574
rect 43168 22510 43220 22516
rect 43180 22030 43208 22510
rect 43364 22438 43392 23598
rect 43456 22642 43484 23752
rect 43548 23730 43576 24210
rect 43536 23724 43588 23730
rect 43588 23684 43668 23712
rect 43536 23666 43588 23672
rect 43444 22636 43496 22642
rect 43444 22578 43496 22584
rect 43352 22432 43404 22438
rect 43352 22374 43404 22380
rect 43364 22166 43392 22374
rect 43352 22160 43404 22166
rect 43352 22102 43404 22108
rect 43168 22024 43220 22030
rect 43168 21966 43220 21972
rect 42892 21548 42944 21554
rect 42892 21490 42944 21496
rect 43076 21548 43128 21554
rect 43076 21490 43128 21496
rect 42616 21072 42668 21078
rect 42616 21014 42668 21020
rect 42628 20942 42656 21014
rect 42904 21010 42932 21490
rect 42892 21004 42944 21010
rect 42892 20946 42944 20952
rect 43088 20942 43116 21490
rect 43168 21344 43220 21350
rect 43168 21286 43220 21292
rect 43260 21344 43312 21350
rect 43260 21286 43312 21292
rect 43180 21146 43208 21286
rect 43272 21146 43300 21286
rect 43168 21140 43220 21146
rect 43168 21082 43220 21088
rect 43260 21140 43312 21146
rect 43260 21082 43312 21088
rect 43364 20942 43392 22102
rect 43640 22030 43668 23684
rect 43536 22024 43588 22030
rect 43536 21966 43588 21972
rect 43628 22024 43680 22030
rect 43628 21966 43680 21972
rect 43548 21690 43576 21966
rect 43536 21684 43588 21690
rect 43536 21626 43588 21632
rect 43640 21554 43668 21966
rect 43444 21548 43496 21554
rect 43444 21490 43496 21496
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 42524 20936 42576 20942
rect 42524 20878 42576 20884
rect 42616 20936 42668 20942
rect 42616 20878 42668 20884
rect 43076 20936 43128 20942
rect 43076 20878 43128 20884
rect 43352 20936 43404 20942
rect 43352 20878 43404 20884
rect 42536 20602 42564 20878
rect 42892 20800 42944 20806
rect 42892 20742 42944 20748
rect 42984 20800 43036 20806
rect 42984 20742 43036 20748
rect 42524 20596 42576 20602
rect 42524 20538 42576 20544
rect 42800 20256 42852 20262
rect 42800 20198 42852 20204
rect 42524 19712 42576 19718
rect 42524 19654 42576 19660
rect 42536 19514 42564 19654
rect 42812 19514 42840 20198
rect 42524 19508 42576 19514
rect 42524 19450 42576 19456
rect 42800 19508 42852 19514
rect 42800 19450 42852 19456
rect 42904 19378 42932 20742
rect 42996 19854 43024 20742
rect 43456 20534 43484 21490
rect 43640 20942 43668 21490
rect 43628 20936 43680 20942
rect 43628 20878 43680 20884
rect 43444 20528 43496 20534
rect 43444 20470 43496 20476
rect 42984 19848 43036 19854
rect 42984 19790 43036 19796
rect 42996 19378 43024 19790
rect 43444 19780 43496 19786
rect 43444 19722 43496 19728
rect 43456 19378 43484 19722
rect 42708 19372 42760 19378
rect 42708 19314 42760 19320
rect 42892 19372 42944 19378
rect 42892 19314 42944 19320
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 43444 19372 43496 19378
rect 43444 19314 43496 19320
rect 43628 19372 43680 19378
rect 43628 19314 43680 19320
rect 42340 18964 42392 18970
rect 42340 18906 42392 18912
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41880 18760 41932 18766
rect 41880 18702 41932 18708
rect 41972 18760 42024 18766
rect 41972 18702 42024 18708
rect 40224 18692 40276 18698
rect 40224 18634 40276 18640
rect 39396 18148 39448 18154
rect 39396 18090 39448 18096
rect 39684 18142 39804 18170
rect 39580 18080 39632 18086
rect 39500 18040 39580 18068
rect 39396 17672 39448 17678
rect 39396 17614 39448 17620
rect 39408 17338 39436 17614
rect 39396 17332 39448 17338
rect 39396 17274 39448 17280
rect 39304 15496 39356 15502
rect 39304 15438 39356 15444
rect 39028 13524 39080 13530
rect 39028 13466 39080 13472
rect 39120 13524 39172 13530
rect 39120 13466 39172 13472
rect 38936 13388 38988 13394
rect 38936 13330 38988 13336
rect 36268 13252 36320 13258
rect 36268 13194 36320 13200
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 38384 13252 38436 13258
rect 38384 13194 38436 13200
rect 38568 13252 38620 13258
rect 38568 13194 38620 13200
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 36280 12782 36308 13194
rect 38580 12850 38608 13194
rect 38660 13184 38712 13190
rect 38660 13126 38712 13132
rect 38672 12968 38700 13126
rect 38856 12986 38884 13194
rect 38844 12980 38896 12986
rect 38672 12940 38792 12968
rect 38568 12844 38620 12850
rect 38568 12786 38620 12792
rect 36268 12776 36320 12782
rect 36268 12718 36320 12724
rect 37556 12776 37608 12782
rect 37556 12718 37608 12724
rect 35912 12406 36032 12434
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 35072 12232 35124 12238
rect 35072 12174 35124 12180
rect 33784 11212 33836 11218
rect 33784 11154 33836 11160
rect 33796 10742 33824 11154
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33508 10600 33560 10606
rect 33508 10542 33560 10548
rect 33520 9042 33548 10542
rect 33980 9450 34008 12174
rect 34532 11914 34560 12174
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34440 11898 34560 11914
rect 34428 11892 34560 11898
rect 34480 11886 34560 11892
rect 34612 11892 34664 11898
rect 34428 11834 34480 11840
rect 34612 11834 34664 11840
rect 34624 11082 34652 11834
rect 34704 11552 34756 11558
rect 34704 11494 34756 11500
rect 34716 11354 34744 11494
rect 34808 11354 34836 12038
rect 35084 11898 35112 12174
rect 35072 11892 35124 11898
rect 35072 11834 35124 11840
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11370 35388 11698
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34796 11348 34848 11354
rect 34796 11290 34848 11296
rect 35268 11342 35388 11370
rect 34612 11076 34664 11082
rect 34612 11018 34664 11024
rect 35072 11076 35124 11082
rect 35072 11018 35124 11024
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 33968 9444 34020 9450
rect 33968 9386 34020 9392
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 33508 9036 33560 9042
rect 33508 8978 33560 8984
rect 34072 8362 34100 9318
rect 34164 8634 34192 9318
rect 34808 8906 34836 10746
rect 35084 10674 35112 11018
rect 35268 10810 35296 11342
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 35256 10804 35308 10810
rect 35256 10746 35308 10752
rect 35072 10668 35124 10674
rect 35072 10610 35124 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 9042 35388 11154
rect 35532 10668 35584 10674
rect 35532 10610 35584 10616
rect 35348 9036 35400 9042
rect 35348 8978 35400 8984
rect 34796 8900 34848 8906
rect 34796 8842 34848 8848
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8634 34560 8774
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34348 7818 34376 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 34336 7812 34388 7818
rect 34336 7754 34388 7760
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33428 6866 33456 7686
rect 33796 7546 33824 7754
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 33324 5636 33376 5642
rect 33324 5578 33376 5584
rect 33232 5296 33284 5302
rect 33232 5238 33284 5244
rect 33336 5030 33364 5578
rect 33796 5302 33824 7482
rect 34348 6934 34376 7754
rect 35360 7750 35388 8978
rect 35440 8900 35492 8906
rect 35440 8842 35492 8848
rect 35452 8634 35480 8842
rect 35440 8628 35492 8634
rect 35440 8570 35492 8576
rect 35544 8430 35572 10610
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35348 7744 35400 7750
rect 35348 7686 35400 7692
rect 35360 7342 35388 7686
rect 35912 7478 35940 7754
rect 36004 7546 36032 12406
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 36096 10674 36124 12038
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 36188 10470 36216 11630
rect 36280 11150 36308 12718
rect 37568 11898 37596 12718
rect 38764 12434 38792 12940
rect 38844 12922 38896 12928
rect 39040 12850 39068 13466
rect 39132 13394 39160 13466
rect 39120 13388 39172 13394
rect 39120 13330 39172 13336
rect 39212 13388 39264 13394
rect 39212 13330 39264 13336
rect 39224 12986 39252 13330
rect 39304 13320 39356 13326
rect 39500 13274 39528 18040
rect 39580 18022 39632 18028
rect 39580 15496 39632 15502
rect 39580 15438 39632 15444
rect 39592 15162 39620 15438
rect 39580 15156 39632 15162
rect 39580 15098 39632 15104
rect 39580 13728 39632 13734
rect 39684 13716 39712 18142
rect 40236 17882 40264 18634
rect 40776 18624 40828 18630
rect 40776 18566 40828 18572
rect 40788 18426 40816 18566
rect 41248 18426 41276 18702
rect 41604 18624 41656 18630
rect 41604 18566 41656 18572
rect 40776 18420 40828 18426
rect 40776 18362 40828 18368
rect 41236 18420 41288 18426
rect 41236 18362 41288 18368
rect 41616 18290 41644 18566
rect 41892 18290 41920 18702
rect 41984 18290 42012 18702
rect 42352 18358 42380 18906
rect 42720 18902 42748 19314
rect 42904 18970 42932 19314
rect 42984 19168 43036 19174
rect 42984 19110 43036 19116
rect 42892 18964 42944 18970
rect 42892 18906 42944 18912
rect 42708 18896 42760 18902
rect 42708 18838 42760 18844
rect 42340 18352 42392 18358
rect 42340 18294 42392 18300
rect 41604 18284 41656 18290
rect 41604 18226 41656 18232
rect 41880 18284 41932 18290
rect 41880 18226 41932 18232
rect 41972 18284 42024 18290
rect 41972 18226 42024 18232
rect 40224 17876 40276 17882
rect 40224 17818 40276 17824
rect 40132 17604 40184 17610
rect 40132 17546 40184 17552
rect 39948 17536 40000 17542
rect 39948 17478 40000 17484
rect 39764 17196 39816 17202
rect 39764 17138 39816 17144
rect 39776 16046 39804 17138
rect 39960 16658 39988 17478
rect 40144 16794 40172 17546
rect 40236 17270 40264 17818
rect 40868 17536 40920 17542
rect 40868 17478 40920 17484
rect 40224 17264 40276 17270
rect 40224 17206 40276 17212
rect 40880 16794 40908 17478
rect 41616 17338 41644 18226
rect 41604 17332 41656 17338
rect 41604 17274 41656 17280
rect 41892 17134 41920 18226
rect 42720 17762 42748 18838
rect 42996 18766 43024 19110
rect 43352 18964 43404 18970
rect 43352 18906 43404 18912
rect 42984 18760 43036 18766
rect 42984 18702 43036 18708
rect 43076 18760 43128 18766
rect 43076 18702 43128 18708
rect 42800 18080 42852 18086
rect 42800 18022 42852 18028
rect 42812 17882 42840 18022
rect 42800 17876 42852 17882
rect 42800 17818 42852 17824
rect 42720 17746 42840 17762
rect 42340 17740 42392 17746
rect 42720 17740 42852 17746
rect 42720 17734 42800 17740
rect 42340 17682 42392 17688
rect 42800 17682 42852 17688
rect 42352 17626 42380 17682
rect 42524 17672 42576 17678
rect 42352 17598 42472 17626
rect 42524 17614 42576 17620
rect 42444 17542 42472 17598
rect 42156 17536 42208 17542
rect 42156 17478 42208 17484
rect 42432 17536 42484 17542
rect 42432 17478 42484 17484
rect 42168 17270 42196 17478
rect 42156 17264 42208 17270
rect 42156 17206 42208 17212
rect 41880 17128 41932 17134
rect 41880 17070 41932 17076
rect 41604 16992 41656 16998
rect 41604 16934 41656 16940
rect 42064 16992 42116 16998
rect 42064 16934 42116 16940
rect 42156 16992 42208 16998
rect 42156 16934 42208 16940
rect 40132 16788 40184 16794
rect 40132 16730 40184 16736
rect 40868 16788 40920 16794
rect 40868 16730 40920 16736
rect 39948 16652 40000 16658
rect 39948 16594 40000 16600
rect 39764 16040 39816 16046
rect 39764 15982 39816 15988
rect 39960 15570 39988 16594
rect 40500 16108 40552 16114
rect 40500 16050 40552 16056
rect 40224 15904 40276 15910
rect 40224 15846 40276 15852
rect 40236 15570 40264 15846
rect 39948 15564 40000 15570
rect 39948 15506 40000 15512
rect 40224 15564 40276 15570
rect 40224 15506 40276 15512
rect 39960 14618 39988 15506
rect 39948 14612 40000 14618
rect 39948 14554 40000 14560
rect 39960 14074 39988 14554
rect 39948 14068 40000 14074
rect 39948 14010 40000 14016
rect 40132 13864 40184 13870
rect 40132 13806 40184 13812
rect 39632 13688 39712 13716
rect 39580 13670 39632 13676
rect 39592 13326 39620 13670
rect 39304 13262 39356 13268
rect 39316 12986 39344 13262
rect 39408 13246 39528 13274
rect 39580 13320 39632 13326
rect 39580 13262 39632 13268
rect 39408 13190 39436 13246
rect 39396 13184 39448 13190
rect 39396 13126 39448 13132
rect 39488 13184 39540 13190
rect 39488 13126 39540 13132
rect 39500 12986 39528 13126
rect 39212 12980 39264 12986
rect 39212 12922 39264 12928
rect 39304 12980 39356 12986
rect 39304 12922 39356 12928
rect 39488 12980 39540 12986
rect 39488 12922 39540 12928
rect 39028 12844 39080 12850
rect 39028 12786 39080 12792
rect 39592 12714 39620 13262
rect 39672 13252 39724 13258
rect 39672 13194 39724 13200
rect 39580 12708 39632 12714
rect 39580 12650 39632 12656
rect 38672 12406 38792 12434
rect 38200 12300 38252 12306
rect 38200 12242 38252 12248
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 36452 11620 36504 11626
rect 36452 11562 36504 11568
rect 36464 11354 36492 11562
rect 36452 11348 36504 11354
rect 36452 11290 36504 11296
rect 37280 11212 37332 11218
rect 37280 11154 37332 11160
rect 36268 11144 36320 11150
rect 36268 11086 36320 11092
rect 36280 10810 36308 11086
rect 36544 11008 36596 11014
rect 36544 10950 36596 10956
rect 36268 10804 36320 10810
rect 36268 10746 36320 10752
rect 36556 10742 36584 10950
rect 37292 10810 37320 11154
rect 38212 11150 38240 12242
rect 38672 11830 38700 12406
rect 39684 12102 39712 13194
rect 40144 12986 40172 13806
rect 40132 12980 40184 12986
rect 40132 12922 40184 12928
rect 40512 12170 40540 16050
rect 40880 15434 40908 16730
rect 41512 16516 41564 16522
rect 41512 16458 41564 16464
rect 41524 15706 41552 16458
rect 41616 16046 41644 16934
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 41512 15700 41564 15706
rect 41512 15642 41564 15648
rect 41616 15502 41644 15982
rect 42076 15502 42104 16934
rect 42168 16046 42196 16934
rect 42444 16538 42472 17478
rect 42536 16658 42564 17614
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 42720 16794 42748 17070
rect 42708 16788 42760 16794
rect 42708 16730 42760 16736
rect 42524 16652 42576 16658
rect 42524 16594 42576 16600
rect 42260 16522 42472 16538
rect 42248 16516 42472 16522
rect 42300 16510 42472 16516
rect 42248 16458 42300 16464
rect 42156 16040 42208 16046
rect 42156 15982 42208 15988
rect 42168 15706 42196 15982
rect 42156 15700 42208 15706
rect 42156 15642 42208 15648
rect 41604 15496 41656 15502
rect 41604 15438 41656 15444
rect 42064 15496 42116 15502
rect 42064 15438 42116 15444
rect 40868 15428 40920 15434
rect 40868 15370 40920 15376
rect 42260 14346 42288 16458
rect 42536 16250 42564 16594
rect 42524 16244 42576 16250
rect 42524 16186 42576 16192
rect 42536 15570 42564 16186
rect 42524 15564 42576 15570
rect 42524 15506 42576 15512
rect 42800 15428 42852 15434
rect 42800 15370 42852 15376
rect 42812 14958 42840 15370
rect 43088 14958 43116 18702
rect 43364 18290 43392 18906
rect 43456 18630 43484 19314
rect 43640 18850 43668 19314
rect 43548 18822 43668 18850
rect 43444 18624 43496 18630
rect 43444 18566 43496 18572
rect 43352 18284 43404 18290
rect 43352 18226 43404 18232
rect 43456 16998 43484 18566
rect 43548 17338 43576 18822
rect 43628 18692 43680 18698
rect 43628 18634 43680 18640
rect 43640 18426 43668 18634
rect 43628 18420 43680 18426
rect 43628 18362 43680 18368
rect 43536 17332 43588 17338
rect 43536 17274 43588 17280
rect 43444 16992 43496 16998
rect 43444 16934 43496 16940
rect 43352 15428 43404 15434
rect 43352 15370 43404 15376
rect 43260 15020 43312 15026
rect 43260 14962 43312 14968
rect 42800 14952 42852 14958
rect 42800 14894 42852 14900
rect 43076 14952 43128 14958
rect 43076 14894 43128 14900
rect 41604 14340 41656 14346
rect 41604 14282 41656 14288
rect 42248 14340 42300 14346
rect 42248 14282 42300 14288
rect 41616 14074 41644 14282
rect 41604 14068 41656 14074
rect 41604 14010 41656 14016
rect 43088 13938 43116 14894
rect 43272 14618 43300 14962
rect 43364 14890 43392 15370
rect 43352 14884 43404 14890
rect 43352 14826 43404 14832
rect 43260 14612 43312 14618
rect 43260 14554 43312 14560
rect 43364 14074 43392 14826
rect 43548 14074 43576 17274
rect 43732 14482 43760 31726
rect 44272 27872 44324 27878
rect 44272 27814 44324 27820
rect 43812 27464 43864 27470
rect 43812 27406 43864 27412
rect 43824 26586 43852 27406
rect 43996 27328 44048 27334
rect 43996 27270 44048 27276
rect 44008 26926 44036 27270
rect 44284 26994 44312 27814
rect 44272 26988 44324 26994
rect 44272 26930 44324 26936
rect 43996 26920 44048 26926
rect 43996 26862 44048 26868
rect 43812 26580 43864 26586
rect 43812 26522 43864 26528
rect 44284 26450 44312 26930
rect 44272 26444 44324 26450
rect 44272 26386 44324 26392
rect 44284 25362 44312 26386
rect 44272 25356 44324 25362
rect 44272 25298 44324 25304
rect 44376 22098 44404 31726
rect 44638 25256 44694 25265
rect 44638 25191 44694 25200
rect 44652 24954 44680 25191
rect 44640 24948 44692 24954
rect 44640 24890 44692 24896
rect 44364 22092 44416 22098
rect 44364 22034 44416 22040
rect 43904 21888 43956 21894
rect 43904 21830 43956 21836
rect 43720 14476 43772 14482
rect 43720 14418 43772 14424
rect 43352 14068 43404 14074
rect 43352 14010 43404 14016
rect 43536 14068 43588 14074
rect 43536 14010 43588 14016
rect 43076 13932 43128 13938
rect 43076 13874 43128 13880
rect 40776 13864 40828 13870
rect 40776 13806 40828 13812
rect 40788 13530 40816 13806
rect 43260 13728 43312 13734
rect 43260 13670 43312 13676
rect 40776 13524 40828 13530
rect 40776 13466 40828 13472
rect 43272 13394 43300 13670
rect 43260 13388 43312 13394
rect 43260 13330 43312 13336
rect 43364 13258 43392 14010
rect 43352 13252 43404 13258
rect 43352 13194 43404 13200
rect 43732 12434 43760 14418
rect 43732 12406 43852 12434
rect 40500 12164 40552 12170
rect 40500 12106 40552 12112
rect 42524 12164 42576 12170
rect 42524 12106 42576 12112
rect 39028 12096 39080 12102
rect 39028 12038 39080 12044
rect 39672 12096 39724 12102
rect 39672 12038 39724 12044
rect 38660 11824 38712 11830
rect 38660 11766 38712 11772
rect 38476 11756 38528 11762
rect 38476 11698 38528 11704
rect 38488 11218 38516 11698
rect 38672 11218 38700 11766
rect 38936 11552 38988 11558
rect 38936 11494 38988 11500
rect 38948 11354 38976 11494
rect 38936 11348 38988 11354
rect 38936 11290 38988 11296
rect 38476 11212 38528 11218
rect 38476 11154 38528 11160
rect 38660 11212 38712 11218
rect 38660 11154 38712 11160
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 38200 11144 38252 11150
rect 38200 11086 38252 11092
rect 38568 11144 38620 11150
rect 38568 11086 38620 11092
rect 37372 11008 37424 11014
rect 37372 10950 37424 10956
rect 37384 10810 37412 10950
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 37372 10804 37424 10810
rect 37372 10746 37424 10752
rect 37660 10742 37688 11086
rect 36544 10736 36596 10742
rect 36544 10678 36596 10684
rect 37648 10736 37700 10742
rect 37648 10678 37700 10684
rect 37280 10668 37332 10674
rect 37332 10628 37412 10656
rect 37280 10610 37332 10616
rect 36912 10600 36964 10606
rect 36912 10542 36964 10548
rect 36176 10464 36228 10470
rect 36176 10406 36228 10412
rect 36924 9178 36952 10542
rect 37188 10532 37240 10538
rect 37240 10492 37320 10520
rect 37188 10474 37240 10480
rect 37292 10266 37320 10492
rect 37384 10470 37412 10628
rect 37372 10464 37424 10470
rect 37372 10406 37424 10412
rect 37280 10260 37332 10266
rect 37280 10202 37332 10208
rect 37660 10062 37688 10678
rect 38120 10266 38148 11086
rect 38580 10538 38608 11086
rect 38568 10532 38620 10538
rect 38568 10474 38620 10480
rect 38108 10260 38160 10266
rect 38108 10202 38160 10208
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 38580 9518 38608 10474
rect 39040 10470 39068 12038
rect 41420 11280 41472 11286
rect 41420 11222 41472 11228
rect 39488 11144 39540 11150
rect 39488 11086 39540 11092
rect 39500 10810 39528 11086
rect 39488 10804 39540 10810
rect 39488 10746 39540 10752
rect 41432 10606 41460 11222
rect 41420 10600 41472 10606
rect 41420 10542 41472 10548
rect 39028 10464 39080 10470
rect 39028 10406 39080 10412
rect 39040 10130 39068 10406
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 40868 9988 40920 9994
rect 40868 9930 40920 9936
rect 40880 9722 40908 9930
rect 40868 9716 40920 9722
rect 40868 9658 40920 9664
rect 42536 9654 42564 12106
rect 42800 11212 42852 11218
rect 42800 11154 42852 11160
rect 42524 9648 42576 9654
rect 42524 9590 42576 9596
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 41512 9512 41564 9518
rect 41512 9454 41564 9460
rect 36912 9172 36964 9178
rect 36912 9114 36964 9120
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 36084 8832 36136 8838
rect 36084 8774 36136 8780
rect 37740 8832 37792 8838
rect 37740 8774 37792 8780
rect 36096 8498 36124 8774
rect 37752 8634 37780 8774
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 37936 8294 37964 8910
rect 41524 8634 41552 9454
rect 41512 8628 41564 8634
rect 41512 8570 41564 8576
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 37924 8288 37976 8294
rect 37924 8230 37976 8236
rect 35992 7540 36044 7546
rect 35992 7482 36044 7488
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 36004 7290 36032 7482
rect 36188 7342 36216 8230
rect 37936 8022 37964 8230
rect 38028 8090 38056 8434
rect 38016 8084 38068 8090
rect 38016 8026 38068 8032
rect 37924 8016 37976 8022
rect 37924 7958 37976 7964
rect 37280 7948 37332 7954
rect 37280 7890 37332 7896
rect 37004 7744 37056 7750
rect 37056 7692 37136 7698
rect 37004 7686 37136 7692
rect 37016 7670 37136 7686
rect 36176 7336 36228 7342
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35256 6996 35308 7002
rect 35360 6984 35388 7278
rect 36004 7262 36124 7290
rect 36176 7278 36228 7284
rect 35308 6956 35388 6984
rect 35256 6938 35308 6944
rect 34336 6928 34388 6934
rect 34336 6870 34388 6876
rect 36096 6798 36124 7262
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 35072 6724 35124 6730
rect 35072 6666 35124 6672
rect 35084 6458 35112 6666
rect 35072 6452 35124 6458
rect 35072 6394 35124 6400
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34152 5568 34204 5574
rect 34152 5510 34204 5516
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33324 5024 33376 5030
rect 33324 4966 33376 4972
rect 34164 4622 34192 5510
rect 34612 5024 34664 5030
rect 34612 4966 34664 4972
rect 34624 4758 34652 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 34152 4616 34204 4622
rect 34152 4558 34204 4564
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34624 4282 34652 4558
rect 34612 4276 34664 4282
rect 34612 4218 34664 4224
rect 36096 4214 36124 6734
rect 37004 6656 37056 6662
rect 37004 6598 37056 6604
rect 37016 6254 37044 6598
rect 37004 6248 37056 6254
rect 37004 6190 37056 6196
rect 36084 4208 36136 4214
rect 36084 4150 36136 4156
rect 37108 4146 37136 7670
rect 37292 6798 37320 7890
rect 37372 7744 37424 7750
rect 37372 7686 37424 7692
rect 37384 7546 37412 7686
rect 37372 7540 37424 7546
rect 37372 7482 37424 7488
rect 37464 7540 37516 7546
rect 37464 7482 37516 7488
rect 37476 6866 37504 7482
rect 38212 6866 38240 8434
rect 38396 8090 38424 8434
rect 42812 8430 42840 11154
rect 43720 9376 43772 9382
rect 43720 9318 43772 9324
rect 43732 8566 43760 9318
rect 43720 8560 43772 8566
rect 43720 8502 43772 8508
rect 42800 8424 42852 8430
rect 42800 8366 42852 8372
rect 38384 8084 38436 8090
rect 38384 8026 38436 8032
rect 38568 7812 38620 7818
rect 38568 7754 38620 7760
rect 38580 7546 38608 7754
rect 42812 7546 42840 8366
rect 43352 7880 43404 7886
rect 43352 7822 43404 7828
rect 43364 7546 43392 7822
rect 38568 7540 38620 7546
rect 38568 7482 38620 7488
rect 42800 7540 42852 7546
rect 42800 7482 42852 7488
rect 43352 7540 43404 7546
rect 43352 7482 43404 7488
rect 38476 7472 38528 7478
rect 38476 7414 38528 7420
rect 38488 7342 38516 7414
rect 43732 7410 43760 8502
rect 43824 7478 43852 12406
rect 43916 11200 43944 21830
rect 44180 18216 44232 18222
rect 44180 18158 44232 18164
rect 44192 17746 44220 18158
rect 44180 17740 44232 17746
rect 44180 17682 44232 17688
rect 44192 17270 44220 17682
rect 44180 17264 44232 17270
rect 44180 17206 44232 17212
rect 44272 16992 44324 16998
rect 44272 16934 44324 16940
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 44008 15162 44036 16050
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44192 15745 44220 15846
rect 44178 15736 44234 15745
rect 44178 15671 44234 15680
rect 44284 15366 44312 16934
rect 44272 15360 44324 15366
rect 44272 15302 44324 15308
rect 43996 15156 44048 15162
rect 43996 15098 44048 15104
rect 44284 15026 44312 15302
rect 44272 15020 44324 15026
rect 44272 14962 44324 14968
rect 44088 13932 44140 13938
rect 44088 13874 44140 13880
rect 44100 13530 44128 13874
rect 44088 13524 44140 13530
rect 44088 13466 44140 13472
rect 43996 11212 44048 11218
rect 43916 11172 43996 11200
rect 43996 11154 44048 11160
rect 44272 11144 44324 11150
rect 44272 11086 44324 11092
rect 44284 9382 44312 11086
rect 44272 9376 44324 9382
rect 44272 9318 44324 9324
rect 43996 8424 44048 8430
rect 43996 8366 44048 8372
rect 44008 8090 44036 8366
rect 43996 8084 44048 8090
rect 43996 8026 44048 8032
rect 43812 7472 43864 7478
rect 43812 7414 43864 7420
rect 43720 7404 43772 7410
rect 43720 7346 43772 7352
rect 44088 7404 44140 7410
rect 44088 7346 44140 7352
rect 38476 7336 38528 7342
rect 38476 7278 38528 7284
rect 38936 7336 38988 7342
rect 38936 7278 38988 7284
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 38200 6860 38252 6866
rect 38200 6802 38252 6808
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 38212 6322 38240 6802
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38948 6254 38976 7278
rect 44100 6905 44128 7346
rect 44086 6896 44142 6905
rect 44086 6831 44142 6840
rect 38936 6248 38988 6254
rect 38936 6190 38988 6196
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 37096 4140 37148 4146
rect 37096 4082 37148 4088
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 29276 3120 29328 3126
rect 29276 3062 29328 3068
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 28828 2514 28856 2926
rect 28816 2508 28868 2514
rect 28816 2450 28868 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 32 800 60 2382
rect 8496 1306 8524 2382
rect 17512 1306 17540 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 8404 1278 8524 1306
rect 17420 1278 17540 1306
rect 8404 800 8432 1278
rect 17420 800 17448 1278
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 25778 0 25834 800
rect 25884 762 25912 870
rect 26160 762 26188 2382
rect 34808 800 34836 4082
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36832 3738 36860 4014
rect 36820 3732 36872 3738
rect 36820 3674 36872 3680
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36556 3194 36584 3470
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 43260 2916 43312 2922
rect 43260 2858 43312 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 43272 2650 43300 2858
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 43180 800 43208 2382
rect 25884 734 26188 762
rect 34794 0 34850 800
rect 43166 0 43222 800
<< via2 >>
rect 1398 45600 1454 45656
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 938 36760 994 36816
rect 938 27240 994 27296
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 938 18400 994 18456
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 10782 42744 10838 42800
rect 10506 30776 10562 30832
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 13910 42744 13966 42800
rect 11886 33516 11942 33552
rect 11886 33496 11888 33516
rect 11888 33496 11940 33516
rect 11940 33496 11942 33516
rect 12346 30640 12402 30696
rect 12990 30540 12992 30560
rect 12992 30540 13044 30560
rect 13044 30540 13046 30560
rect 12990 30504 13046 30540
rect 12990 30252 13046 30288
rect 12990 30232 12992 30252
rect 12992 30232 13044 30252
rect 13044 30232 13046 30252
rect 10782 16088 10838 16144
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4802 6332 4804 6352
rect 4804 6332 4856 6352
rect 4856 6332 4858 6352
rect 4802 6296 4858 6332
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 8206 6332 8208 6352
rect 8208 6332 8260 6352
rect 8260 6332 8262 6352
rect 8206 6296 8262 6332
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 10046 11892 10102 11928
rect 10046 11872 10048 11892
rect 10048 11872 10100 11892
rect 10100 11872 10102 11892
rect 9862 11212 9918 11248
rect 9862 11192 9864 11212
rect 9864 11192 9916 11212
rect 9916 11192 9918 11212
rect 10046 11328 10102 11384
rect 10414 10956 10416 10976
rect 10416 10956 10468 10976
rect 10468 10956 10470 10976
rect 10414 10920 10470 10956
rect 10874 11328 10930 11384
rect 10782 9036 10838 9072
rect 10782 9016 10784 9036
rect 10784 9016 10836 9036
rect 10836 9016 10838 9036
rect 10598 7112 10654 7168
rect 10506 6840 10562 6896
rect 10414 4256 10470 4312
rect 13450 33496 13506 33552
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 14462 42744 14518 42800
rect 13358 30232 13414 30288
rect 13910 30540 13912 30560
rect 13912 30540 13964 30560
rect 13964 30540 13966 30560
rect 13910 30504 13966 30540
rect 14094 30660 14150 30696
rect 14094 30640 14096 30660
rect 14096 30640 14148 30660
rect 14148 30640 14150 30660
rect 17222 32836 17278 32872
rect 17222 32816 17224 32836
rect 17224 32816 17276 32836
rect 17276 32816 17278 32836
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 17958 32816 18014 32872
rect 11794 13252 11850 13288
rect 11794 13232 11796 13252
rect 11796 13232 11848 13252
rect 11848 13232 11850 13252
rect 11886 12960 11942 13016
rect 11334 11464 11390 11520
rect 11334 11076 11390 11112
rect 11334 11056 11336 11076
rect 11336 11056 11388 11076
rect 11388 11056 11390 11076
rect 11518 9172 11574 9208
rect 11518 9152 11520 9172
rect 11520 9152 11572 9172
rect 11572 9152 11574 9172
rect 11518 8744 11574 8800
rect 11978 12688 12034 12744
rect 11702 9696 11758 9752
rect 11978 10240 12034 10296
rect 12162 9696 12218 9752
rect 11702 7112 11758 7168
rect 11426 4120 11482 4176
rect 11886 6432 11942 6488
rect 11886 5480 11942 5536
rect 11886 4936 11942 4992
rect 14094 13776 14150 13832
rect 12530 11328 12586 11384
rect 12622 10240 12678 10296
rect 12530 9016 12586 9072
rect 12254 6024 12310 6080
rect 13266 9580 13322 9616
rect 13266 9560 13268 9580
rect 13268 9560 13320 9580
rect 13320 9560 13322 9580
rect 13174 9288 13230 9344
rect 12254 3984 12310 4040
rect 8758 3068 8760 3088
rect 8760 3068 8812 3088
rect 8812 3068 8814 3088
rect 8758 3032 8814 3068
rect 13634 9424 13690 9480
rect 14094 12164 14150 12200
rect 14094 12144 14096 12164
rect 14096 12144 14148 12164
rect 14148 12144 14150 12164
rect 13910 10920 13966 10976
rect 13358 6160 13414 6216
rect 12898 4020 12900 4040
rect 12900 4020 12952 4040
rect 12952 4020 12954 4040
rect 12898 3984 12954 4020
rect 12254 3460 12310 3496
rect 12254 3440 12256 3460
rect 12256 3440 12308 3460
rect 12308 3440 12310 3460
rect 13266 3848 13322 3904
rect 14186 9424 14242 9480
rect 13910 8880 13966 8936
rect 14186 8744 14242 8800
rect 13542 5888 13598 5944
rect 13726 6060 13728 6080
rect 13728 6060 13780 6080
rect 13780 6060 13782 6080
rect 13726 6024 13782 6060
rect 13542 5652 13544 5672
rect 13544 5652 13596 5672
rect 13596 5652 13598 5672
rect 13542 5616 13598 5652
rect 13910 5480 13966 5536
rect 13818 3848 13874 3904
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 20074 31628 20076 31648
rect 20076 31628 20128 31648
rect 20128 31628 20130 31648
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19246 30640 19302 30696
rect 19890 30912 19946 30968
rect 19798 30776 19854 30832
rect 20074 31592 20130 31628
rect 20166 30776 20222 30832
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19338 30252 19394 30288
rect 19338 30232 19340 30252
rect 19340 30232 19392 30252
rect 19392 30232 19394 30252
rect 19798 30096 19854 30152
rect 20258 30540 20260 30560
rect 20260 30540 20312 30560
rect 20312 30540 20314 30560
rect 20258 30504 20314 30540
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20994 31628 20996 31648
rect 20996 31628 21048 31648
rect 21048 31628 21050 31648
rect 20994 31592 21050 31628
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 21086 30932 21142 30968
rect 21086 30912 21088 30932
rect 21088 30912 21140 30932
rect 21140 30912 21142 30932
rect 20902 30640 20958 30696
rect 21546 30368 21602 30424
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19522 23044 19578 23080
rect 19522 23024 19524 23044
rect 19524 23024 19576 23044
rect 19576 23024 19578 23044
rect 19338 22888 19394 22944
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19890 22616 19946 22672
rect 19706 22500 19762 22536
rect 19706 22480 19708 22500
rect 19708 22480 19760 22500
rect 19760 22480 19762 22500
rect 19430 22344 19486 22400
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 16302 16088 16358 16144
rect 16486 14476 16542 14512
rect 16486 14456 16488 14476
rect 16488 14456 16540 14476
rect 16540 14456 16542 14476
rect 14738 12844 14794 12880
rect 14738 12824 14740 12844
rect 14740 12824 14792 12844
rect 14792 12824 14794 12844
rect 15382 12552 15438 12608
rect 14922 11872 14978 11928
rect 14554 11056 14610 11112
rect 15198 11192 15254 11248
rect 14646 9596 14648 9616
rect 14648 9596 14700 9616
rect 14700 9596 14702 9616
rect 14646 9560 14702 9596
rect 15658 12144 15714 12200
rect 15842 9460 15844 9480
rect 15844 9460 15896 9480
rect 15896 9460 15898 9480
rect 15842 9424 15898 9460
rect 15290 9288 15346 9344
rect 14922 8916 14924 8936
rect 14924 8916 14976 8936
rect 14976 8916 14978 8936
rect 14922 8880 14978 8916
rect 14922 6296 14978 6352
rect 15106 6432 15162 6488
rect 15014 5344 15070 5400
rect 15566 6160 15622 6216
rect 17406 12688 17462 12744
rect 16486 9460 16488 9480
rect 16488 9460 16540 9480
rect 16540 9460 16542 9480
rect 16486 9424 16542 9460
rect 15750 6568 15806 6624
rect 15566 4392 15622 4448
rect 14922 4276 14978 4312
rect 14922 4256 14924 4276
rect 14924 4256 14976 4276
rect 14976 4256 14978 4276
rect 14830 3476 14832 3496
rect 14832 3476 14884 3496
rect 14884 3476 14886 3496
rect 14830 3440 14886 3476
rect 16486 4392 16542 4448
rect 17314 9696 17370 9752
rect 17590 9052 17592 9072
rect 17592 9052 17644 9072
rect 17644 9052 17646 9072
rect 17590 9016 17646 9052
rect 16762 5480 16818 5536
rect 17130 6024 17186 6080
rect 17314 6432 17370 6488
rect 17590 6316 17646 6352
rect 17590 6296 17592 6316
rect 17592 6296 17644 6316
rect 17644 6296 17646 6316
rect 17130 5344 17186 5400
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20166 23024 20222 23080
rect 19890 19388 19892 19408
rect 19892 19388 19944 19408
rect 19944 19388 19946 19408
rect 18602 14456 18658 14512
rect 18234 12960 18290 13016
rect 18050 11056 18106 11112
rect 18234 9052 18236 9072
rect 18236 9052 18288 9072
rect 18288 9052 18290 9072
rect 18234 9016 18290 9052
rect 18050 6160 18106 6216
rect 17866 6024 17922 6080
rect 17498 5616 17554 5672
rect 16946 3884 16948 3904
rect 16948 3884 17000 3904
rect 17000 3884 17002 3904
rect 16946 3848 17002 3884
rect 17866 4392 17922 4448
rect 17590 4120 17646 4176
rect 19890 19352 19946 19388
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 18786 9696 18842 9752
rect 18878 9016 18934 9072
rect 18142 5480 18198 5536
rect 18234 4936 18290 4992
rect 18326 4140 18382 4176
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19522 11464 19578 11520
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 5908 19394 5944
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19338 5888 19340 5908
rect 19340 5888 19392 5908
rect 19392 5888 19394 5908
rect 19338 5616 19394 5672
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 18326 4120 18328 4140
rect 18328 4120 18380 4140
rect 18380 4120 18382 4140
rect 18142 3984 18198 4040
rect 19062 4120 19118 4176
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21546 15408 21602 15464
rect 21270 11092 21272 11112
rect 21272 11092 21324 11112
rect 21324 11092 21326 11112
rect 21270 11056 21326 11092
rect 22006 13232 22062 13288
rect 22006 12960 22062 13016
rect 22098 12280 22154 12336
rect 22098 10920 22154 10976
rect 22098 10668 22154 10704
rect 22098 10648 22100 10668
rect 22100 10648 22152 10668
rect 22152 10648 22154 10668
rect 22466 12960 22522 13016
rect 23386 22344 23442 22400
rect 23846 22480 23902 22536
rect 23202 15428 23258 15464
rect 23202 15408 23204 15428
rect 23204 15408 23256 15428
rect 23256 15408 23258 15428
rect 23386 13096 23442 13152
rect 22558 10920 22614 10976
rect 23018 10648 23074 10704
rect 25502 20576 25558 20632
rect 25778 20032 25834 20088
rect 25502 19372 25558 19408
rect 25502 19352 25504 19372
rect 25504 19352 25556 19372
rect 25556 19352 25558 19372
rect 25502 12980 25558 13016
rect 25502 12960 25504 12980
rect 25504 12960 25556 12980
rect 25556 12960 25558 12980
rect 24950 12824 25006 12880
rect 26146 12824 26202 12880
rect 25318 7248 25374 7304
rect 18694 3052 18750 3088
rect 18694 3032 18696 3052
rect 18696 3032 18748 3052
rect 18748 3032 18750 3052
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 22926 4120 22982 4176
rect 28078 30368 28134 30424
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 28262 19760 28318 19816
rect 29826 22636 29882 22672
rect 29826 22616 29828 22636
rect 29828 22616 29880 22636
rect 29880 22616 29882 22636
rect 29826 20324 29882 20360
rect 29826 20304 29828 20324
rect 29828 20304 29880 20324
rect 29880 20304 29882 20324
rect 30562 20576 30618 20632
rect 30378 19760 30434 19816
rect 30286 16108 30342 16144
rect 30286 16088 30288 16108
rect 30288 16088 30340 16108
rect 30340 16088 30342 16108
rect 30838 15988 30840 16008
rect 30840 15988 30892 16008
rect 30892 15988 30894 16008
rect 30838 15952 30894 15988
rect 31206 28192 31262 28248
rect 31390 28484 31446 28520
rect 31390 28464 31392 28484
rect 31392 28464 31444 28484
rect 31444 28464 31446 28484
rect 31298 20304 31354 20360
rect 31206 20032 31262 20088
rect 31298 15952 31354 16008
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 32310 28212 32366 28248
rect 32310 28192 32312 28212
rect 32312 28192 32364 28212
rect 32364 28192 32366 28212
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 32218 16108 32274 16144
rect 32218 16088 32220 16108
rect 32220 16088 32272 16108
rect 32272 16088 32274 16108
rect 31850 15972 31906 16008
rect 26974 13096 27030 13152
rect 27618 11056 27674 11112
rect 26790 7248 26846 7304
rect 24490 4120 24546 4176
rect 28722 7420 28724 7440
rect 28724 7420 28776 7440
rect 28776 7420 28778 7440
rect 28722 7384 28778 7420
rect 29458 7420 29460 7440
rect 29460 7420 29512 7440
rect 29512 7420 29514 7440
rect 29458 7384 29514 7420
rect 31850 15952 31852 15972
rect 31852 15952 31904 15972
rect 31904 15952 31906 15972
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34518 28464 34574 28520
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34150 22616 34206 22672
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 31482 12824 31538 12880
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 44638 43560 44694 43616
rect 40314 41540 40370 41576
rect 40314 41520 40316 41540
rect 40316 41520 40368 41540
rect 40368 41520 40370 41540
rect 41602 41520 41658 41576
rect 44638 34060 44694 34096
rect 44638 34040 44640 34060
rect 44640 34040 44692 34060
rect 44692 34040 44694 34060
rect 31114 5480 31170 5536
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 44638 25200 44694 25256
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 44178 15680 44234 15736
rect 44086 6840 44142 6896
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 19570 45728 19886 45729
rect 0 45658 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 1393 45658 1459 45661
rect 0 45656 1459 45658
rect 0 45600 1398 45656
rect 1454 45600 1459 45656
rect 0 45598 1459 45600
rect 0 45568 800 45598
rect 1393 45595 1459 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 44633 43618 44699 43621
rect 44933 43618 45733 43648
rect 44633 43616 45733 43618
rect 44633 43560 44638 43616
rect 44694 43560 45733 43616
rect 44633 43558 45733 43560
rect 44633 43555 44699 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 44933 43528 45733 43558
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 10777 42802 10843 42805
rect 13905 42802 13971 42805
rect 14457 42802 14523 42805
rect 10777 42800 14523 42802
rect 10777 42744 10782 42800
rect 10838 42744 13910 42800
rect 13966 42744 14462 42800
rect 14518 42744 14523 42800
rect 10777 42742 14523 42744
rect 10777 42739 10843 42742
rect 13905 42739 13971 42742
rect 14457 42739 14523 42742
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 40309 41578 40375 41581
rect 41597 41578 41663 41581
rect 40309 41576 41663 41578
rect 40309 41520 40314 41576
rect 40370 41520 41602 41576
rect 41658 41520 41663 41576
rect 40309 41518 41663 41520
rect 40309 41515 40375 41518
rect 41597 41515 41663 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 44633 34098 44699 34101
rect 44933 34098 45733 34128
rect 44633 34096 45733 34098
rect 44633 34040 44638 34096
rect 44694 34040 45733 34096
rect 44633 34038 45733 34040
rect 44633 34035 44699 34038
rect 44933 34008 45733 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 11881 33554 11947 33557
rect 13445 33554 13511 33557
rect 11881 33552 13511 33554
rect 11881 33496 11886 33552
rect 11942 33496 13450 33552
rect 13506 33496 13511 33552
rect 11881 33494 13511 33496
rect 11881 33491 11947 33494
rect 13445 33491 13511 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 17217 32874 17283 32877
rect 17953 32874 18019 32877
rect 17217 32872 18019 32874
rect 17217 32816 17222 32872
rect 17278 32816 17958 32872
rect 18014 32816 18019 32872
rect 17217 32814 18019 32816
rect 17217 32811 17283 32814
rect 17953 32811 18019 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 20069 31650 20135 31653
rect 20989 31650 21055 31653
rect 20069 31648 21055 31650
rect 20069 31592 20074 31648
rect 20130 31592 20994 31648
rect 21050 31592 21055 31648
rect 20069 31590 21055 31592
rect 20069 31587 20135 31590
rect 20989 31587 21055 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19885 30970 19951 30973
rect 21081 30970 21147 30973
rect 19885 30968 21147 30970
rect 19885 30912 19890 30968
rect 19946 30912 21086 30968
rect 21142 30912 21147 30968
rect 19885 30910 21147 30912
rect 19885 30907 19951 30910
rect 21081 30907 21147 30910
rect 10501 30834 10567 30837
rect 19793 30834 19859 30837
rect 20161 30836 20227 30837
rect 20110 30834 20116 30836
rect 10501 30832 19859 30834
rect 10501 30776 10506 30832
rect 10562 30776 19798 30832
rect 19854 30776 19859 30832
rect 10501 30774 19859 30776
rect 20070 30774 20116 30834
rect 20180 30832 20227 30836
rect 20222 30776 20227 30832
rect 10501 30771 10567 30774
rect 19793 30771 19859 30774
rect 20110 30772 20116 30774
rect 20180 30772 20227 30776
rect 20161 30771 20227 30772
rect 12341 30698 12407 30701
rect 14089 30698 14155 30701
rect 12341 30696 14155 30698
rect 12341 30640 12346 30696
rect 12402 30640 14094 30696
rect 14150 30640 14155 30696
rect 12341 30638 14155 30640
rect 12341 30635 12407 30638
rect 14089 30635 14155 30638
rect 19241 30698 19307 30701
rect 20897 30698 20963 30701
rect 19241 30696 20963 30698
rect 19241 30640 19246 30696
rect 19302 30640 20902 30696
rect 20958 30640 20963 30696
rect 19241 30638 20963 30640
rect 19241 30635 19307 30638
rect 20897 30635 20963 30638
rect 12985 30562 13051 30565
rect 13905 30562 13971 30565
rect 12985 30560 13971 30562
rect 12985 30504 12990 30560
rect 13046 30504 13910 30560
rect 13966 30504 13971 30560
rect 12985 30502 13971 30504
rect 12985 30499 13051 30502
rect 13905 30499 13971 30502
rect 20253 30562 20319 30565
rect 20253 30560 20914 30562
rect 20253 30504 20258 30560
rect 20314 30504 20914 30560
rect 20253 30502 20914 30504
rect 20253 30499 20319 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 12985 30290 13051 30293
rect 13353 30290 13419 30293
rect 12985 30288 13419 30290
rect 12985 30232 12990 30288
rect 13046 30232 13358 30288
rect 13414 30232 13419 30288
rect 12985 30230 13419 30232
rect 12985 30227 13051 30230
rect 13353 30227 13419 30230
rect 19333 30290 19399 30293
rect 20854 30290 20914 30502
rect 21541 30426 21607 30429
rect 28073 30426 28139 30429
rect 21541 30424 28139 30426
rect 21541 30368 21546 30424
rect 21602 30368 28078 30424
rect 28134 30368 28139 30424
rect 21541 30366 28139 30368
rect 21541 30363 21607 30366
rect 28073 30363 28139 30366
rect 19333 30288 20914 30290
rect 19333 30232 19338 30288
rect 19394 30232 20914 30288
rect 19333 30230 20914 30232
rect 19333 30227 19399 30230
rect 19793 30154 19859 30157
rect 20110 30154 20116 30156
rect 19793 30152 20116 30154
rect 19793 30096 19798 30152
rect 19854 30096 20116 30152
rect 19793 30094 20116 30096
rect 19793 30091 19859 30094
rect 20110 30092 20116 30094
rect 20180 30092 20186 30156
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 31385 28522 31451 28525
rect 34513 28522 34579 28525
rect 31385 28520 34579 28522
rect 31385 28464 31390 28520
rect 31446 28464 34518 28520
rect 34574 28464 34579 28520
rect 31385 28462 34579 28464
rect 31385 28459 31451 28462
rect 34513 28459 34579 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 31201 28250 31267 28253
rect 32305 28250 32371 28253
rect 31201 28248 32371 28250
rect 31201 28192 31206 28248
rect 31262 28192 32310 28248
rect 32366 28192 32371 28248
rect 31201 28190 32371 28192
rect 31201 28187 31267 28190
rect 32305 28187 32371 28190
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27298 800 27328
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 0 27208 800 27238
rect 933 27235 999 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 44633 25258 44699 25261
rect 44933 25258 45733 25288
rect 44633 25256 45733 25258
rect 44633 25200 44638 25256
rect 44694 25200 45733 25256
rect 44633 25198 45733 25200
rect 44633 25195 44699 25198
rect 44933 25168 45733 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19517 23082 19583 23085
rect 20161 23082 20227 23085
rect 19517 23080 20227 23082
rect 19517 23024 19522 23080
rect 19578 23024 20166 23080
rect 20222 23024 20227 23080
rect 19517 23022 20227 23024
rect 19517 23019 19583 23022
rect 20161 23019 20227 23022
rect 19333 22946 19399 22949
rect 19333 22944 19442 22946
rect 19333 22888 19338 22944
rect 19394 22888 19442 22944
rect 19333 22883 19442 22888
rect 19382 22674 19442 22883
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 19885 22674 19951 22677
rect 19382 22672 19951 22674
rect 19382 22616 19890 22672
rect 19946 22616 19951 22672
rect 19382 22614 19951 22616
rect 19885 22611 19951 22614
rect 29821 22674 29887 22677
rect 34145 22674 34211 22677
rect 29821 22672 34211 22674
rect 29821 22616 29826 22672
rect 29882 22616 34150 22672
rect 34206 22616 34211 22672
rect 29821 22614 34211 22616
rect 29821 22611 29887 22614
rect 34145 22611 34211 22614
rect 19701 22538 19767 22541
rect 23841 22538 23907 22541
rect 19701 22536 23907 22538
rect 19701 22480 19706 22536
rect 19762 22480 23846 22536
rect 23902 22480 23907 22536
rect 19701 22478 23907 22480
rect 19701 22475 19767 22478
rect 23841 22475 23907 22478
rect 19425 22402 19491 22405
rect 23381 22402 23447 22405
rect 19425 22400 23447 22402
rect 19425 22344 19430 22400
rect 19486 22344 23386 22400
rect 23442 22344 23447 22400
rect 19425 22342 23447 22344
rect 19425 22339 19491 22342
rect 23381 22339 23447 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 25497 20634 25563 20637
rect 30557 20634 30623 20637
rect 25497 20632 30623 20634
rect 25497 20576 25502 20632
rect 25558 20576 30562 20632
rect 30618 20576 30623 20632
rect 25497 20574 30623 20576
rect 25497 20571 25563 20574
rect 30557 20571 30623 20574
rect 29821 20362 29887 20365
rect 31293 20362 31359 20365
rect 29821 20360 31359 20362
rect 29821 20304 29826 20360
rect 29882 20304 31298 20360
rect 31354 20304 31359 20360
rect 29821 20302 31359 20304
rect 29821 20299 29887 20302
rect 31293 20299 31359 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 25773 20090 25839 20093
rect 31201 20090 31267 20093
rect 25773 20088 31267 20090
rect 25773 20032 25778 20088
rect 25834 20032 31206 20088
rect 31262 20032 31267 20088
rect 25773 20030 31267 20032
rect 25773 20027 25839 20030
rect 31201 20027 31267 20030
rect 28257 19818 28323 19821
rect 30373 19818 30439 19821
rect 28257 19816 30439 19818
rect 28257 19760 28262 19816
rect 28318 19760 30378 19816
rect 30434 19760 30439 19816
rect 28257 19758 30439 19760
rect 28257 19755 28323 19758
rect 30373 19755 30439 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 19885 19410 19951 19413
rect 25497 19410 25563 19413
rect 19885 19408 25563 19410
rect 19885 19352 19890 19408
rect 19946 19352 25502 19408
rect 25558 19352 25563 19408
rect 19885 19350 25563 19352
rect 19885 19347 19951 19350
rect 25497 19347 25563 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 10777 16146 10843 16149
rect 16297 16146 16363 16149
rect 10777 16144 16363 16146
rect 10777 16088 10782 16144
rect 10838 16088 16302 16144
rect 16358 16088 16363 16144
rect 10777 16086 16363 16088
rect 10777 16083 10843 16086
rect 16297 16083 16363 16086
rect 30281 16146 30347 16149
rect 32213 16146 32279 16149
rect 30281 16144 32279 16146
rect 30281 16088 30286 16144
rect 30342 16088 32218 16144
rect 32274 16088 32279 16144
rect 30281 16086 32279 16088
rect 30281 16083 30347 16086
rect 32213 16083 32279 16086
rect 30833 16010 30899 16013
rect 31293 16010 31359 16013
rect 31845 16010 31911 16013
rect 30833 16008 31911 16010
rect 30833 15952 30838 16008
rect 30894 15952 31298 16008
rect 31354 15952 31850 16008
rect 31906 15952 31911 16008
rect 30833 15950 31911 15952
rect 30833 15947 30899 15950
rect 31293 15947 31359 15950
rect 31845 15947 31911 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 44173 15738 44239 15741
rect 44933 15738 45733 15768
rect 44173 15736 45733 15738
rect 44173 15680 44178 15736
rect 44234 15680 45733 15736
rect 44173 15678 45733 15680
rect 44173 15675 44239 15678
rect 44933 15648 45733 15678
rect 21541 15466 21607 15469
rect 23197 15466 23263 15469
rect 21541 15464 23263 15466
rect 21541 15408 21546 15464
rect 21602 15408 23202 15464
rect 23258 15408 23263 15464
rect 21541 15406 23263 15408
rect 21541 15403 21607 15406
rect 23197 15403 23263 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 16481 14514 16547 14517
rect 18597 14514 18663 14517
rect 16481 14512 18663 14514
rect 16481 14456 16486 14512
rect 16542 14456 18602 14512
rect 18658 14456 18663 14512
rect 16481 14454 18663 14456
rect 16481 14451 16547 14454
rect 18597 14451 18663 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 14089 13834 14155 13837
rect 17902 13834 17908 13836
rect 14089 13832 17908 13834
rect 14089 13776 14094 13832
rect 14150 13776 17908 13832
rect 14089 13774 17908 13776
rect 14089 13771 14155 13774
rect 17902 13772 17908 13774
rect 17972 13772 17978 13836
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 11789 13290 11855 13293
rect 22001 13290 22067 13293
rect 11789 13288 22067 13290
rect 11789 13232 11794 13288
rect 11850 13232 22006 13288
rect 22062 13232 22067 13288
rect 11789 13230 22067 13232
rect 11789 13227 11855 13230
rect 22001 13227 22067 13230
rect 23381 13154 23447 13157
rect 26969 13154 27035 13157
rect 23381 13152 27035 13154
rect 23381 13096 23386 13152
rect 23442 13096 26974 13152
rect 27030 13096 27035 13152
rect 23381 13094 27035 13096
rect 23381 13091 23447 13094
rect 26969 13091 27035 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 11881 13018 11947 13021
rect 18229 13018 18295 13021
rect 11881 13016 18295 13018
rect 11881 12960 11886 13016
rect 11942 12960 18234 13016
rect 18290 12960 18295 13016
rect 11881 12958 18295 12960
rect 11881 12955 11947 12958
rect 18229 12955 18295 12958
rect 22001 13018 22067 13021
rect 22461 13018 22527 13021
rect 25497 13018 25563 13021
rect 22001 13016 25563 13018
rect 22001 12960 22006 13016
rect 22062 12960 22466 13016
rect 22522 12960 25502 13016
rect 25558 12960 25563 13016
rect 22001 12958 25563 12960
rect 22001 12955 22067 12958
rect 22461 12955 22527 12958
rect 25497 12955 25563 12958
rect 14733 12882 14799 12885
rect 24945 12882 25011 12885
rect 26141 12882 26207 12885
rect 14733 12880 26207 12882
rect 14733 12824 14738 12880
rect 14794 12824 24950 12880
rect 25006 12824 26146 12880
rect 26202 12824 26207 12880
rect 14733 12822 26207 12824
rect 14733 12819 14799 12822
rect 24945 12819 25011 12822
rect 26141 12819 26207 12822
rect 31150 12820 31156 12884
rect 31220 12882 31226 12884
rect 31477 12882 31543 12885
rect 31220 12880 31543 12882
rect 31220 12824 31482 12880
rect 31538 12824 31543 12880
rect 31220 12822 31543 12824
rect 31220 12820 31226 12822
rect 31477 12819 31543 12822
rect 11973 12746 12039 12749
rect 17401 12746 17467 12749
rect 11973 12744 17467 12746
rect 11973 12688 11978 12744
rect 12034 12688 17406 12744
rect 17462 12688 17467 12744
rect 11973 12686 17467 12688
rect 11973 12683 12039 12686
rect 17401 12683 17467 12686
rect 15142 12548 15148 12612
rect 15212 12610 15218 12612
rect 15377 12610 15443 12613
rect 15212 12608 15443 12610
rect 15212 12552 15382 12608
rect 15438 12552 15443 12608
rect 15212 12550 15443 12552
rect 15212 12548 15218 12550
rect 15377 12547 15443 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 17902 12276 17908 12340
rect 17972 12338 17978 12340
rect 22093 12338 22159 12341
rect 17972 12336 22159 12338
rect 17972 12280 22098 12336
rect 22154 12280 22159 12336
rect 17972 12278 22159 12280
rect 17972 12276 17978 12278
rect 22093 12275 22159 12278
rect 14089 12202 14155 12205
rect 15653 12202 15719 12205
rect 14089 12200 15719 12202
rect 14089 12144 14094 12200
rect 14150 12144 15658 12200
rect 15714 12144 15719 12200
rect 14089 12142 15719 12144
rect 14089 12139 14155 12142
rect 15653 12139 15719 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 10041 11930 10107 11933
rect 14917 11930 14983 11933
rect 10041 11928 14983 11930
rect 10041 11872 10046 11928
rect 10102 11872 14922 11928
rect 14978 11872 14983 11928
rect 10041 11870 14983 11872
rect 10041 11867 10107 11870
rect 14917 11867 14983 11870
rect 11329 11522 11395 11525
rect 19517 11522 19583 11525
rect 11329 11520 19583 11522
rect 11329 11464 11334 11520
rect 11390 11464 19522 11520
rect 19578 11464 19583 11520
rect 11329 11462 19583 11464
rect 11329 11459 11395 11462
rect 19517 11459 19583 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 10041 11386 10107 11389
rect 10869 11386 10935 11389
rect 12525 11386 12591 11389
rect 10041 11384 12591 11386
rect 10041 11328 10046 11384
rect 10102 11328 10874 11384
rect 10930 11328 12530 11384
rect 12586 11328 12591 11384
rect 10041 11326 12591 11328
rect 10041 11323 10107 11326
rect 10869 11323 10935 11326
rect 12525 11323 12591 11326
rect 9857 11250 9923 11253
rect 10542 11250 10548 11252
rect 9857 11248 10548 11250
rect 9857 11192 9862 11248
rect 9918 11192 10548 11248
rect 9857 11190 10548 11192
rect 9857 11187 9923 11190
rect 10542 11188 10548 11190
rect 10612 11250 10618 11252
rect 15193 11250 15259 11253
rect 10612 11248 15259 11250
rect 10612 11192 15198 11248
rect 15254 11192 15259 11248
rect 10612 11190 15259 11192
rect 10612 11188 10618 11190
rect 15193 11187 15259 11190
rect 11329 11114 11395 11117
rect 14549 11114 14615 11117
rect 18045 11114 18111 11117
rect 11329 11112 18111 11114
rect 11329 11056 11334 11112
rect 11390 11056 14554 11112
rect 14610 11056 18050 11112
rect 18106 11056 18111 11112
rect 11329 11054 18111 11056
rect 11329 11051 11395 11054
rect 14549 11051 14615 11054
rect 18045 11051 18111 11054
rect 21265 11114 21331 11117
rect 27613 11114 27679 11117
rect 21265 11112 27679 11114
rect 21265 11056 21270 11112
rect 21326 11056 27618 11112
rect 27674 11056 27679 11112
rect 21265 11054 27679 11056
rect 21265 11051 21331 11054
rect 27613 11051 27679 11054
rect 10409 10978 10475 10981
rect 13905 10978 13971 10981
rect 10409 10976 13971 10978
rect 10409 10920 10414 10976
rect 10470 10920 13910 10976
rect 13966 10920 13971 10976
rect 10409 10918 13971 10920
rect 10409 10915 10475 10918
rect 13905 10915 13971 10918
rect 22093 10978 22159 10981
rect 22553 10978 22619 10981
rect 22093 10976 22619 10978
rect 22093 10920 22098 10976
rect 22154 10920 22558 10976
rect 22614 10920 22619 10976
rect 22093 10918 22619 10920
rect 22093 10915 22159 10918
rect 22553 10915 22619 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 22093 10706 22159 10709
rect 23013 10706 23079 10709
rect 22093 10704 23079 10706
rect 22093 10648 22098 10704
rect 22154 10648 23018 10704
rect 23074 10648 23079 10704
rect 22093 10646 23079 10648
rect 22093 10643 22159 10646
rect 23013 10643 23079 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 11973 10298 12039 10301
rect 12617 10298 12683 10301
rect 11973 10296 12683 10298
rect 11973 10240 11978 10296
rect 12034 10240 12622 10296
rect 12678 10240 12683 10296
rect 11973 10238 12683 10240
rect 11973 10235 12039 10238
rect 12617 10235 12683 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 11697 9754 11763 9757
rect 11830 9754 11836 9756
rect 11697 9752 11836 9754
rect 11697 9696 11702 9752
rect 11758 9696 11836 9752
rect 11697 9694 11836 9696
rect 11697 9691 11763 9694
rect 11830 9692 11836 9694
rect 11900 9692 11906 9756
rect 12157 9754 12223 9757
rect 17309 9754 17375 9757
rect 18781 9754 18847 9757
rect 12157 9752 18847 9754
rect 12157 9696 12162 9752
rect 12218 9696 17314 9752
rect 17370 9696 18786 9752
rect 18842 9696 18847 9752
rect 12157 9694 18847 9696
rect 12157 9691 12223 9694
rect 17309 9691 17375 9694
rect 18781 9691 18847 9694
rect 13261 9618 13327 9621
rect 14641 9618 14707 9621
rect 13261 9616 14707 9618
rect 13261 9560 13266 9616
rect 13322 9560 14646 9616
rect 14702 9560 14707 9616
rect 13261 9558 14707 9560
rect 13261 9555 13327 9558
rect 14641 9555 14707 9558
rect 13629 9482 13695 9485
rect 14181 9482 14247 9485
rect 13629 9480 14247 9482
rect 13629 9424 13634 9480
rect 13690 9424 14186 9480
rect 14242 9424 14247 9480
rect 13629 9422 14247 9424
rect 13629 9419 13695 9422
rect 14181 9419 14247 9422
rect 15837 9482 15903 9485
rect 16481 9482 16547 9485
rect 15837 9480 16547 9482
rect 15837 9424 15842 9480
rect 15898 9424 16486 9480
rect 16542 9424 16547 9480
rect 15837 9422 16547 9424
rect 15837 9419 15903 9422
rect 16481 9419 16547 9422
rect 13169 9346 13235 9349
rect 15285 9346 15351 9349
rect 13169 9344 15351 9346
rect 13169 9288 13174 9344
rect 13230 9288 15290 9344
rect 15346 9288 15351 9344
rect 13169 9286 15351 9288
rect 13169 9283 13235 9286
rect 15285 9283 15351 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 11513 9210 11579 9213
rect 15142 9210 15148 9212
rect 11513 9208 15148 9210
rect 11513 9152 11518 9208
rect 11574 9152 15148 9208
rect 11513 9150 15148 9152
rect 11513 9147 11579 9150
rect 15142 9148 15148 9150
rect 15212 9148 15218 9212
rect 10777 9074 10843 9077
rect 12525 9074 12591 9077
rect 10777 9072 12591 9074
rect 10777 9016 10782 9072
rect 10838 9016 12530 9072
rect 12586 9016 12591 9072
rect 10777 9014 12591 9016
rect 10777 9011 10843 9014
rect 12525 9011 12591 9014
rect 17585 9074 17651 9077
rect 18086 9074 18092 9076
rect 17585 9072 18092 9074
rect 17585 9016 17590 9072
rect 17646 9016 18092 9072
rect 17585 9014 18092 9016
rect 17585 9011 17651 9014
rect 18086 9012 18092 9014
rect 18156 9074 18162 9076
rect 18229 9074 18295 9077
rect 18873 9074 18939 9077
rect 18156 9072 18939 9074
rect 18156 9016 18234 9072
rect 18290 9016 18878 9072
rect 18934 9016 18939 9072
rect 18156 9014 18939 9016
rect 18156 9012 18162 9014
rect 18229 9011 18295 9014
rect 18873 9011 18939 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 13905 8938 13971 8941
rect 14917 8938 14983 8941
rect 13905 8936 14983 8938
rect 13905 8880 13910 8936
rect 13966 8880 14922 8936
rect 14978 8880 14983 8936
rect 13905 8878 14983 8880
rect 13905 8875 13971 8878
rect 14917 8875 14983 8878
rect 11513 8802 11579 8805
rect 14181 8802 14247 8805
rect 11513 8800 14247 8802
rect 11513 8744 11518 8800
rect 11574 8744 14186 8800
rect 14242 8744 14247 8800
rect 11513 8742 14247 8744
rect 11513 8739 11579 8742
rect 14181 8739 14247 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 28717 7442 28783 7445
rect 29453 7442 29519 7445
rect 28717 7440 29519 7442
rect 28717 7384 28722 7440
rect 28778 7384 29458 7440
rect 29514 7384 29519 7440
rect 28717 7382 29519 7384
rect 28717 7379 28783 7382
rect 29453 7379 29519 7382
rect 25313 7306 25379 7309
rect 26785 7306 26851 7309
rect 25313 7304 26851 7306
rect 25313 7248 25318 7304
rect 25374 7248 26790 7304
rect 26846 7248 26851 7304
rect 25313 7246 26851 7248
rect 25313 7243 25379 7246
rect 26785 7243 26851 7246
rect 10593 7170 10659 7173
rect 11697 7170 11763 7173
rect 10593 7168 11763 7170
rect 10593 7112 10598 7168
rect 10654 7112 11702 7168
rect 11758 7112 11763 7168
rect 10593 7110 11763 7112
rect 10593 7107 10659 7110
rect 11697 7107 11763 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 10501 6900 10567 6901
rect 10501 6898 10548 6900
rect 10456 6896 10548 6898
rect 10612 6898 10618 6900
rect 44081 6898 44147 6901
rect 44933 6898 45733 6928
rect 10456 6840 10506 6896
rect 10456 6838 10548 6840
rect 10501 6836 10548 6838
rect 10612 6838 12450 6898
rect 10612 6836 10618 6838
rect 10501 6835 10567 6836
rect 12390 6626 12450 6838
rect 44081 6896 45733 6898
rect 44081 6840 44086 6896
rect 44142 6840 45733 6896
rect 44081 6838 45733 6840
rect 44081 6835 44147 6838
rect 44933 6808 45733 6838
rect 15745 6626 15811 6629
rect 12390 6624 15811 6626
rect 12390 6568 15750 6624
rect 15806 6568 15811 6624
rect 12390 6566 15811 6568
rect 15745 6563 15811 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 11881 6490 11947 6493
rect 15101 6490 15167 6493
rect 17309 6490 17375 6493
rect 11881 6488 17375 6490
rect 11881 6432 11886 6488
rect 11942 6432 15106 6488
rect 15162 6432 17314 6488
rect 17370 6432 17375 6488
rect 11881 6430 17375 6432
rect 11881 6427 11947 6430
rect 15101 6427 15167 6430
rect 17309 6427 17375 6430
rect 4797 6354 4863 6357
rect 8201 6354 8267 6357
rect 4797 6352 8267 6354
rect 4797 6296 4802 6352
rect 4858 6296 8206 6352
rect 8262 6296 8267 6352
rect 4797 6294 8267 6296
rect 4797 6291 4863 6294
rect 8201 6291 8267 6294
rect 14917 6354 14983 6357
rect 17585 6354 17651 6357
rect 14917 6352 17651 6354
rect 14917 6296 14922 6352
rect 14978 6296 17590 6352
rect 17646 6296 17651 6352
rect 14917 6294 17651 6296
rect 14917 6291 14983 6294
rect 17585 6291 17651 6294
rect 13353 6218 13419 6221
rect 15561 6218 15627 6221
rect 18045 6218 18111 6221
rect 13353 6216 18111 6218
rect 13353 6160 13358 6216
rect 13414 6160 15566 6216
rect 15622 6160 18050 6216
rect 18106 6160 18111 6216
rect 13353 6158 18111 6160
rect 13353 6155 13419 6158
rect 15561 6155 15627 6158
rect 18045 6155 18111 6158
rect 12249 6082 12315 6085
rect 13721 6082 13787 6085
rect 12249 6080 13787 6082
rect 12249 6024 12254 6080
rect 12310 6024 13726 6080
rect 13782 6024 13787 6080
rect 12249 6022 13787 6024
rect 12249 6019 12315 6022
rect 13721 6019 13787 6022
rect 17125 6082 17191 6085
rect 17861 6082 17927 6085
rect 17125 6080 17927 6082
rect 17125 6024 17130 6080
rect 17186 6024 17866 6080
rect 17922 6024 17927 6080
rect 17125 6022 17927 6024
rect 17125 6019 17191 6022
rect 17861 6019 17927 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 13537 5946 13603 5949
rect 19333 5946 19399 5949
rect 13537 5944 19399 5946
rect 13537 5888 13542 5944
rect 13598 5888 19338 5944
rect 19394 5888 19399 5944
rect 13537 5886 19399 5888
rect 13537 5883 13603 5886
rect 19333 5883 19399 5886
rect 13537 5674 13603 5677
rect 17493 5674 17559 5677
rect 19333 5674 19399 5677
rect 13537 5672 19399 5674
rect 13537 5616 13542 5672
rect 13598 5616 17498 5672
rect 17554 5616 19338 5672
rect 19394 5616 19399 5672
rect 13537 5614 19399 5616
rect 13537 5611 13603 5614
rect 17493 5611 17559 5614
rect 19333 5611 19399 5614
rect 11881 5540 11947 5541
rect 11830 5476 11836 5540
rect 11900 5538 11947 5540
rect 13905 5538 13971 5541
rect 16757 5538 16823 5541
rect 18137 5540 18203 5541
rect 18086 5538 18092 5540
rect 11900 5536 11992 5538
rect 11942 5480 11992 5536
rect 11900 5478 11992 5480
rect 13905 5536 16823 5538
rect 13905 5480 13910 5536
rect 13966 5480 16762 5536
rect 16818 5480 16823 5536
rect 13905 5478 16823 5480
rect 18046 5478 18092 5538
rect 18156 5536 18203 5540
rect 31109 5540 31175 5541
rect 31109 5538 31156 5540
rect 18198 5480 18203 5536
rect 11900 5476 11947 5478
rect 11881 5475 11947 5476
rect 13905 5475 13971 5478
rect 16757 5475 16823 5478
rect 18086 5476 18092 5478
rect 18156 5476 18203 5480
rect 31064 5536 31156 5538
rect 31064 5480 31114 5536
rect 31064 5478 31156 5480
rect 18137 5475 18203 5476
rect 31109 5476 31156 5478
rect 31220 5476 31226 5540
rect 31109 5475 31175 5476
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 15009 5402 15075 5405
rect 15142 5402 15148 5404
rect 15009 5400 15148 5402
rect 15009 5344 15014 5400
rect 15070 5344 15148 5400
rect 15009 5342 15148 5344
rect 15009 5339 15075 5342
rect 15142 5340 15148 5342
rect 15212 5402 15218 5404
rect 17125 5402 17191 5405
rect 15212 5400 17191 5402
rect 15212 5344 17130 5400
rect 17186 5344 17191 5400
rect 15212 5342 17191 5344
rect 15212 5340 15218 5342
rect 17125 5339 17191 5342
rect 11881 4994 11947 4997
rect 18229 4994 18295 4997
rect 11881 4992 18295 4994
rect 11881 4936 11886 4992
rect 11942 4936 18234 4992
rect 18290 4936 18295 4992
rect 11881 4934 18295 4936
rect 11881 4931 11947 4934
rect 18229 4931 18295 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 15561 4450 15627 4453
rect 16481 4450 16547 4453
rect 17861 4450 17927 4453
rect 15561 4448 17927 4450
rect 15561 4392 15566 4448
rect 15622 4392 16486 4448
rect 16542 4392 17866 4448
rect 17922 4392 17927 4448
rect 15561 4390 17927 4392
rect 15561 4387 15627 4390
rect 16481 4387 16547 4390
rect 17861 4387 17927 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 10409 4314 10475 4317
rect 14917 4314 14983 4317
rect 10409 4312 14983 4314
rect 10409 4256 10414 4312
rect 10470 4256 14922 4312
rect 14978 4256 14983 4312
rect 10409 4254 14983 4256
rect 10409 4251 10475 4254
rect 14917 4251 14983 4254
rect 11421 4178 11487 4181
rect 17585 4178 17651 4181
rect 11421 4176 17651 4178
rect 11421 4120 11426 4176
rect 11482 4120 17590 4176
rect 17646 4120 17651 4176
rect 11421 4118 17651 4120
rect 11421 4115 11487 4118
rect 17585 4115 17651 4118
rect 18321 4178 18387 4181
rect 19057 4178 19123 4181
rect 18321 4176 19123 4178
rect 18321 4120 18326 4176
rect 18382 4120 19062 4176
rect 19118 4120 19123 4176
rect 18321 4118 19123 4120
rect 18321 4115 18387 4118
rect 19057 4115 19123 4118
rect 22921 4178 22987 4181
rect 24485 4178 24551 4181
rect 22921 4176 24551 4178
rect 22921 4120 22926 4176
rect 22982 4120 24490 4176
rect 24546 4120 24551 4176
rect 22921 4118 24551 4120
rect 22921 4115 22987 4118
rect 24485 4115 24551 4118
rect 12249 4042 12315 4045
rect 12893 4042 12959 4045
rect 18137 4042 18203 4045
rect 12249 4040 18203 4042
rect 12249 3984 12254 4040
rect 12310 3984 12898 4040
rect 12954 3984 18142 4040
rect 18198 3984 18203 4040
rect 12249 3982 18203 3984
rect 12249 3979 12315 3982
rect 12893 3979 12959 3982
rect 18137 3979 18203 3982
rect 13261 3906 13327 3909
rect 13813 3906 13879 3909
rect 16941 3906 17007 3909
rect 13261 3904 17007 3906
rect 13261 3848 13266 3904
rect 13322 3848 13818 3904
rect 13874 3848 16946 3904
rect 17002 3848 17007 3904
rect 13261 3846 17007 3848
rect 13261 3843 13327 3846
rect 13813 3843 13879 3846
rect 16941 3843 17007 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 12249 3498 12315 3501
rect 14825 3498 14891 3501
rect 12249 3496 14891 3498
rect 12249 3440 12254 3496
rect 12310 3440 14830 3496
rect 14886 3440 14891 3496
rect 12249 3438 14891 3440
rect 12249 3435 12315 3438
rect 14825 3435 14891 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 8753 3090 8819 3093
rect 18689 3090 18755 3093
rect 8753 3088 18755 3090
rect 8753 3032 8758 3088
rect 8814 3032 18694 3088
rect 18750 3032 18755 3088
rect 8753 3030 18755 3032
rect 8753 3027 8819 3030
rect 18689 3027 18755 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 20116 30832 20180 30836
rect 20116 30776 20166 30832
rect 20166 30776 20180 30832
rect 20116 30772 20180 30776
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 20116 30092 20180 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 17908 13772 17972 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 31156 12820 31220 12884
rect 15148 12548 15212 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 17908 12276 17972 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 10548 11188 10612 11252
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 11836 9692 11900 9756
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 15148 9148 15212 9212
rect 18092 9012 18156 9076
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 10548 6896 10612 6900
rect 10548 6840 10562 6896
rect 10562 6840 10612 6896
rect 10548 6836 10612 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 11836 5536 11900 5540
rect 11836 5480 11886 5536
rect 11886 5480 11900 5536
rect 11836 5476 11900 5480
rect 18092 5536 18156 5540
rect 18092 5480 18142 5536
rect 18142 5480 18156 5536
rect 18092 5476 18156 5480
rect 31156 5536 31220 5540
rect 31156 5480 31170 5536
rect 31170 5480 31220 5536
rect 31156 5476 31220 5480
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 15148 5340 15212 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 45184 4528 45744
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 19568 45728 19888 45744
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 34928 45184 35248 45744
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 20115 30836 20181 30837
rect 20115 30772 20116 30836
rect 20180 30772 20181 30836
rect 20115 30771 20181 30772
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 20118 30157 20178 30771
rect 20115 30156 20181 30157
rect 20115 30092 20116 30156
rect 20180 30092 20181 30156
rect 20115 30091 20181 30092
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 17907 13836 17973 13837
rect 17907 13772 17908 13836
rect 17972 13772 17973 13836
rect 17907 13771 17973 13772
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 15147 12612 15213 12613
rect 15147 12548 15148 12612
rect 15212 12548 15213 12612
rect 15147 12547 15213 12548
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 10547 11252 10613 11253
rect 10547 11188 10548 11252
rect 10612 11188 10613 11252
rect 10547 11187 10613 11188
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 10550 6901 10610 11187
rect 11835 9756 11901 9757
rect 11835 9692 11836 9756
rect 11900 9692 11901 9756
rect 11835 9691 11901 9692
rect 10547 6900 10613 6901
rect 10547 6836 10548 6900
rect 10612 6836 10613 6900
rect 10547 6835 10613 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 11838 5541 11898 9691
rect 15150 9213 15210 12547
rect 17910 12341 17970 13771
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 19568 12000 19888 13024
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 31155 12884 31221 12885
rect 31155 12820 31156 12884
rect 31220 12820 31221 12884
rect 31155 12819 31221 12820
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 15147 9212 15213 9213
rect 15147 9148 15148 9212
rect 15212 9148 15213 9212
rect 15147 9147 15213 9148
rect 11835 5540 11901 5541
rect 11835 5476 11836 5540
rect 11900 5476 11901 5540
rect 11835 5475 11901 5476
rect 15150 5405 15210 9147
rect 18091 9076 18157 9077
rect 18091 9012 18092 9076
rect 18156 9012 18157 9076
rect 18091 9011 18157 9012
rect 18094 5541 18154 9011
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 18091 5540 18157 5541
rect 18091 5476 18092 5540
rect 18156 5476 18157 5540
rect 18091 5475 18157 5476
rect 19568 5472 19888 6496
rect 31158 5541 31218 12819
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 31155 5540 31221 5541
rect 31155 5476 31156 5540
rect 31220 5476 31221 5540
rect 31155 5475 31221 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 15147 5404 15213 5405
rect 15147 5340 15148 5404
rect 15212 5340 15213 5404
rect 15147 5339 15213 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__and3_1  _1239_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38640 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1240_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36156 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1241_
timestamp 1688980957
transform -1 0 34868 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1242_
timestamp 1688980957
transform -1 0 36248 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1243_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35604 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1244_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28520 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1246_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27600 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1247_
timestamp 1688980957
transform -1 0 26496 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1248_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1249_
timestamp 1688980957
transform 1 0 34684 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1250_
timestamp 1688980957
transform -1 0 28060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1251_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_1  _1252_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36432 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1253_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36248 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1254_
timestamp 1688980957
transform -1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1688980957
transform -1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1256_
timestamp 1688980957
transform 1 0 36064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1688980957
transform -1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1258_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1688980957
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1260_
timestamp 1688980957
transform 1 0 18400 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1688980957
transform -1 0 19780 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1262_
timestamp 1688980957
transform 1 0 36156 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1688980957
transform -1 0 36984 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1264_
timestamp 1688980957
transform 1 0 5612 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1688980957
transform -1 0 6624 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1266_
timestamp 1688980957
transform 1 0 31556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1267_
timestamp 1688980957
transform 1 0 31648 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1268_
timestamp 1688980957
transform 1 0 25576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1269_
timestamp 1688980957
transform -1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1270_
timestamp 1688980957
transform -1 0 5428 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1272_
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1688980957
transform -1 0 25208 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1274_
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1688980957
transform -1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1276_
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1688980957
transform -1 0 2852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1278_
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1688980957
transform -1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1280_
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1688980957
transform -1 0 43608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1282_
timestamp 1688980957
transform 1 0 1748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1688980957
transform -1 0 2944 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1284_
timestamp 1688980957
transform 1 0 43332 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1688980957
transform 1 0 43332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1286_
timestamp 1688980957
transform -1 0 43792 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1688980957
transform -1 0 43608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1688980957
transform -1 0 34132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34408 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1290_
timestamp 1688980957
transform -1 0 36984 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35328 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36432 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1688980957
transform -1 0 35788 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1294_
timestamp 1688980957
transform -1 0 34960 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1688980957
transform 1 0 35052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1296_
timestamp 1688980957
transform 1 0 34776 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1297_
timestamp 1688980957
transform -1 0 35880 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1298_
timestamp 1688980957
transform -1 0 36340 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36524 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1301_
timestamp 1688980957
transform 1 0 37720 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1302_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43148 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1303_
timestamp 1688980957
transform 1 0 40020 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1304_
timestamp 1688980957
transform 1 0 41216 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40296 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42412 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41032 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1308_
timestamp 1688980957
transform -1 0 40848 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1309_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35972 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1310_
timestamp 1688980957
transform 1 0 37812 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1311_
timestamp 1688980957
transform 1 0 37996 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1688980957
transform 1 0 37720 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1688980957
transform -1 0 38548 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _1314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 41032 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1315_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1316_
timestamp 1688980957
transform -1 0 38272 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1317_
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1688980957
transform 1 0 40112 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1319_
timestamp 1688980957
transform -1 0 40296 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1320_
timestamp 1688980957
transform -1 0 40480 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1688980957
transform 1 0 40480 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1322_
timestamp 1688980957
transform -1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1323_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 39100 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1324_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 39560 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1325_
timestamp 1688980957
transform -1 0 39560 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1327_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1328_
timestamp 1688980957
transform -1 0 40664 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1329_
timestamp 1688980957
transform 1 0 40664 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1330_
timestamp 1688980957
transform 1 0 40020 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1688980957
transform 1 0 40572 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1688980957
transform 1 0 41400 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1333_
timestamp 1688980957
transform 1 0 41952 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1334_
timestamp 1688980957
transform 1 0 41860 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1688980957
transform -1 0 42320 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1336_
timestamp 1688980957
transform -1 0 44344 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1337_
timestamp 1688980957
transform -1 0 43056 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1338_
timestamp 1688980957
transform -1 0 43424 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1688980957
transform -1 0 43516 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1340_
timestamp 1688980957
transform -1 0 43700 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1341_
timestamp 1688980957
transform -1 0 42412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1342_
timestamp 1688980957
transform -1 0 39376 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1343_
timestamp 1688980957
transform -1 0 39744 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1344_
timestamp 1688980957
transform -1 0 40296 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1345_
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1346_
timestamp 1688980957
transform 1 0 40296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1347_
timestamp 1688980957
transform -1 0 41032 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1348_
timestamp 1688980957
transform -1 0 40388 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1349_
timestamp 1688980957
transform 1 0 41308 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 1688980957
transform 1 0 41860 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1351_
timestamp 1688980957
transform -1 0 43056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1352_
timestamp 1688980957
transform -1 0 43608 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1688980957
transform -1 0 42320 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1688980957
transform -1 0 43240 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1355_
timestamp 1688980957
transform 1 0 42044 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1688980957
transform -1 0 41860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1357_
timestamp 1688980957
transform 1 0 42412 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1358_
timestamp 1688980957
transform -1 0 37168 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1359_
timestamp 1688980957
transform 1 0 33672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361_
timestamp 1688980957
transform -1 0 43424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1362_
timestamp 1688980957
transform -1 0 43240 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1363_
timestamp 1688980957
transform -1 0 43700 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1364_
timestamp 1688980957
transform -1 0 43424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1365_
timestamp 1688980957
transform -1 0 42504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1366_
timestamp 1688980957
transform -1 0 42044 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1367_
timestamp 1688980957
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1688980957
transform -1 0 42044 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1369_
timestamp 1688980957
transform 1 0 39652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1370_
timestamp 1688980957
transform -1 0 40296 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1371_
timestamp 1688980957
transform 1 0 39376 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1688980957
transform -1 0 39376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1373_
timestamp 1688980957
transform -1 0 39376 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1688980957
transform -1 0 37904 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1375_
timestamp 1688980957
transform -1 0 38364 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 1688980957
transform -1 0 37076 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1377_
timestamp 1688980957
transform -1 0 37904 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1378_
timestamp 1688980957
transform -1 0 36708 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1379_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1688980957
transform -1 0 25944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1381_
timestamp 1688980957
transform -1 0 25484 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1382_
timestamp 1688980957
transform 1 0 31924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1383_
timestamp 1688980957
transform -1 0 35880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1384_
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1385_
timestamp 1688980957
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1386_
timestamp 1688980957
transform -1 0 37168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1688980957
transform -1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1388_
timestamp 1688980957
transform -1 0 35696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1389_
timestamp 1688980957
transform -1 0 34592 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1390_
timestamp 1688980957
transform -1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1391_
timestamp 1688980957
transform -1 0 35144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1392_
timestamp 1688980957
transform 1 0 34684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1393_
timestamp 1688980957
transform 1 0 34960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1394_
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1395_
timestamp 1688980957
transform -1 0 34960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1688980957
transform 1 0 35328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1397_
timestamp 1688980957
transform -1 0 20976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1688980957
transform 1 0 9292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1399_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1400_
timestamp 1688980957
transform 1 0 11868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1401_
timestamp 1688980957
transform -1 0 22080 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1402_
timestamp 1688980957
transform 1 0 10396 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1403_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1688980957
transform -1 0 11500 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1405_
timestamp 1688980957
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1406_
timestamp 1688980957
transform 1 0 10948 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1407_
timestamp 1688980957
transform 1 0 11500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1688980957
transform -1 0 12604 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1409_
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1410_
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1411_
timestamp 1688980957
transform 1 0 15088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412_
timestamp 1688980957
transform -1 0 16468 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1688980957
transform -1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1414_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1688980957
transform -1 0 15548 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1688980957
transform 1 0 18768 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1688980957
transform -1 0 14628 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1418_
timestamp 1688980957
transform 1 0 14168 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1688980957
transform -1 0 14996 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1420_
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1688980957
transform 1 0 11224 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1422_
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1688980957
transform 1 0 11592 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1688980957
transform -1 0 19228 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1425_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1426_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14260 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1427_
timestamp 1688980957
transform -1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428_
timestamp 1688980957
transform 1 0 11960 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1429_
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1430_
timestamp 1688980957
transform -1 0 13156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1431_
timestamp 1688980957
transform 1 0 13616 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1432_
timestamp 1688980957
transform 1 0 14996 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1433_
timestamp 1688980957
transform -1 0 13616 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1434_
timestamp 1688980957
transform -1 0 12880 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1435_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1436_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1437_
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1438_
timestamp 1688980957
transform -1 0 10764 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 1688980957
transform -1 0 9292 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1440_
timestamp 1688980957
transform 1 0 9844 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1442_
timestamp 1688980957
transform 1 0 9016 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1443_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 1688980957
transform -1 0 9016 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1688980957
transform -1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1446_
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1688980957
transform 1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1688980957
transform -1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1449_
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1688980957
transform -1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1688980957
transform -1 0 6900 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1452_
timestamp 1688980957
transform -1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1688980957
transform -1 0 5888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1454_
timestamp 1688980957
transform -1 0 7360 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1455_
timestamp 1688980957
transform -1 0 6256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1456_
timestamp 1688980957
transform 1 0 5336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1457_
timestamp 1688980957
transform -1 0 6624 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1458_
timestamp 1688980957
transform -1 0 6164 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1459_
timestamp 1688980957
transform -1 0 5888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1688980957
transform -1 0 5612 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 1688980957
transform 1 0 5704 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1463_
timestamp 1688980957
transform 1 0 5336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 1688980957
transform 1 0 5888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1466_
timestamp 1688980957
transform 1 0 6624 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1467_
timestamp 1688980957
transform -1 0 7544 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1468_
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1688980957
transform 1 0 7544 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1471_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1472_
timestamp 1688980957
transform 1 0 8004 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1688980957
transform -1 0 8556 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1474_
timestamp 1688980957
transform 1 0 8280 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1475_
timestamp 1688980957
transform 1 0 7636 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1476_
timestamp 1688980957
transform 1 0 7820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1477_
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1478_
timestamp 1688980957
transform -1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1479_
timestamp 1688980957
transform 1 0 8280 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1688980957
transform -1 0 6256 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1481_
timestamp 1688980957
transform -1 0 6808 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1482_
timestamp 1688980957
transform -1 0 5796 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1483_
timestamp 1688980957
transform -1 0 5704 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1688980957
transform 1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1485_
timestamp 1688980957
transform -1 0 6072 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1487_
timestamp 1688980957
transform 1 0 5428 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1688980957
transform 1 0 5888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1489_
timestamp 1688980957
transform -1 0 7268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1490_
timestamp 1688980957
transform -1 0 6348 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1491_
timestamp 1688980957
transform 1 0 4968 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1492_
timestamp 1688980957
transform 1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1688980957
transform -1 0 8556 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1494_
timestamp 1688980957
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1495_
timestamp 1688980957
transform -1 0 8096 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1497_
timestamp 1688980957
transform 1 0 8096 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1498_
timestamp 1688980957
transform -1 0 9660 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1499_
timestamp 1688980957
transform -1 0 8648 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1500_
timestamp 1688980957
transform -1 0 9016 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1501_
timestamp 1688980957
transform -1 0 9292 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 1688980957
transform -1 0 40848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1503_
timestamp 1688980957
transform 1 0 39100 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1504_
timestamp 1688980957
transform 1 0 39100 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1688980957
transform -1 0 39836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1506_
timestamp 1688980957
transform -1 0 39560 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1507_
timestamp 1688980957
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1508_
timestamp 1688980957
transform -1 0 5980 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1509_
timestamp 1688980957
transform -1 0 6164 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1510_
timestamp 1688980957
transform 1 0 5336 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1511_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 1688980957
transform -1 0 37996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1513_
timestamp 1688980957
transform 1 0 33396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1515_
timestamp 1688980957
transform -1 0 34500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1688980957
transform 1 0 33672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1517_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43424 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1519_
timestamp 1688980957
transform -1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1688980957
transform -1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1521_
timestamp 1688980957
transform 1 0 20240 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1522_
timestamp 1688980957
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1523_
timestamp 1688980957
transform -1 0 20792 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20056 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1525_
timestamp 1688980957
transform 1 0 12052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1526_
timestamp 1688980957
transform 1 0 12328 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1688980957
transform -1 0 12972 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1528_
timestamp 1688980957
transform 1 0 14904 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1529_
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1530_
timestamp 1688980957
transform 1 0 12420 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1531_
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 1688980957
transform 1 0 12972 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1534_
timestamp 1688980957
transform -1 0 11684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1535_
timestamp 1688980957
transform -1 0 12052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1536_
timestamp 1688980957
transform -1 0 14352 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1537_
timestamp 1688980957
transform 1 0 12420 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1538_
timestamp 1688980957
transform 1 0 13156 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1539_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1540_
timestamp 1688980957
transform -1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1541_
timestamp 1688980957
transform 1 0 20884 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1542_
timestamp 1688980957
transform -1 0 22356 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1688980957
transform -1 0 21712 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1688980957
transform -1 0 20976 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1545_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1546_
timestamp 1688980957
transform -1 0 20700 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1547_
timestamp 1688980957
transform 1 0 19780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1548_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 1688980957
transform -1 0 20608 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1550_
timestamp 1688980957
transform -1 0 20148 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1551_
timestamp 1688980957
transform 1 0 19872 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1688980957
transform -1 0 21436 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1553_
timestamp 1688980957
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1554_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1555_
timestamp 1688980957
transform 1 0 20608 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1556_
timestamp 1688980957
transform -1 0 19228 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1557_
timestamp 1688980957
transform -1 0 19136 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1558_
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1559_
timestamp 1688980957
transform -1 0 19872 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1560_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1561_
timestamp 1688980957
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1562_
timestamp 1688980957
transform -1 0 12420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1563_
timestamp 1688980957
transform -1 0 13984 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1564_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13708 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1565_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_2  _1566_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1567_
timestamp 1688980957
transform -1 0 21344 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1568_
timestamp 1688980957
transform -1 0 20884 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1569_
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1570_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1571_
timestamp 1688980957
transform -1 0 20884 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1572_
timestamp 1688980957
transform 1 0 19412 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_2  _1573_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21712 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1574_
timestamp 1688980957
transform 1 0 41492 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1575_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 1688980957
transform -1 0 41492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1577_
timestamp 1688980957
transform 1 0 40848 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1578_
timestamp 1688980957
transform 1 0 39008 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1579_
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1580_
timestamp 1688980957
transform -1 0 39008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1581_
timestamp 1688980957
transform -1 0 40480 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _1582_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1583_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1584_
timestamp 1688980957
transform 1 0 40480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40388 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1586_
timestamp 1688980957
transform 1 0 42780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1587_
timestamp 1688980957
transform -1 0 43332 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1588_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42320 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1589_
timestamp 1688980957
transform 1 0 43332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1590_
timestamp 1688980957
transform -1 0 43240 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1591_
timestamp 1688980957
transform 1 0 43240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1592_
timestamp 1688980957
transform 1 0 42780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_2  _1593_
timestamp 1688980957
transform 1 0 41676 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1594_
timestamp 1688980957
transform -1 0 42964 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1595_
timestamp 1688980957
transform -1 0 42872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1596_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43056 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1597_
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1598_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42964 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1599_
timestamp 1688980957
transform 1 0 43056 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1600_
timestamp 1688980957
transform -1 0 43056 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1601_
timestamp 1688980957
transform -1 0 42136 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1688980957
transform -1 0 41952 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1603_
timestamp 1688980957
transform -1 0 42044 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1688980957
transform -1 0 41584 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1605_
timestamp 1688980957
transform -1 0 40388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1606_
timestamp 1688980957
transform 1 0 39376 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1607_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 40296 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1688980957
transform 1 0 39100 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1609_
timestamp 1688980957
transform 1 0 39376 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1610_
timestamp 1688980957
transform -1 0 39192 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1611_
timestamp 1688980957
transform -1 0 38548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1612_
timestamp 1688980957
transform 1 0 38824 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1613_
timestamp 1688980957
transform -1 0 39100 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1614_
timestamp 1688980957
transform 1 0 38732 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1615_
timestamp 1688980957
transform -1 0 39836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38088 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1617_
timestamp 1688980957
transform 1 0 29900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1619_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1620_
timestamp 1688980957
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1621_
timestamp 1688980957
transform 1 0 32660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1622_
timestamp 1688980957
transform -1 0 39100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1623_
timestamp 1688980957
transform 1 0 40848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1624_
timestamp 1688980957
transform -1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1625_
timestamp 1688980957
transform -1 0 22724 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1626_
timestamp 1688980957
transform -1 0 22540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1627_
timestamp 1688980957
transform -1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1628_
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_2  _1629_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33764 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1630_
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1631_
timestamp 1688980957
transform -1 0 24104 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1632_
timestamp 1688980957
transform -1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1633_
timestamp 1688980957
transform -1 0 26404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1634_
timestamp 1688980957
transform -1 0 26680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 1688980957
transform -1 0 24932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1636_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23920 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1637_
timestamp 1688980957
transform 1 0 23276 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1638_
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1639_
timestamp 1688980957
transform 1 0 22908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1640_
timestamp 1688980957
transform 1 0 22356 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1641_
timestamp 1688980957
transform -1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23000 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1643_
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1644_
timestamp 1688980957
transform 1 0 22080 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1645_
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1646_
timestamp 1688980957
transform 1 0 23368 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1647_
timestamp 1688980957
transform 1 0 33672 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1648_
timestamp 1688980957
transform -1 0 35144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1649_
timestamp 1688980957
transform -1 0 34868 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1650_
timestamp 1688980957
transform -1 0 35052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1651_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1652_
timestamp 1688980957
transform 1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1653_
timestamp 1688980957
transform -1 0 32660 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1654_
timestamp 1688980957
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1688980957
transform 1 0 33028 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1656_
timestamp 1688980957
transform -1 0 33856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1657_
timestamp 1688980957
transform 1 0 33856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1658_
timestamp 1688980957
transform -1 0 35328 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1660_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1688980957
transform -1 0 35604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1662_
timestamp 1688980957
transform -1 0 31832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1663_
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1664_
timestamp 1688980957
transform 1 0 33672 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1665_
timestamp 1688980957
transform 1 0 33396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1667_
timestamp 1688980957
transform 1 0 34224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1668_
timestamp 1688980957
transform 1 0 34132 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1669_
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1670_
timestamp 1688980957
transform -1 0 34684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1671_
timestamp 1688980957
transform -1 0 33028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1672_
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1673_
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1674_
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1675_
timestamp 1688980957
transform -1 0 34500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1676_
timestamp 1688980957
transform 1 0 34500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1677_
timestamp 1688980957
transform 1 0 33672 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1678_
timestamp 1688980957
transform -1 0 36064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1679_
timestamp 1688980957
transform 1 0 32660 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1680_
timestamp 1688980957
transform 1 0 33396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1681_
timestamp 1688980957
transform -1 0 34408 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1682_
timestamp 1688980957
transform -1 0 34500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1683_
timestamp 1688980957
transform 1 0 25668 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1684_
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1685_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1686_
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1687_
timestamp 1688980957
transform -1 0 34592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1688_
timestamp 1688980957
transform 1 0 35328 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1689_
timestamp 1688980957
transform 1 0 33580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1688980957
transform -1 0 34776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1691_
timestamp 1688980957
transform 1 0 33488 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1688980957
transform -1 0 34408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1693_
timestamp 1688980957
transform 1 0 25944 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1694_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25668 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1695_
timestamp 1688980957
transform 1 0 32200 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1696_
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1697_
timestamp 1688980957
transform 1 0 33396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1698_
timestamp 1688980957
transform -1 0 33580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1688980957
transform -1 0 32016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1700_
timestamp 1688980957
transform 1 0 25484 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1701_
timestamp 1688980957
transform -1 0 27692 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1702_
timestamp 1688980957
transform 1 0 27048 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1703_
timestamp 1688980957
transform -1 0 31188 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1704_
timestamp 1688980957
transform 1 0 31188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1705_
timestamp 1688980957
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1706_
timestamp 1688980957
transform 1 0 33120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1707_
timestamp 1688980957
transform -1 0 34224 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1708_
timestamp 1688980957
transform 1 0 32568 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1709_
timestamp 1688980957
transform -1 0 32660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1710_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32660 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1711_
timestamp 1688980957
transform -1 0 30268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1712_
timestamp 1688980957
transform -1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1713_
timestamp 1688980957
transform 1 0 29256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1715_
timestamp 1688980957
transform -1 0 26496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1716_
timestamp 1688980957
transform 1 0 26496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1717_
timestamp 1688980957
transform -1 0 29900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1718_
timestamp 1688980957
transform 1 0 28980 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1719_
timestamp 1688980957
transform 1 0 30360 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1720_
timestamp 1688980957
transform 1 0 30084 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1721_
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1722_
timestamp 1688980957
transform -1 0 31740 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1723_
timestamp 1688980957
transform 1 0 29532 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1724_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30360 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1725_
timestamp 1688980957
transform -1 0 31188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1726_
timestamp 1688980957
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1727_
timestamp 1688980957
transform -1 0 26404 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1728_
timestamp 1688980957
transform -1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1729_
timestamp 1688980957
transform 1 0 25576 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1730_
timestamp 1688980957
transform 1 0 28704 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1731_
timestamp 1688980957
transform -1 0 30452 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1732_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29992 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1733_
timestamp 1688980957
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1734_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29164 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1735_
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1736_
timestamp 1688980957
transform 1 0 25576 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1737_
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1738_
timestamp 1688980957
transform 1 0 28244 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp 1688980957
transform 1 0 29532 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1740_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1741_
timestamp 1688980957
transform -1 0 29348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1742_
timestamp 1688980957
transform 1 0 28336 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1743_
timestamp 1688980957
transform -1 0 28980 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1744_
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1745_
timestamp 1688980957
transform 1 0 24656 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1746_
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1747_
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1748_
timestamp 1688980957
transform 1 0 30084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1749_
timestamp 1688980957
transform -1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_4  _1750_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28980 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1751_
timestamp 1688980957
transform -1 0 32384 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1752_
timestamp 1688980957
transform -1 0 30544 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1753_
timestamp 1688980957
transform 1 0 29348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1754_
timestamp 1688980957
transform 1 0 25852 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1755_
timestamp 1688980957
transform 1 0 25208 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1756_
timestamp 1688980957
transform 1 0 26772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1757_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1758_
timestamp 1688980957
transform 1 0 30544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1759_
timestamp 1688980957
transform 1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1760_
timestamp 1688980957
transform -1 0 31648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1761_
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1762_
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1688980957
transform -1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1764_
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1765_
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1688980957
transform -1 0 31832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1767_
timestamp 1688980957
transform 1 0 25392 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1768_
timestamp 1688980957
transform 1 0 27600 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1769_
timestamp 1688980957
transform 1 0 26864 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1770_
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1771_
timestamp 1688980957
transform 1 0 28520 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1772_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1773_
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1774_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29348 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1775_
timestamp 1688980957
transform -1 0 29808 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1776_
timestamp 1688980957
transform -1 0 29808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1777_
timestamp 1688980957
transform 1 0 28796 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1778_
timestamp 1688980957
transform 1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1779_
timestamp 1688980957
transform -1 0 26404 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1780_
timestamp 1688980957
transform 1 0 26220 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1781_
timestamp 1688980957
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1782_
timestamp 1688980957
transform 1 0 28152 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1783_
timestamp 1688980957
transform 1 0 28888 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1784_
timestamp 1688980957
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1785_
timestamp 1688980957
transform 1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1786_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1787_
timestamp 1688980957
transform 1 0 32752 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1788_
timestamp 1688980957
transform 1 0 25668 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1789_
timestamp 1688980957
transform 1 0 25576 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1790_
timestamp 1688980957
transform 1 0 31464 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1791_
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1792_
timestamp 1688980957
transform -1 0 32384 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp 1688980957
transform -1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1794_
timestamp 1688980957
transform -1 0 29348 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1795_
timestamp 1688980957
transform -1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1796_
timestamp 1688980957
transform -1 0 30912 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1797_
timestamp 1688980957
transform -1 0 31188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1798_
timestamp 1688980957
transform 1 0 29716 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1799_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 1688980957
transform 1 0 27876 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1801_
timestamp 1688980957
transform 1 0 27232 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1802_
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1803_
timestamp 1688980957
transform -1 0 32016 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1804_
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1805_
timestamp 1688980957
transform 1 0 31280 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1806_
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1807_
timestamp 1688980957
transform -1 0 33304 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1808_
timestamp 1688980957
transform 1 0 32752 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1809_
timestamp 1688980957
transform -1 0 34132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1810_
timestamp 1688980957
transform -1 0 28152 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1811_
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1812_
timestamp 1688980957
transform 1 0 33488 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1813_
timestamp 1688980957
transform 1 0 33396 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1814_
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1815_
timestamp 1688980957
transform 1 0 31188 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1816_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1817_
timestamp 1688980957
transform -1 0 33212 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1818_
timestamp 1688980957
transform -1 0 33488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1819_
timestamp 1688980957
transform 1 0 25852 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1820_
timestamp 1688980957
transform 1 0 32200 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1821_
timestamp 1688980957
transform 1 0 35144 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp 1688980957
transform -1 0 33764 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1823_
timestamp 1688980957
transform 1 0 27232 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1824_
timestamp 1688980957
transform 1 0 29072 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1825_
timestamp 1688980957
transform 1 0 30084 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1826_
timestamp 1688980957
transform 1 0 33856 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1827_
timestamp 1688980957
transform 1 0 34408 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1828_
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1829_
timestamp 1688980957
transform 1 0 35052 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1830_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30176 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1831_
timestamp 1688980957
transform 1 0 34408 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1832_
timestamp 1688980957
transform 1 0 35236 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1833_
timestamp 1688980957
transform -1 0 35328 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1834_
timestamp 1688980957
transform -1 0 34500 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1835_
timestamp 1688980957
transform 1 0 33856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1836_
timestamp 1688980957
transform -1 0 33488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1837_
timestamp 1688980957
transform -1 0 34408 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1838_
timestamp 1688980957
transform 1 0 34960 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1839_
timestamp 1688980957
transform 1 0 36156 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1840_
timestamp 1688980957
transform -1 0 33948 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1841_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1842_
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1843_
timestamp 1688980957
transform 1 0 35052 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1844_
timestamp 1688980957
transform 1 0 34040 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1845_
timestamp 1688980957
transform -1 0 30360 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1846_
timestamp 1688980957
transform -1 0 33304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1688980957
transform -1 0 34224 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1848_
timestamp 1688980957
transform 1 0 33304 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1849_
timestamp 1688980957
transform 1 0 34040 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1850_
timestamp 1688980957
transform -1 0 33672 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1851_
timestamp 1688980957
transform 1 0 33396 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1852_
timestamp 1688980957
transform -1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1853_
timestamp 1688980957
transform -1 0 33580 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1854_
timestamp 1688980957
transform -1 0 33856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1855_
timestamp 1688980957
transform 1 0 32844 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1856_
timestamp 1688980957
transform -1 0 33396 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1857_
timestamp 1688980957
transform -1 0 34316 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1858_
timestamp 1688980957
transform -1 0 34040 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1859_
timestamp 1688980957
transform 1 0 32660 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1860_
timestamp 1688980957
transform -1 0 33580 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1861_
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1862_
timestamp 1688980957
transform -1 0 33488 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1863_
timestamp 1688980957
transform 1 0 33304 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1864_
timestamp 1688980957
transform -1 0 31556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1865_
timestamp 1688980957
transform 1 0 31556 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1866_
timestamp 1688980957
transform -1 0 32016 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1867_
timestamp 1688980957
transform 1 0 32200 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1868_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32844 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1869_
timestamp 1688980957
transform 1 0 30544 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1870_
timestamp 1688980957
transform -1 0 24932 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1871_
timestamp 1688980957
transform -1 0 31740 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1872_
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1873_
timestamp 1688980957
transform -1 0 31004 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1874_
timestamp 1688980957
transform 1 0 29624 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1875_
timestamp 1688980957
transform 1 0 32292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_1  _1876_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32752 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1877_
timestamp 1688980957
transform -1 0 31280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1878_
timestamp 1688980957
transform 1 0 29992 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1879_
timestamp 1688980957
transform 1 0 30728 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1880_
timestamp 1688980957
transform -1 0 32568 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1881_
timestamp 1688980957
transform 1 0 32108 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1882_
timestamp 1688980957
transform 1 0 32568 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1883_
timestamp 1688980957
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1884_
timestamp 1688980957
transform -1 0 31648 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1885_
timestamp 1688980957
transform -1 0 31372 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1886_
timestamp 1688980957
transform 1 0 30912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1887_
timestamp 1688980957
transform 1 0 31004 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1888_
timestamp 1688980957
transform -1 0 31924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1889_
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1891_
timestamp 1688980957
transform -1 0 32292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1892_
timestamp 1688980957
transform 1 0 36432 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1893_
timestamp 1688980957
transform -1 0 39560 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1894_
timestamp 1688980957
transform 1 0 38272 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1895_
timestamp 1688980957
transform 1 0 38364 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1896_
timestamp 1688980957
transform 1 0 38732 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1897_
timestamp 1688980957
transform -1 0 38548 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1898_
timestamp 1688980957
transform -1 0 36340 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1899_
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1900_
timestamp 1688980957
transform -1 0 16560 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1901_
timestamp 1688980957
transform 1 0 13524 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1902_
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1903_
timestamp 1688980957
transform 1 0 17112 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1904_
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1905_
timestamp 1688980957
transform -1 0 26772 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1906_
timestamp 1688980957
transform -1 0 25760 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1907_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1908_
timestamp 1688980957
transform 1 0 24656 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1909_
timestamp 1688980957
transform 1 0 19228 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1910_
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1911_
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1912_
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1913_
timestamp 1688980957
transform 1 0 16560 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1914_
timestamp 1688980957
transform -1 0 25116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1915_
timestamp 1688980957
transform -1 0 25668 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1916_
timestamp 1688980957
transform 1 0 17112 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1917_
timestamp 1688980957
transform 1 0 18768 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1918_
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1919_
timestamp 1688980957
transform 1 0 17020 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1920_
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1921_
timestamp 1688980957
transform 1 0 12972 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1922_
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1923_
timestamp 1688980957
transform -1 0 12788 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1924_
timestamp 1688980957
transform 1 0 10948 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1925_
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1926_
timestamp 1688980957
transform -1 0 18400 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1927_
timestamp 1688980957
transform 1 0 12420 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1928_
timestamp 1688980957
transform 1 0 12972 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1929_
timestamp 1688980957
transform 1 0 12880 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1930_
timestamp 1688980957
transform 1 0 14904 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1931_
timestamp 1688980957
transform 1 0 15640 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1932_
timestamp 1688980957
transform 1 0 16652 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1933_
timestamp 1688980957
transform 1 0 17572 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1934_
timestamp 1688980957
transform 1 0 18308 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1935_
timestamp 1688980957
transform 1 0 17940 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1936_
timestamp 1688980957
transform 1 0 20792 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1937_
timestamp 1688980957
transform 1 0 17112 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1938_
timestamp 1688980957
transform 1 0 23460 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1939_
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1940_
timestamp 1688980957
transform 1 0 23736 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1941_
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1942_
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1943_
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1944_
timestamp 1688980957
transform 1 0 29072 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1945_
timestamp 1688980957
transform -1 0 29072 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1946_
timestamp 1688980957
transform 1 0 28336 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1947_
timestamp 1688980957
transform -1 0 29440 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1948_
timestamp 1688980957
transform -1 0 28520 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1949_
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1950_
timestamp 1688980957
transform -1 0 28244 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1951_
timestamp 1688980957
transform -1 0 27968 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1952_
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1953_
timestamp 1688980957
transform -1 0 27600 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1954_
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 1688980957
transform -1 0 27968 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1956_
timestamp 1688980957
transform 1 0 27232 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1957_
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1958_
timestamp 1688980957
transform -1 0 42320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1959_
timestamp 1688980957
transform 1 0 42688 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1960_
timestamp 1688980957
transform -1 0 42320 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1961_
timestamp 1688980957
transform -1 0 43240 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1962_
timestamp 1688980957
transform 1 0 43976 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1963_
timestamp 1688980957
transform -1 0 43240 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1964_
timestamp 1688980957
transform -1 0 43516 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1965_
timestamp 1688980957
transform 1 0 40940 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1966_
timestamp 1688980957
transform -1 0 40480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1967_
timestamp 1688980957
transform 1 0 39008 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1968_
timestamp 1688980957
transform -1 0 39100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1969_
timestamp 1688980957
transform 1 0 37536 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1970_
timestamp 1688980957
transform 1 0 37352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1971_
timestamp 1688980957
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1972_
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1973_
timestamp 1688980957
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1974_
timestamp 1688980957
transform 1 0 36432 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1975_
timestamp 1688980957
transform 1 0 37812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1976_
timestamp 1688980957
transform 1 0 36432 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1977_
timestamp 1688980957
transform -1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1978_
timestamp 1688980957
transform 1 0 37812 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1979_
timestamp 1688980957
transform -1 0 38272 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1980_
timestamp 1688980957
transform 1 0 40572 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1981_
timestamp 1688980957
transform 1 0 41308 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1982_
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1983_
timestamp 1688980957
transform -1 0 41492 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1984_
timestamp 1688980957
transform 1 0 40480 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1985_
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1986_
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1987_
timestamp 1688980957
transform 1 0 36432 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1988_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1989_
timestamp 1688980957
transform 1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1990_
timestamp 1688980957
transform -1 0 22448 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1991_
timestamp 1688980957
transform -1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1992_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1993_
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1994_
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1995_
timestamp 1688980957
transform 1 0 20792 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1996_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1997_
timestamp 1688980957
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1998_
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1999_
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2000_
timestamp 1688980957
transform -1 0 26772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2001_
timestamp 1688980957
transform -1 0 27232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2002_
timestamp 1688980957
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2003_
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2004_
timestamp 1688980957
transform -1 0 23184 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2005_
timestamp 1688980957
transform -1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2006_
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2007_
timestamp 1688980957
transform -1 0 10948 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2008_
timestamp 1688980957
transform 1 0 10488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2009_
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2010_
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2011_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2012_
timestamp 1688980957
transform 1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2013_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2014_
timestamp 1688980957
transform -1 0 13340 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 1688980957
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2016_
timestamp 1688980957
transform -1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2017_
timestamp 1688980957
transform 1 0 22080 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2018_
timestamp 1688980957
transform -1 0 22448 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2019_
timestamp 1688980957
transform -1 0 24840 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2020_
timestamp 1688980957
transform -1 0 24656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2021_
timestamp 1688980957
transform -1 0 24288 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2022_
timestamp 1688980957
transform -1 0 24656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2023_
timestamp 1688980957
transform -1 0 24104 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2024_
timestamp 1688980957
transform 1 0 23552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2025_
timestamp 1688980957
transform -1 0 23644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2026_
timestamp 1688980957
transform -1 0 23368 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2027_
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2028_
timestamp 1688980957
transform -1 0 11316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2029_
timestamp 1688980957
transform -1 0 11132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2030_
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2031_
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2032_
timestamp 1688980957
transform 1 0 11316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2033_
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2034_
timestamp 1688980957
transform 1 0 12052 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2035_
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2036_
timestamp 1688980957
transform 1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2037_
timestamp 1688980957
transform -1 0 15640 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2038_
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _2039_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2040_
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2041_
timestamp 1688980957
transform -1 0 11316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2043_
timestamp 1688980957
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2044_
timestamp 1688980957
transform -1 0 13892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2045_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2047_
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2048_
timestamp 1688980957
transform -1 0 9200 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2049_
timestamp 1688980957
transform -1 0 16928 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _2050_
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2051_
timestamp 1688980957
transform -1 0 15732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2052_
timestamp 1688980957
transform -1 0 18860 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2053_
timestamp 1688980957
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2054_
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2055_
timestamp 1688980957
transform 1 0 14260 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2056_
timestamp 1688980957
transform 1 0 15088 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2057_
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2058_
timestamp 1688980957
transform -1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _2059_
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2060_
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2061_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2062_
timestamp 1688980957
transform 1 0 18032 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2063_
timestamp 1688980957
transform -1 0 18032 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2064_
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2065_
timestamp 1688980957
transform -1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2066_
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2067_
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2068_
timestamp 1688980957
transform 1 0 10396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2069_
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2070_
timestamp 1688980957
transform -1 0 11408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _2071_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _2072_
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2073_
timestamp 1688980957
transform 1 0 31004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2074_
timestamp 1688980957
transform 1 0 31004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2075_
timestamp 1688980957
transform 1 0 30728 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2076_
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _2077_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30544 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__and2b_1  _2078_
timestamp 1688980957
transform -1 0 33212 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2079_
timestamp 1688980957
transform 1 0 31372 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2080_
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2081_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2082_
timestamp 1688980957
transform 1 0 30820 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2083_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_2  _2084_
timestamp 1688980957
transform 1 0 32016 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2085_
timestamp 1688980957
transform -1 0 32384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2086_
timestamp 1688980957
transform -1 0 31464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2087_
timestamp 1688980957
transform -1 0 31832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2088_
timestamp 1688980957
transform -1 0 31372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2089_
timestamp 1688980957
transform -1 0 32016 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2090_
timestamp 1688980957
transform 1 0 29256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2091_
timestamp 1688980957
transform -1 0 31832 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2092_
timestamp 1688980957
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _2093_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30360 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_2  _2094_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _2095_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2096_
timestamp 1688980957
transform -1 0 29532 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2097_
timestamp 1688980957
transform -1 0 30912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2098_
timestamp 1688980957
transform -1 0 29992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2099_
timestamp 1688980957
transform -1 0 29624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2100_
timestamp 1688980957
transform -1 0 31832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _2101_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2102_
timestamp 1688980957
transform -1 0 29992 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2103_
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2104_
timestamp 1688980957
transform 1 0 25852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2105_
timestamp 1688980957
transform 1 0 31280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2106_
timestamp 1688980957
transform 1 0 28980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2107_
timestamp 1688980957
transform -1 0 27784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2108_
timestamp 1688980957
transform -1 0 31372 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2109_
timestamp 1688980957
transform -1 0 28520 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2110_
timestamp 1688980957
transform 1 0 27784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2111_
timestamp 1688980957
transform -1 0 30544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2112_
timestamp 1688980957
transform 1 0 28704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _2113_
timestamp 1688980957
transform -1 0 28428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2114_
timestamp 1688980957
transform 1 0 26496 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2115_
timestamp 1688980957
transform -1 0 24288 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2116_
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2117_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _2118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2119_
timestamp 1688980957
transform -1 0 31648 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2120_
timestamp 1688980957
transform -1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2122_
timestamp 1688980957
transform -1 0 30360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2123_
timestamp 1688980957
transform 1 0 30084 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2124_
timestamp 1688980957
transform -1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2125_
timestamp 1688980957
transform -1 0 31004 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2126_
timestamp 1688980957
transform 1 0 25300 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2127_
timestamp 1688980957
transform -1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2128_
timestamp 1688980957
transform -1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2129_
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2130_
timestamp 1688980957
transform -1 0 28888 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _2131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28244 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2132_
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2133_
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2134_
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2135_
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2136_
timestamp 1688980957
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2137_
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2138_
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2139_
timestamp 1688980957
transform -1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _2140_
timestamp 1688980957
transform 1 0 15640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2141_
timestamp 1688980957
transform -1 0 18400 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2142_
timestamp 1688980957
transform -1 0 15640 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _2143_
timestamp 1688980957
transform 1 0 14720 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2144_
timestamp 1688980957
transform 1 0 11316 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2145_
timestamp 1688980957
transform 1 0 15364 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2146_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2147_
timestamp 1688980957
transform -1 0 17572 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _2148_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _2149_
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2150_
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2151_
timestamp 1688980957
transform -1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2152_
timestamp 1688980957
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2153_
timestamp 1688980957
transform -1 0 18308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2154_
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2155_
timestamp 1688980957
transform -1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2156_
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2157_
timestamp 1688980957
transform -1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2158_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__a31o_1  _2159_
timestamp 1688980957
transform 1 0 29624 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2160_
timestamp 1688980957
transform -1 0 28888 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2161_
timestamp 1688980957
transform 1 0 25668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2162_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2163_
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2164_
timestamp 1688980957
transform -1 0 22172 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _2165_
timestamp 1688980957
transform -1 0 27784 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  _2166_
timestamp 1688980957
transform -1 0 22816 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2167_
timestamp 1688980957
transform -1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2168_
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2169_
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2170_
timestamp 1688980957
transform 1 0 20976 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2171_
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2172_
timestamp 1688980957
transform -1 0 28244 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2173_
timestamp 1688980957
transform 1 0 25668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2174_
timestamp 1688980957
transform 1 0 24288 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2175_
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2176_
timestamp 1688980957
transform 1 0 23184 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2177_
timestamp 1688980957
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2178_
timestamp 1688980957
transform -1 0 19136 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2179_
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2180_
timestamp 1688980957
transform -1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2181_
timestamp 1688980957
transform -1 0 19044 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2182_
timestamp 1688980957
transform -1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2183_
timestamp 1688980957
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2184_
timestamp 1688980957
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2185_
timestamp 1688980957
transform -1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2186_
timestamp 1688980957
transform -1 0 18768 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _2187_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2188_
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2189_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2190_
timestamp 1688980957
transform 1 0 17112 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2191_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2192_
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2193_
timestamp 1688980957
transform -1 0 28704 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2194_
timestamp 1688980957
transform 1 0 25760 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2195_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2196_
timestamp 1688980957
transform 1 0 25024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2197_
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2198_
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2199_
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2200_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2201_
timestamp 1688980957
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2202_
timestamp 1688980957
transform -1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _2203_
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2204_
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _2205_
timestamp 1688980957
transform -1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2206_
timestamp 1688980957
transform -1 0 17480 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _2207_
timestamp 1688980957
transform 1 0 16376 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _2208_
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2209_
timestamp 1688980957
transform -1 0 21712 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2210_
timestamp 1688980957
transform 1 0 20884 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2211_
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2212_
timestamp 1688980957
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _2213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2214_
timestamp 1688980957
transform -1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2215_
timestamp 1688980957
transform -1 0 19780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2216_
timestamp 1688980957
transform 1 0 10120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2217_
timestamp 1688980957
transform 1 0 19228 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2218_
timestamp 1688980957
transform -1 0 20148 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2219_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2220_
timestamp 1688980957
transform -1 0 13984 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2221_
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2222_
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _2223_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2224_
timestamp 1688980957
transform 1 0 10488 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2225_
timestamp 1688980957
transform -1 0 14076 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2226_
timestamp 1688980957
transform 1 0 28704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2227_
timestamp 1688980957
transform 1 0 28428 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2228_
timestamp 1688980957
transform -1 0 28428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2229_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2230_
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2231_
timestamp 1688980957
transform -1 0 21712 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2232_
timestamp 1688980957
transform -1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2233_
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2234_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2235_
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2236_
timestamp 1688980957
transform 1 0 15824 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2237_
timestamp 1688980957
transform 1 0 15088 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2238_
timestamp 1688980957
transform -1 0 16376 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2239_
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2240_
timestamp 1688980957
transform 1 0 16928 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2241_
timestamp 1688980957
transform -1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2242_
timestamp 1688980957
transform -1 0 16928 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2243_
timestamp 1688980957
transform 1 0 10304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2244_
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2245_
timestamp 1688980957
transform -1 0 16468 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2246_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2247_
timestamp 1688980957
transform -1 0 16560 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2248_
timestamp 1688980957
transform -1 0 22908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2249_
timestamp 1688980957
transform 1 0 26036 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2250_
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2251_
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2252_
timestamp 1688980957
transform -1 0 22632 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2253_
timestamp 1688980957
transform 1 0 22356 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2254_
timestamp 1688980957
transform -1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2255_
timestamp 1688980957
transform 1 0 31004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2256_
timestamp 1688980957
transform 1 0 29624 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2257_
timestamp 1688980957
transform -1 0 29992 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2258_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2259_
timestamp 1688980957
transform -1 0 25116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2260_
timestamp 1688980957
transform 1 0 24472 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2261_
timestamp 1688980957
transform 1 0 23920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2262_
timestamp 1688980957
transform -1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2263_
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2264_
timestamp 1688980957
transform 1 0 14628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2265_
timestamp 1688980957
transform -1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2266_
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2267_
timestamp 1688980957
transform 1 0 9844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _2268_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2269_
timestamp 1688980957
transform -1 0 17204 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2270_
timestamp 1688980957
transform -1 0 19136 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2271_
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2272_
timestamp 1688980957
transform -1 0 18584 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2273_
timestamp 1688980957
transform 1 0 17940 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2274_
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2275_
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2276_
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _2277_
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2278_
timestamp 1688980957
transform -1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _2279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2280_
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2281_
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2282_
timestamp 1688980957
transform -1 0 13340 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2283_
timestamp 1688980957
transform 1 0 12328 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__a311o_1  _2284_
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2285_
timestamp 1688980957
transform 1 0 27508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2286_
timestamp 1688980957
transform -1 0 28336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2287_
timestamp 1688980957
transform 1 0 25484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2288_
timestamp 1688980957
transform -1 0 22632 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2289_
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2290_
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2291_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2292_
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2293_
timestamp 1688980957
transform -1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2294_
timestamp 1688980957
transform 1 0 14076 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2295_
timestamp 1688980957
transform 1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2296_
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2297_
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2298_
timestamp 1688980957
transform 1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2299_
timestamp 1688980957
transform -1 0 14628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2300_
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2301_
timestamp 1688980957
transform 1 0 15180 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2302_
timestamp 1688980957
transform -1 0 13432 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _2303_
timestamp 1688980957
transform 1 0 13432 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _2304_
timestamp 1688980957
transform -1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2305_
timestamp 1688980957
transform 1 0 27876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2306_
timestamp 1688980957
transform 1 0 26680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2307_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2308_
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2309_
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2310_
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2311_
timestamp 1688980957
transform -1 0 21804 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2312_
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2313_
timestamp 1688980957
transform -1 0 11408 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2314_
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2315_
timestamp 1688980957
transform 1 0 10580 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2316_
timestamp 1688980957
transform -1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2317_
timestamp 1688980957
transform -1 0 11408 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2318_
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2319_
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2320_
timestamp 1688980957
transform -1 0 11132 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2321_
timestamp 1688980957
transform -1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2322_
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _2323_
timestamp 1688980957
transform -1 0 12604 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2324_
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2325_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29256 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2326_
timestamp 1688980957
transform -1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2327_
timestamp 1688980957
transform 1 0 25852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2328_
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _2329_
timestamp 1688980957
transform -1 0 11868 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2330_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2331_
timestamp 1688980957
transform 1 0 10672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2332_
timestamp 1688980957
transform 1 0 23276 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2333_
timestamp 1688980957
transform 1 0 23920 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2334_
timestamp 1688980957
transform 1 0 22816 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2335_
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2336_
timestamp 1688980957
transform -1 0 11040 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2337_
timestamp 1688980957
transform 1 0 11868 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2338_
timestamp 1688980957
transform -1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2339_
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2340_
timestamp 1688980957
transform -1 0 13984 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2341_
timestamp 1688980957
transform 1 0 12880 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2342_
timestamp 1688980957
transform -1 0 12788 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2343_
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2344_
timestamp 1688980957
transform 1 0 12696 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2345_
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2346_
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2347_
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2348_
timestamp 1688980957
transform -1 0 11776 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2349_
timestamp 1688980957
transform -1 0 11316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2350_
timestamp 1688980957
transform -1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2351_
timestamp 1688980957
transform 1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2352_
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2353_
timestamp 1688980957
transform -1 0 11408 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__or3_1  _2354_
timestamp 1688980957
transform 1 0 26404 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2355_
timestamp 1688980957
transform -1 0 27324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2356_
timestamp 1688980957
transform -1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2357_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2358_
timestamp 1688980957
transform 1 0 11960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2359_
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2360_
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2361_
timestamp 1688980957
transform 1 0 12328 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _2362_
timestamp 1688980957
transform 1 0 12972 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2363_
timestamp 1688980957
transform -1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2364_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2365_
timestamp 1688980957
transform -1 0 13800 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2366_
timestamp 1688980957
transform -1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2367_
timestamp 1688980957
transform 1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2368_
timestamp 1688980957
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2369_
timestamp 1688980957
transform 1 0 21988 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2370_
timestamp 1688980957
transform 1 0 22080 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2371_
timestamp 1688980957
transform -1 0 14628 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2372_
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2373_
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2374_
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2375_
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2376_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _2377_
timestamp 1688980957
transform -1 0 12052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2378_
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2379_
timestamp 1688980957
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2380_
timestamp 1688980957
transform -1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2381_
timestamp 1688980957
transform -1 0 16376 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2382_
timestamp 1688980957
transform -1 0 16744 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2383_
timestamp 1688980957
transform 1 0 15548 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2384_
timestamp 1688980957
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2385_
timestamp 1688980957
transform -1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2386_
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2387_
timestamp 1688980957
transform -1 0 17204 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2388_
timestamp 1688980957
transform -1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _2389_
timestamp 1688980957
transform -1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2390_
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2391_
timestamp 1688980957
transform -1 0 22816 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2392_
timestamp 1688980957
transform 1 0 21896 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2393_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2394_
timestamp 1688980957
transform -1 0 19872 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2395_
timestamp 1688980957
transform -1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2396_
timestamp 1688980957
transform -1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2397_
timestamp 1688980957
transform -1 0 19228 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2398_
timestamp 1688980957
transform -1 0 23552 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 1688980957
transform 1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2400_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2401_
timestamp 1688980957
transform -1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2402_
timestamp 1688980957
transform -1 0 18676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 1688980957
transform -1 0 20056 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2404_
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2405_
timestamp 1688980957
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2406_
timestamp 1688980957
transform 1 0 23276 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2407_
timestamp 1688980957
transform 1 0 23000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2408_
timestamp 1688980957
transform 1 0 22448 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2409_
timestamp 1688980957
transform -1 0 22448 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2410_
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _2411_
timestamp 1688980957
transform -1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2412_
timestamp 1688980957
transform -1 0 22172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2413_
timestamp 1688980957
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2414_
timestamp 1688980957
transform 1 0 14536 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2415_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2416_
timestamp 1688980957
transform 1 0 21160 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2417_
timestamp 1688980957
transform 1 0 20792 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2418_
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2419_
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2420_
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2421_
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2422_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2423_
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2424_
timestamp 1688980957
transform 1 0 16928 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2425_
timestamp 1688980957
transform 1 0 17572 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2426_
timestamp 1688980957
transform -1 0 16560 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2427_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2428_
timestamp 1688980957
transform 1 0 18124 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2429_
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2430_
timestamp 1688980957
transform 1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2431_
timestamp 1688980957
transform -1 0 19596 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2432_
timestamp 1688980957
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2433_
timestamp 1688980957
transform 1 0 10948 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2434_
timestamp 1688980957
transform 1 0 10580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2435_
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2436_
timestamp 1688980957
transform 1 0 12052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2437_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2438_
timestamp 1688980957
transform 1 0 10304 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2439_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2440_
timestamp 1688980957
transform -1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2441_
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2442_
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2443_
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2444_
timestamp 1688980957
transform -1 0 16928 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2445_
timestamp 1688980957
transform -1 0 17572 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2446_
timestamp 1688980957
transform 1 0 23460 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2447_
timestamp 1688980957
transform -1 0 22632 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2448_
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2449_
timestamp 1688980957
transform -1 0 24288 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2450_
timestamp 1688980957
transform 1 0 22632 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2451_
timestamp 1688980957
transform -1 0 22356 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2452_
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2453_
timestamp 1688980957
transform 1 0 17112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2454_
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2455_
timestamp 1688980957
transform 1 0 23552 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2456_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2457_
timestamp 1688980957
transform 1 0 23552 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2458_
timestamp 1688980957
transform 1 0 18308 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2459_
timestamp 1688980957
transform -1 0 17296 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2460_
timestamp 1688980957
transform 1 0 12972 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2461_
timestamp 1688980957
transform 1 0 9384 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2462_
timestamp 1688980957
transform -1 0 10212 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2463_
timestamp 1688980957
transform -1 0 11408 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2464_
timestamp 1688980957
transform 1 0 13432 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2465_
timestamp 1688980957
transform 1 0 17480 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2466_
timestamp 1688980957
transform 1 0 18584 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2467_
timestamp 1688980957
transform 1 0 19136 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2468_
timestamp 1688980957
transform -1 0 22356 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2469_
timestamp 1688980957
transform 1 0 22080 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2470_
timestamp 1688980957
transform 1 0 12328 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2471_
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2472_
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2473_
timestamp 1688980957
transform -1 0 14352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2474_
timestamp 1688980957
transform 1 0 14444 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2475_
timestamp 1688980957
transform -1 0 13984 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2476_
timestamp 1688980957
transform 1 0 16744 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2477_
timestamp 1688980957
transform -1 0 16560 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2478_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2479_
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2480_
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2481_
timestamp 1688980957
transform 1 0 14720 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2482_
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2483_
timestamp 1688980957
transform 1 0 15824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2484_
timestamp 1688980957
transform -1 0 16560 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2485_
timestamp 1688980957
transform -1 0 15272 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2486_
timestamp 1688980957
transform 1 0 15272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2487_
timestamp 1688980957
transform 1 0 7636 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2488_
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2489_
timestamp 1688980957
transform 1 0 7636 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2490_
timestamp 1688980957
transform 1 0 7084 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2491_
timestamp 1688980957
transform 1 0 8648 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2492_
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2493_
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2494_
timestamp 1688980957
transform 1 0 10948 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2495_
timestamp 1688980957
transform -1 0 10212 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2496_
timestamp 1688980957
transform 1 0 9660 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2497_
timestamp 1688980957
transform 1 0 8004 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2498_
timestamp 1688980957
transform 1 0 7728 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2499_
timestamp 1688980957
transform -1 0 16100 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2500_
timestamp 1688980957
transform 1 0 16100 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2501_
timestamp 1688980957
transform -1 0 17112 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2502_
timestamp 1688980957
transform 1 0 17848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 1688980957
transform 1 0 15732 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2504_
timestamp 1688980957
transform -1 0 13984 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2505_
timestamp 1688980957
transform -1 0 23552 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 1688980957
transform 1 0 14996 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2507_
timestamp 1688980957
transform -1 0 14904 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 1688980957
transform -1 0 20884 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2509_
timestamp 1688980957
transform 1 0 21252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 17664 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2511_
timestamp 1688980957
transform -1 0 17112 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2512_
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2513_
timestamp 1688980957
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2514_
timestamp 1688980957
transform -1 0 23184 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2515_
timestamp 1688980957
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2516_
timestamp 1688980957
transform -1 0 18400 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2517_
timestamp 1688980957
transform 1 0 18032 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform 1 0 22172 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2519_
timestamp 1688980957
transform -1 0 21712 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2521_
timestamp 1688980957
transform -1 0 19136 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 1688980957
transform -1 0 20332 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2523_
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2524_
timestamp 1688980957
transform 1 0 13064 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2525_
timestamp 1688980957
transform 1 0 12512 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2526_
timestamp 1688980957
transform 1 0 10672 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2527_
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2528_
timestamp 1688980957
transform 1 0 10488 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2529_
timestamp 1688980957
transform 1 0 10028 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2530_
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2531_
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2532_
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2533_
timestamp 1688980957
transform 1 0 13432 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2534_
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2535_
timestamp 1688980957
transform -1 0 16100 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2536_
timestamp 1688980957
transform 1 0 19964 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2537_
timestamp 1688980957
transform -1 0 18400 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 19504 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 1688980957
transform -1 0 19136 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2541_
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2543_
timestamp 1688980957
transform 1 0 21160 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2544_
timestamp 1688980957
transform 1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2545_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2546_
timestamp 1688980957
transform -1 0 8280 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _2547_
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2548_
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2549_
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2550_
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2551_
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2552_
timestamp 1688980957
transform -1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2553_
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2554_
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2555_
timestamp 1688980957
transform -1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2556_
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 1688980957
transform -1 0 7912 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2558_
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2559_
timestamp 1688980957
transform -1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2560_
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2561_
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2562_
timestamp 1688980957
transform -1 0 8556 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2563_
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2564_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34776 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2565_
timestamp 1688980957
transform -1 0 39284 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2566_
timestamp 1688980957
transform 1 0 35328 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2567_
timestamp 1688980957
transform 1 0 35052 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2568_
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2569_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2570_
timestamp 1688980957
transform -1 0 36524 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2571_
timestamp 1688980957
transform 1 0 35052 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2572_
timestamp 1688980957
transform -1 0 40480 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2573_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37812 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2574_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7268 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2575_
timestamp 1688980957
transform -1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2576_
timestamp 1688980957
transform 1 0 3312 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2577_
timestamp 1688980957
transform -1 0 6164 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2578_
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2579_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2580_
timestamp 1688980957
transform -1 0 8556 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2581_
timestamp 1688980957
transform 1 0 7636 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2582_
timestamp 1688980957
transform -1 0 10764 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2583_
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2584_
timestamp 1688980957
transform -1 0 8924 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2585_
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2586_
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2587_
timestamp 1688980957
transform -1 0 5888 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2588_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2589_
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2590_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _2591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2592_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2593_
timestamp 1688980957
transform 1 0 32660 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2594_
timestamp 1688980957
transform 1 0 34684 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2595_
timestamp 1688980957
transform 1 0 35328 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2596_
timestamp 1688980957
transform 1 0 34224 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2597_
timestamp 1688980957
transform 1 0 34960 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2598_
timestamp 1688980957
transform 1 0 35052 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2599_
timestamp 1688980957
transform 1 0 37076 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2600_
timestamp 1688980957
transform -1 0 39100 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2602_
timestamp 1688980957
transform 1 0 38456 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2604_
timestamp 1688980957
transform 1 0 38916 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2605_
timestamp 1688980957
transform 1 0 39836 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2606_
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2607_
timestamp 1688980957
transform 1 0 42504 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2608_
timestamp 1688980957
transform -1 0 44252 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2609_
timestamp 1688980957
transform 1 0 37812 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 1688980957
transform 1 0 39376 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2611_
timestamp 1688980957
transform 1 0 39284 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 1688980957
transform -1 0 44252 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 1688980957
transform -1 0 44344 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 1688980957
transform -1 0 44344 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2617_
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2618_
timestamp 1688980957
transform -1 0 34592 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2619_
timestamp 1688980957
transform 1 0 32384 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2620_
timestamp 1688980957
transform 1 0 32752 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2621_
timestamp 1688980957
transform 1 0 32844 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2622_
timestamp 1688980957
transform -1 0 38364 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2623_
timestamp 1688980957
transform 1 0 28520 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2624_
timestamp 1688980957
transform -1 0 32476 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2625_
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2626_
timestamp 1688980957
transform 1 0 28888 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2627_
timestamp 1688980957
transform -1 0 38088 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2628_
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2629_
timestamp 1688980957
transform -1 0 34040 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2630_
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2631_
timestamp 1688980957
transform 1 0 8924 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2632_
timestamp 1688980957
transform 1 0 27416 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2633_
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2634_
timestamp 1688980957
transform 1 0 8280 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2635_
timestamp 1688980957
transform 1 0 20148 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2636_
timestamp 1688980957
transform -1 0 39468 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2637_
timestamp 1688980957
transform 1 0 32200 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2638_
timestamp 1688980957
transform -1 0 44344 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2639_
timestamp 1688980957
transform 1 0 36064 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2640_
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2641_
timestamp 1688980957
transform -1 0 37168 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2642_
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 1688980957
transform 1 0 19872 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2644_
timestamp 1688980957
transform -1 0 37168 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2645_
timestamp 1688980957
transform 1 0 6716 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2646_
timestamp 1688980957
transform 1 0 31280 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 1688980957
transform 1 0 26956 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 1688980957
transform 1 0 5796 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2649_
timestamp 1688980957
transform 1 0 25024 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2650_
timestamp 1688980957
transform 1 0 2760 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2651_
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2652_
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2653_
timestamp 1688980957
transform -1 0 44344 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2654_
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2655_
timestamp 1688980957
transform 1 0 42504 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2656_
timestamp 1688980957
transform 1 0 40480 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 1688980957
transform 1 0 32752 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2658_
timestamp 1688980957
transform -1 0 37168 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 1688980957
transform 1 0 34868 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 1688980957
transform -1 0 36156 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2661_
timestamp 1688980957
transform 1 0 32752 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2662_
timestamp 1688980957
transform -1 0 32384 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2663_
timestamp 1688980957
transform 1 0 27600 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 1688980957
transform 1 0 30820 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2665_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2666_
timestamp 1688980957
transform -1 0 28612 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2667_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2668_
timestamp 1688980957
transform -1 0 33948 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2669_
timestamp 1688980957
transform -1 0 28796 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2670_
timestamp 1688980957
transform -1 0 33948 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2671_
timestamp 1688980957
transform 1 0 28612 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2672_
timestamp 1688980957
transform 1 0 33304 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2673_
timestamp 1688980957
transform 1 0 31280 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2674_
timestamp 1688980957
transform 1 0 35512 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2675_
timestamp 1688980957
transform -1 0 39100 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2676_
timestamp 1688980957
transform -1 0 36432 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2677_
timestamp 1688980957
transform 1 0 32108 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2678_
timestamp 1688980957
transform -1 0 32108 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2679_
timestamp 1688980957
transform 1 0 29624 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2680_
timestamp 1688980957
transform 1 0 28612 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2681_
timestamp 1688980957
transform 1 0 29256 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2682_
timestamp 1688980957
transform 1 0 28244 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 37076 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 38456 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 1688980957
transform 1 0 38732 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 1688980957
transform -1 0 40756 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform -1 0 40940 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 35604 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 1688980957
transform 1 0 34868 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2691_
timestamp 1688980957
transform 1 0 27508 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 1688980957
transform -1 0 27508 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 24840 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform -1 0 26404 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform 1 0 24196 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 1688980957
transform -1 0 25668 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2697_
timestamp 1688980957
transform -1 0 20424 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 1688980957
transform -1 0 18308 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 1688980957
transform -1 0 14628 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 1688980957
transform 1 0 11500 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 1688980957
transform -1 0 13708 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 13064 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2703_
timestamp 1688980957
transform 1 0 14904 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2704_
timestamp 1688980957
transform -1 0 18676 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2705_
timestamp 1688980957
transform 1 0 19044 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2706_
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 1688980957
transform 1 0 24472 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 1688980957
transform 1 0 33488 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2710_
timestamp 1688980957
transform 1 0 26404 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2711_
timestamp 1688980957
transform 1 0 27968 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2712_
timestamp 1688980957
transform 1 0 26036 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 1688980957
transform 1 0 26220 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2714_
timestamp 1688980957
transform 1 0 26680 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2715_
timestamp 1688980957
transform 1 0 42044 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2716_
timestamp 1688980957
transform 1 0 42228 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2717_
timestamp 1688980957
transform -1 0 44344 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2718_
timestamp 1688980957
transform -1 0 44252 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2719_
timestamp 1688980957
transform 1 0 40480 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 1688980957
transform 1 0 39100 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 1688980957
transform 1 0 36984 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2722_
timestamp 1688980957
transform 1 0 36156 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 1688980957
transform 1 0 40296 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 1688980957
transform 1 0 40848 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 1688980957
transform 1 0 40388 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 1688980957
transform 1 0 41676 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 1688980957
transform 1 0 38088 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 1688980957
transform 1 0 36340 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 1688980957
transform 1 0 35328 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 1688980957
transform 1 0 35880 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 1688980957
transform 1 0 42320 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 1688980957
transform 1 0 42504 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 1688980957
transform 1 0 42504 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2736_
timestamp 1688980957
transform 1 0 40940 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2737_
timestamp 1688980957
transform 1 0 39928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2738_
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2739_
timestamp 1688980957
transform 1 0 36984 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2740_
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _2741_
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2742_
timestamp 1688980957
transform -1 0 11040 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2743_
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2744_
timestamp 1688980957
transform 1 0 9292 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2745_
timestamp 1688980957
transform 1 0 6624 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2746_
timestamp 1688980957
transform 1 0 4692 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2747_
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2748_
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2749_
timestamp 1688980957
transform 1 0 5428 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2750_
timestamp 1688980957
transform 1 0 7728 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2751_
timestamp 1688980957
transform 1 0 6900 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2752_
timestamp 1688980957
transform 1 0 9292 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2753_
timestamp 1688980957
transform 1 0 3864 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2754_
timestamp 1688980957
transform 1 0 4324 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2755_
timestamp 1688980957
transform 1 0 5704 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2756_
timestamp 1688980957
transform 1 0 6900 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 1688980957
transform 1 0 9660 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 1688980957
transform 1 0 9016 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2759_
timestamp 1688980957
transform 1 0 17848 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2760_
timestamp 1688980957
transform 1 0 22540 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2761_
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2762_
timestamp 1688980957
transform 1 0 20516 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2763_
timestamp 1688980957
transform 1 0 18400 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2764_
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2765_
timestamp 1688980957
transform -1 0 27876 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2766_
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2767_
timestamp 1688980957
transform -1 0 25116 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2768_
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2769_
timestamp 1688980957
transform 1 0 12420 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2770_
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2771_
timestamp 1688980957
transform 1 0 13340 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2772_
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2773_
timestamp 1688980957
transform 1 0 22448 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2774_
timestamp 1688980957
transform 1 0 24656 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2775_
timestamp 1688980957
transform 1 0 25024 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2776_
timestamp 1688980957
transform 1 0 23368 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 1688980957
transform 1 0 17296 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 1688980957
transform 1 0 15916 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 1688980957
transform 1 0 20056 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 1688980957
transform 1 0 17848 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 1688980957
transform 1 0 24932 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 1688980957
transform 1 0 13248 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2785_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2786_
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2787_
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2788_
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2789_
timestamp 1688980957
transform 1 0 12144 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2790_
timestamp 1688980957
transform 1 0 14720 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2791_
timestamp 1688980957
transform 1 0 20976 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2792_
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 1688980957
transform 1 0 13524 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 1688980957
transform 1 0 19872 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2797_
timestamp 1688980957
transform 1 0 15364 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2798_
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2799_
timestamp 1688980957
transform 1 0 17940 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 1688980957
transform 1 0 11868 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2803_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 1688980957
transform 1 0 9844 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2806_
timestamp 1688980957
transform 1 0 9476 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2807_
timestamp 1688980957
transform 1 0 11040 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2808_
timestamp 1688980957
transform 1 0 13800 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2810_
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2811_
timestamp 1688980957
transform 1 0 24104 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2812_
timestamp 1688980957
transform 1 0 22172 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2813_
timestamp 1688980957
transform 1 0 19320 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2814_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2815_
timestamp 1688980957
transform -1 0 23644 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2816_
timestamp 1688980957
transform -1 0 23828 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2817_
timestamp 1688980957
transform 1 0 15732 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2818_
timestamp 1688980957
transform -1 0 23552 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2819_
timestamp 1688980957
transform 1 0 17020 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2820_
timestamp 1688980957
transform 1 0 17020 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2821_
timestamp 1688980957
transform -1 0 14076 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2822_
timestamp 1688980957
transform 1 0 9384 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2823_
timestamp 1688980957
transform 1 0 9108 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2824_
timestamp 1688980957
transform 1 0 10580 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2825_
timestamp 1688980957
transform 1 0 12696 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2826_
timestamp 1688980957
transform 1 0 15272 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2827_
timestamp 1688980957
transform 1 0 18124 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2828_
timestamp 1688980957
transform 1 0 18492 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2829_
timestamp 1688980957
transform -1 0 24012 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2830_
timestamp 1688980957
transform 1 0 21804 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2831_
timestamp 1688980957
transform 1 0 11592 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2832_
timestamp 1688980957
transform 1 0 14076 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2833_
timestamp 1688980957
transform 1 0 13984 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2834_
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2835_
timestamp 1688980957
transform 1 0 10672 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2836_
timestamp 1688980957
transform 1 0 14444 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2837_
timestamp 1688980957
transform 1 0 15640 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2838_
timestamp 1688980957
transform 1 0 14260 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2839_
timestamp 1688980957
transform 1 0 6532 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2840_
timestamp 1688980957
transform 1 0 6440 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2841_
timestamp 1688980957
transform 1 0 6808 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2842_
timestamp 1688980957
transform 1 0 10212 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2843_
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2844_
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2845_
timestamp 1688980957
transform 1 0 15272 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2846_
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2847_
timestamp 1688980957
transform 1 0 14260 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2848_
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2849_
timestamp 1688980957
transform -1 0 21252 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2850_
timestamp 1688980957
transform 1 0 17112 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2851_
timestamp 1688980957
transform 1 0 21620 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2852_
timestamp 1688980957
transform -1 0 23644 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2853_
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2854_
timestamp 1688980957
transform -1 0 23644 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2855_
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2856_
timestamp 1688980957
transform -1 0 21068 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2857_
timestamp 1688980957
transform 1 0 11776 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2858_
timestamp 1688980957
transform 1 0 9568 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2859_
timestamp 1688980957
transform 1 0 9568 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2860_
timestamp 1688980957
transform 1 0 10212 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2861_
timestamp 1688980957
transform 1 0 13064 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2862_
timestamp 1688980957
transform 1 0 16100 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2863_
timestamp 1688980957
transform 1 0 19228 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2864_
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2865_
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2866_
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2867_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2868_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _2869_
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2870_
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2871_
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2872_
timestamp 1688980957
transform 1 0 7912 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2873_
timestamp 1688980957
transform 1 0 41308 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26496 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform -1 0 33028 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform -1 0 14812 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 33764 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1688980957
transform 1 0 10948 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1688980957
transform -1 0 18860 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1688980957
transform -1 0 18032 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1688980957
transform -1 0 11224 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1688980957
transform -1 0 8188 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1688980957
transform 1 0 6900 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1688980957
transform 1 0 9108 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1688980957
transform 1 0 13892 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1688980957
transform -1 0 21068 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1688980957
transform -1 0 17480 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1688980957
transform 1 0 23000 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1688980957
transform 1 0 27140 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1688980957
transform -1 0 27232 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1688980957
transform -1 0 32660 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1688980957
transform -1 0 38272 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1688980957
transform 1 0 42504 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1688980957
transform 1 0 42504 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1688980957
transform -1 0 32016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1688980957
transform 1 0 35144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1688980957
transform -1 0 39100 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1688980957
transform 1 0 40480 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1688980957
transform 1 0 37904 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1688980957
transform 1 0 42504 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1688980957
transform -1 0 37168 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_clk
timestamp 1688980957
transform -1 0 34684 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1688980957
transform -1 0 28796 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1688980957
transform 1 0 18124 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1688980957
transform -1 0 21712 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1688980957
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1688980957
transform -1 0 7268 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_37_clk
timestamp 1688980957
transform -1 0 8188 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1688980957
transform -1 0 7268 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1688980957
transform 1 0 7268 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1688980957
transform -1 0 7544 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1688980957
transform 1 0 6440 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 1688980957
transform -1 0 16560 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1688980957
transform 1 0 15364 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1688980957
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1688980957
transform 1 0 35236 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1688980957
transform 1 0 35696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 1688980957
transform 1 0 28612 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1688980957
transform 1 0 36156 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1688980957
transform -1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1688980957
transform -1 0 8004 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1688980957
transform -1 0 6992 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1688980957
transform -1 0 16376 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1688980957
transform -1 0 18032 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1688980957
transform 1 0 6992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1688980957
transform 1 0 9200 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1688980957
transform -1 0 8464 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1688980957
transform -1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1688980957
transform -1 0 14628 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1688980957
transform 1 0 19320 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1688980957
transform 1 0 8464 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1688980957
transform -1 0 31004 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1688980957
transform -1 0 26772 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1688980957
transform -1 0 35696 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1688980957
transform -1 0 39652 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1688980957
transform 1 0 37536 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1688980957
transform 1 0 37444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1688980957
transform -1 0 26864 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1688980957
transform 1 0 36616 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 1688980957
transform -1 0 35236 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1688980957
transform -1 0 35420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1688980957
transform 1 0 27324 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_197 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_211
timestamp 1688980957
transform 1 0 20516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_275 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_469
timestamp 1688980957
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_129
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_141
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_154
timestamp 1688980957
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_160
timestamp 1688980957
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_178
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_190
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_197
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp 1688980957
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 1688980957
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_239
timestamp 1688980957
transform 1 0 23092 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_247
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1688980957
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_297
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_318
timestamp 1688980957
transform 1 0 30360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_330
timestamp 1688980957
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_379
timestamp 1688980957
transform 1 0 35972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_386
timestamp 1688980957
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_469
timestamp 1688980957
transform 1 0 44252 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_116
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_154
timestamp 1688980957
transform 1 0 15272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_160
timestamp 1688980957
transform 1 0 15824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_192
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_200
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_208
timestamp 1688980957
transform 1 0 20240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_243
timestamp 1688980957
transform 1 0 23460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_273
timestamp 1688980957
transform 1 0 26220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_383
timestamp 1688980957
transform 1 0 36340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_395
timestamp 1688980957
transform 1 0 37444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_407
timestamp 1688980957
transform 1 0 38548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_63
timestamp 1688980957
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_85
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_102
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_120
timestamp 1688980957
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_196
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_238
timestamp 1688980957
transform 1 0 23000 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_259
timestamp 1688980957
transform 1 0 24932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_271
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_301
timestamp 1688980957
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_325
timestamp 1688980957
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_369
timestamp 1688980957
transform 1 0 35052 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_469
timestamp 1688980957
transform 1 0 44252 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_61
timestamp 1688980957
transform 1 0 6716 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_67
timestamp 1688980957
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_117
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_124
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_162
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_174
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_186
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_205
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_217
timestamp 1688980957
transform 1 0 21068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_229
timestamp 1688980957
transform 1 0 22172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_241
timestamp 1688980957
transform 1 0 23276 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp 1688980957
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_276
timestamp 1688980957
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_341
timestamp 1688980957
transform 1 0 32476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_347
timestamp 1688980957
transform 1 0 33028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_371
timestamp 1688980957
transform 1 0 35236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_383
timestamp 1688980957
transform 1 0 36340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_395
timestamp 1688980957
transform 1 0 37444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_407
timestamp 1688980957
transform 1 0 38548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_78
timestamp 1688980957
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_88
timestamp 1688980957
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_99
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_118
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_126
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_134
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_153
timestamp 1688980957
transform 1 0 15180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_234
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_246
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_258
timestamp 1688980957
transform 1 0 24840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_266
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_304
timestamp 1688980957
transform 1 0 29072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_316
timestamp 1688980957
transform 1 0 30176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_324
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_334
timestamp 1688980957
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_340
timestamp 1688980957
transform 1 0 32384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_344
timestamp 1688980957
transform 1 0 32752 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_365
timestamp 1688980957
transform 1 0 34684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_377
timestamp 1688980957
transform 1 0 35788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_389
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_469
timestamp 1688980957
transform 1 0 44252 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_159
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_168
timestamp 1688980957
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_180
timestamp 1688980957
transform 1 0 17664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_188
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_203
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_237
timestamp 1688980957
transform 1 0 22908 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_266
timestamp 1688980957
transform 1 0 25576 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_278
timestamp 1688980957
transform 1 0 26680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_290
timestamp 1688980957
transform 1 0 27784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_302
timestamp 1688980957
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_339
timestamp 1688980957
transform 1 0 32292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_360
timestamp 1688980957
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_23
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_46
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_91
timestamp 1688980957
transform 1 0 9476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_97
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_136
timestamp 1688980957
transform 1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_147
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_235
timestamp 1688980957
transform 1 0 22724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_247
timestamp 1688980957
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_259
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_271
timestamp 1688980957
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_287
timestamp 1688980957
transform 1 0 27508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_295
timestamp 1688980957
transform 1 0 28244 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_306
timestamp 1688980957
transform 1 0 29256 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_318
timestamp 1688980957
transform 1 0 30360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_330
timestamp 1688980957
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_378
timestamp 1688980957
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_390
timestamp 1688980957
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_400
timestamp 1688980957
transform 1 0 37904 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_412
timestamp 1688980957
transform 1 0 39008 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_424
timestamp 1688980957
transform 1 0 40112 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_436
timestamp 1688980957
transform 1 0 41216 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_469
timestamp 1688980957
transform 1 0 44252 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_115
timestamp 1688980957
transform 1 0 11684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_125
timestamp 1688980957
transform 1 0 12604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_130
timestamp 1688980957
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_152
timestamp 1688980957
transform 1 0 15088 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_160
timestamp 1688980957
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_166
timestamp 1688980957
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_178
timestamp 1688980957
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_259
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_290
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 1688980957
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_314
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_386
timestamp 1688980957
transform 1 0 36616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_390
timestamp 1688980957
transform 1 0 36984 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_402
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_414
timestamp 1688980957
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_100
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_127
timestamp 1688980957
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_139
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_151
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_196
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_208
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_245
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_272
timestamp 1688980957
transform 1 0 26128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_295
timestamp 1688980957
transform 1 0 28244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_330
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_365
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_371
timestamp 1688980957
transform 1 0 35236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_415
timestamp 1688980957
transform 1 0 39284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_427
timestamp 1688980957
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_439
timestamp 1688980957
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_457
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_465
timestamp 1688980957
transform 1 0 43884 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_66
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_120
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_124
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_128
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_135
timestamp 1688980957
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_185
timestamp 1688980957
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_206
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_218
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_228
timestamp 1688980957
transform 1 0 22080 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_239
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_262
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_268
timestamp 1688980957
transform 1 0 25760 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_278
timestamp 1688980957
transform 1 0 26680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_290
timestamp 1688980957
transform 1 0 27784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_298
timestamp 1688980957
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_306
timestamp 1688980957
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_318
timestamp 1688980957
transform 1 0 30360 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_334
timestamp 1688980957
transform 1 0 31832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_342
timestamp 1688980957
transform 1 0 32568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_371
timestamp 1688980957
transform 1 0 35236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_392
timestamp 1688980957
transform 1 0 37168 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_408
timestamp 1688980957
transform 1 0 38640 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_462
timestamp 1688980957
transform 1 0 43608 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_90
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_98
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_136
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_178
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_186
timestamp 1688980957
transform 1 0 18216 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_208
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_229
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_258
timestamp 1688980957
transform 1 0 24840 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_266
timestamp 1688980957
transform 1 0 25576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_276
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_290
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_340
timestamp 1688980957
transform 1 0 32384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_366
timestamp 1688980957
transform 1 0 34776 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_372
timestamp 1688980957
transform 1 0 35328 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_57
timestamp 1688980957
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_98
timestamp 1688980957
transform 1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_116
timestamp 1688980957
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_127
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_152
timestamp 1688980957
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_160
timestamp 1688980957
transform 1 0 15824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_179
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_205
timestamp 1688980957
transform 1 0 19964 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_212
timestamp 1688980957
transform 1 0 20608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_220
timestamp 1688980957
transform 1 0 21344 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_237
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_262
timestamp 1688980957
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_266
timestamp 1688980957
transform 1 0 25576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_285
timestamp 1688980957
transform 1 0 27324 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_295
timestamp 1688980957
transform 1 0 28244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_332
timestamp 1688980957
transform 1 0 31648 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_400
timestamp 1688980957
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_412
timestamp 1688980957
transform 1 0 39008 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_146
timestamp 1688980957
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_158
timestamp 1688980957
transform 1 0 15640 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_201
timestamp 1688980957
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_213
timestamp 1688980957
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1688980957
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_229
timestamp 1688980957
transform 1 0 22172 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_267
timestamp 1688980957
transform 1 0 25668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1688980957
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_311
timestamp 1688980957
transform 1 0 29716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_319
timestamp 1688980957
transform 1 0 30452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_324
timestamp 1688980957
transform 1 0 30912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_334
timestamp 1688980957
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_340
timestamp 1688980957
transform 1 0 32384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_352
timestamp 1688980957
transform 1 0 33488 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_360
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_372
timestamp 1688980957
transform 1 0 35328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_384
timestamp 1688980957
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_429
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_440
timestamp 1688980957
transform 1 0 41584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_46
timestamp 1688980957
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_58
timestamp 1688980957
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_70
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_103
timestamp 1688980957
transform 1 0 10580 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_167
timestamp 1688980957
transform 1 0 16468 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_179
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_191
timestamp 1688980957
transform 1 0 18676 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_205
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_217
timestamp 1688980957
transform 1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_225
timestamp 1688980957
transform 1 0 21804 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_234
timestamp 1688980957
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_317
timestamp 1688980957
transform 1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_325
timestamp 1688980957
transform 1 0 31004 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_347
timestamp 1688980957
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_359
timestamp 1688980957
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_417
timestamp 1688980957
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1688980957
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_469
timestamp 1688980957
transform 1 0 44252 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_78
timestamp 1688980957
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_90
timestamp 1688980957
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_102
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1688980957
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_127
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_139
timestamp 1688980957
transform 1 0 13892 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_151
timestamp 1688980957
transform 1 0 14996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_158
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1688980957
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_182
timestamp 1688980957
transform 1 0 17848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_191
timestamp 1688980957
transform 1 0 18676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_215
timestamp 1688980957
transform 1 0 20884 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_236
timestamp 1688980957
transform 1 0 22816 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_251
timestamp 1688980957
transform 1 0 24196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_270
timestamp 1688980957
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_297
timestamp 1688980957
transform 1 0 28428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_303
timestamp 1688980957
transform 1 0 28980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_309
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_346
timestamp 1688980957
transform 1 0 32936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_376
timestamp 1688980957
transform 1 0 35696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_384
timestamp 1688980957
transform 1 0 36432 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_421
timestamp 1688980957
transform 1 0 39836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_433
timestamp 1688980957
transform 1 0 40940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_445
timestamp 1688980957
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_461
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_469
timestamp 1688980957
transform 1 0 44252 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_111
timestamp 1688980957
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_125
timestamp 1688980957
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_134
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_169
timestamp 1688980957
transform 1 0 16652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_181
timestamp 1688980957
transform 1 0 17756 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_203
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_215
timestamp 1688980957
transform 1 0 20884 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_239
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_257
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_273
timestamp 1688980957
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_285
timestamp 1688980957
transform 1 0 27324 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_294
timestamp 1688980957
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_306
timestamp 1688980957
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_314
timestamp 1688980957
transform 1 0 29992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_322
timestamp 1688980957
transform 1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_349
timestamp 1688980957
transform 1 0 33212 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_393
timestamp 1688980957
transform 1 0 37260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_410
timestamp 1688980957
transform 1 0 38824 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_90
timestamp 1688980957
transform 1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_98
timestamp 1688980957
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_124
timestamp 1688980957
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_155
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1688980957
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_189
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_201
timestamp 1688980957
transform 1 0 19596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_213
timestamp 1688980957
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_245
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_253
timestamp 1688980957
transform 1 0 24380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_260
timestamp 1688980957
transform 1 0 25024 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_272
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_290
timestamp 1688980957
transform 1 0 27784 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_302
timestamp 1688980957
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_314
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_326
timestamp 1688980957
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_330
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_334
timestamp 1688980957
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_383
timestamp 1688980957
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_397
timestamp 1688980957
transform 1 0 37628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_401
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_411
timestamp 1688980957
transform 1 0 38916 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_423
timestamp 1688980957
transform 1 0 40020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_435
timestamp 1688980957
transform 1 0 41124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_469
timestamp 1688980957
transform 1 0 44252 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_108
timestamp 1688980957
transform 1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_119
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 1688980957
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_161
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_169
timestamp 1688980957
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_175
timestamp 1688980957
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_187
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_207
timestamp 1688980957
transform 1 0 20148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_219
timestamp 1688980957
transform 1 0 21252 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_231
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_243
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_262
timestamp 1688980957
transform 1 0 25208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_268
timestamp 1688980957
transform 1 0 25760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_296
timestamp 1688980957
transform 1 0 28336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_304
timestamp 1688980957
transform 1 0 29072 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_370
timestamp 1688980957
transform 1 0 35144 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_381
timestamp 1688980957
transform 1 0 36156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_393
timestamp 1688980957
transform 1 0 37260 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_399
timestamp 1688980957
transform 1 0 37812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_469
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1688980957
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_73
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_95
timestamp 1688980957
transform 1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_152
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_159
timestamp 1688980957
transform 1 0 15732 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_206
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_235
timestamp 1688980957
transform 1 0 22724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_257
timestamp 1688980957
transform 1 0 24748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_274
timestamp 1688980957
transform 1 0 26312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_289
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_297
timestamp 1688980957
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_320
timestamp 1688980957
transform 1 0 30544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_330
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_367
timestamp 1688980957
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_382
timestamp 1688980957
transform 1 0 36248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_390
timestamp 1688980957
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_421
timestamp 1688980957
transform 1 0 39836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_433
timestamp 1688980957
transform 1 0 40940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_445
timestamp 1688980957
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_461
timestamp 1688980957
transform 1 0 43516 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_469
timestamp 1688980957
transform 1 0 44252 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_108
timestamp 1688980957
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_117
timestamp 1688980957
transform 1 0 11868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_129
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_151
timestamp 1688980957
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_163
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_167
timestamp 1688980957
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_236
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_261
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_273
timestamp 1688980957
transform 1 0 26220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_285
timestamp 1688980957
transform 1 0 27324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_337
timestamp 1688980957
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_418
timestamp 1688980957
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_435
timestamp 1688980957
transform 1 0 41124 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_447
timestamp 1688980957
transform 1 0 42228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_468
timestamp 1688980957
transform 1 0 44160 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_31
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_75
timestamp 1688980957
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_99
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_117
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_122
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_126
timestamp 1688980957
transform 1 0 12696 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_147
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_159
timestamp 1688980957
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_176
timestamp 1688980957
transform 1 0 17296 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_190
timestamp 1688980957
transform 1 0 18584 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_199
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_211
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_387
timestamp 1688980957
transform 1 0 36708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_405
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_460
timestamp 1688980957
transform 1 0 43424 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_469
timestamp 1688980957
transform 1 0 44252 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_45
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_54
timestamp 1688980957
transform 1 0 6072 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_66
timestamp 1688980957
transform 1 0 7176 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_78
timestamp 1688980957
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_151
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_170
timestamp 1688980957
transform 1 0 16744 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_182
timestamp 1688980957
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_261
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_269
timestamp 1688980957
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_291
timestamp 1688980957
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_303
timestamp 1688980957
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_330
timestamp 1688980957
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_342
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_354
timestamp 1688980957
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_362
timestamp 1688980957
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_374
timestamp 1688980957
transform 1 0 35512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_392
timestamp 1688980957
transform 1 0 37168 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_404
timestamp 1688980957
transform 1 0 38272 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_416
timestamp 1688980957
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_464
timestamp 1688980957
transform 1 0 43792 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_23
timestamp 1688980957
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_45
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_104
timestamp 1688980957
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_202
timestamp 1688980957
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_210
timestamp 1688980957
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_229
timestamp 1688980957
transform 1 0 22172 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_240
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_252
timestamp 1688980957
transform 1 0 24288 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_258
timestamp 1688980957
transform 1 0 24840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_289
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_301
timestamp 1688980957
transform 1 0 28796 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_313
timestamp 1688980957
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_325
timestamp 1688980957
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_333
timestamp 1688980957
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_343
timestamp 1688980957
transform 1 0 32660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_364
timestamp 1688980957
transform 1 0 34592 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_368
timestamp 1688980957
transform 1 0 34960 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_389
timestamp 1688980957
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_420
timestamp 1688980957
transform 1 0 39744 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_432
timestamp 1688980957
transform 1 0 40848 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_444
timestamp 1688980957
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_458
timestamp 1688980957
transform 1 0 43240 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_67
timestamp 1688980957
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_128
timestamp 1688980957
transform 1 0 12880 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_150
timestamp 1688980957
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_162
timestamp 1688980957
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_174
timestamp 1688980957
transform 1 0 17112 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_186
timestamp 1688980957
transform 1 0 18216 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_226
timestamp 1688980957
transform 1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_269
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_287
timestamp 1688980957
transform 1 0 27508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_317
timestamp 1688980957
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_340
timestamp 1688980957
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_344
timestamp 1688980957
transform 1 0 32752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_355
timestamp 1688980957
transform 1 0 33764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_362
timestamp 1688980957
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_371
timestamp 1688980957
transform 1 0 35236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_375
timestamp 1688980957
transform 1 0 35604 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_381
timestamp 1688980957
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_402
timestamp 1688980957
transform 1 0 38088 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_418
timestamp 1688980957
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_445
timestamp 1688980957
transform 1 0 42044 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_449
timestamp 1688980957
transform 1 0 42412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_36
timestamp 1688980957
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_63
timestamp 1688980957
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_120
timestamp 1688980957
transform 1 0 12144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_130
timestamp 1688980957
transform 1 0 13064 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1688980957
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_172
timestamp 1688980957
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_183
timestamp 1688980957
transform 1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_213
timestamp 1688980957
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1688980957
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_266
timestamp 1688980957
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_284
timestamp 1688980957
transform 1 0 27232 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_296
timestamp 1688980957
transform 1 0 28336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_304
timestamp 1688980957
transform 1 0 29072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_369
timestamp 1688980957
transform 1 0 35052 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_381
timestamp 1688980957
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_389
timestamp 1688980957
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1688980957
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_417
timestamp 1688980957
transform 1 0 39468 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_426
timestamp 1688980957
transform 1 0 40296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_457
timestamp 1688980957
transform 1 0 43148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_465
timestamp 1688980957
transform 1 0 43884 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1688980957
transform 1 0 11316 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_155
timestamp 1688980957
transform 1 0 15364 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_181
timestamp 1688980957
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1688980957
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_206
timestamp 1688980957
transform 1 0 20056 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_218
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_234
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_242
timestamp 1688980957
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_262
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_274
timestamp 1688980957
transform 1 0 26312 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_323
timestamp 1688980957
transform 1 0 30820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_335
timestamp 1688980957
transform 1 0 31924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_351
timestamp 1688980957
transform 1 0 33396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_359
timestamp 1688980957
transform 1 0 34132 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1688980957
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1688980957
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_416
timestamp 1688980957
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_425
timestamp 1688980957
transform 1 0 40204 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_430
timestamp 1688980957
transform 1 0 40664 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_453
timestamp 1688980957
transform 1 0 42780 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_465
timestamp 1688980957
transform 1 0 43884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_469
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_91
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_122
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_134
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_186
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_211
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_265
timestamp 1688980957
transform 1 0 25484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_294
timestamp 1688980957
transform 1 0 28152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_306
timestamp 1688980957
transform 1 0 29256 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_321
timestamp 1688980957
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_333
timestamp 1688980957
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_366
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_378
timestamp 1688980957
transform 1 0 35880 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_390
timestamp 1688980957
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_420
timestamp 1688980957
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_426
timestamp 1688980957
transform 1 0 40296 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_437
timestamp 1688980957
transform 1 0 41308 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_463
timestamp 1688980957
transform 1 0 43700 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_469
timestamp 1688980957
transform 1 0 44252 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_147
timestamp 1688980957
transform 1 0 14628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_159
timestamp 1688980957
transform 1 0 15732 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_184
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_241
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_292
timestamp 1688980957
transform 1 0 27968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_300
timestamp 1688980957
transform 1 0 28704 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_323
timestamp 1688980957
transform 1 0 30820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_335
timestamp 1688980957
transform 1 0 31924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_341
timestamp 1688980957
transform 1 0 32476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_349
timestamp 1688980957
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_361
timestamp 1688980957
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_369
timestamp 1688980957
transform 1 0 35052 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_410
timestamp 1688980957
transform 1 0 38824 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_441
timestamp 1688980957
transform 1 0 41676 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_23
timestamp 1688980957
transform 1 0 3220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_45
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_77
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_101
timestamp 1688980957
transform 1 0 10396 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_158
timestamp 1688980957
transform 1 0 15640 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_164
timestamp 1688980957
transform 1 0 16192 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_190
timestamp 1688980957
transform 1 0 18584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_202
timestamp 1688980957
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_276
timestamp 1688980957
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_309
timestamp 1688980957
transform 1 0 29532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_320
timestamp 1688980957
transform 1 0 30544 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_332
timestamp 1688980957
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_387
timestamp 1688980957
transform 1 0 36708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_400
timestamp 1688980957
transform 1 0 37904 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_421
timestamp 1688980957
transform 1 0 39836 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_433
timestamp 1688980957
transform 1 0 40940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_444
timestamp 1688980957
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_6
timestamp 1688980957
transform 1 0 1656 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_13
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_25
timestamp 1688980957
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_130
timestamp 1688980957
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_172
timestamp 1688980957
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_214
timestamp 1688980957
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_222
timestamp 1688980957
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_256
timestamp 1688980957
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_275
timestamp 1688980957
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_287
timestamp 1688980957
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_299
timestamp 1688980957
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_355
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_380
timestamp 1688980957
transform 1 0 36064 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_392
timestamp 1688980957
transform 1 0 37168 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_405
timestamp 1688980957
transform 1 0 38364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_429
timestamp 1688980957
transform 1 0 40572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_455
timestamp 1688980957
transform 1 0 42964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_460
timestamp 1688980957
transform 1 0 43424 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_468
timestamp 1688980957
transform 1 0 44160 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_76
timestamp 1688980957
transform 1 0 8096 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_88
timestamp 1688980957
transform 1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_177
timestamp 1688980957
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_213
timestamp 1688980957
transform 1 0 20700 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_232
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_256
timestamp 1688980957
transform 1 0 24656 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_264
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_274
timestamp 1688980957
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_314
timestamp 1688980957
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_333
timestamp 1688980957
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_345
timestamp 1688980957
transform 1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_353
timestamp 1688980957
transform 1 0 33580 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_366
timestamp 1688980957
transform 1 0 34776 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_378
timestamp 1688980957
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_390
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_421
timestamp 1688980957
transform 1 0 39836 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_433
timestamp 1688980957
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_445
timestamp 1688980957
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_463
timestamp 1688980957
transform 1 0 43700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_469
timestamp 1688980957
transform 1 0 44252 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_70
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_82
timestamp 1688980957
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_119
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_150
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_206
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_210
timestamp 1688980957
transform 1 0 20424 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_231
timestamp 1688980957
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_243
timestamp 1688980957
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_272
timestamp 1688980957
transform 1 0 26128 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_284
timestamp 1688980957
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_288
timestamp 1688980957
transform 1 0 27600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_318
timestamp 1688980957
transform 1 0 30360 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_327
timestamp 1688980957
transform 1 0 31188 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_341
timestamp 1688980957
transform 1 0 32476 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_349
timestamp 1688980957
transform 1 0 33212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_360
timestamp 1688980957
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_418
timestamp 1688980957
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_428
timestamp 1688980957
transform 1 0 40480 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_440
timestamp 1688980957
transform 1 0 41584 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_448
timestamp 1688980957
transform 1 0 42320 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_455
timestamp 1688980957
transform 1 0 42964 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_467
timestamp 1688980957
transform 1 0 44068 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_101
timestamp 1688980957
transform 1 0 10396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_122
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_133
timestamp 1688980957
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_141
timestamp 1688980957
transform 1 0 14076 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_151
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1688980957
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_212
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_248
timestamp 1688980957
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_260
timestamp 1688980957
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_272
timestamp 1688980957
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_324
timestamp 1688980957
transform 1 0 30912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_333
timestamp 1688980957
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_365
timestamp 1688980957
transform 1 0 34684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_390
timestamp 1688980957
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_420
timestamp 1688980957
transform 1 0 39744 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_432
timestamp 1688980957
transform 1 0 40848 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_444
timestamp 1688980957
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_454
timestamp 1688980957
transform 1 0 42872 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_466
timestamp 1688980957
transform 1 0 43976 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_105
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_117
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_129
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1688980957
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_150
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_162
timestamp 1688980957
transform 1 0 16008 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_168
timestamp 1688980957
transform 1 0 16560 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_178
timestamp 1688980957
transform 1 0 17480 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_186
timestamp 1688980957
transform 1 0 18216 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_190
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_222
timestamp 1688980957
transform 1 0 21528 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_230
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_293
timestamp 1688980957
transform 1 0 28060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_319
timestamp 1688980957
transform 1 0 30452 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_325
timestamp 1688980957
transform 1 0 31004 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_347
timestamp 1688980957
transform 1 0 33028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_373
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_387
timestamp 1688980957
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_399
timestamp 1688980957
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_429
timestamp 1688980957
transform 1 0 40572 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_435
timestamp 1688980957
transform 1 0 41124 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_439
timestamp 1688980957
transform 1 0 41492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_463
timestamp 1688980957
transform 1 0 43700 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_77
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_89
timestamp 1688980957
transform 1 0 9292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_101
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_126
timestamp 1688980957
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_156
timestamp 1688980957
transform 1 0 15456 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_163
timestamp 1688980957
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_235
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_242
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_272
timestamp 1688980957
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_287
timestamp 1688980957
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_303
timestamp 1688980957
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_353
timestamp 1688980957
transform 1 0 33580 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_363
timestamp 1688980957
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_375
timestamp 1688980957
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_387
timestamp 1688980957
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_414
timestamp 1688980957
transform 1 0 39192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_418
timestamp 1688980957
transform 1 0 39560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_426
timestamp 1688980957
transform 1 0 40296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_433
timestamp 1688980957
transform 1 0 40940 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_446
timestamp 1688980957
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_462
timestamp 1688980957
transform 1 0 43608 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_93
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_115
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_176
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_188
timestamp 1688980957
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_215
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_236
timestamp 1688980957
transform 1 0 22816 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_271
timestamp 1688980957
transform 1 0 26036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 1688980957
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_317
timestamp 1688980957
transform 1 0 30268 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_326
timestamp 1688980957
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_338
timestamp 1688980957
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_350
timestamp 1688980957
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_362
timestamp 1688980957
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_375
timestamp 1688980957
transform 1 0 35604 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_387
timestamp 1688980957
transform 1 0 36708 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_399
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_411
timestamp 1688980957
transform 1 0 38916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_443
timestamp 1688980957
transform 1 0 41860 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_447
timestamp 1688980957
transform 1 0 42228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_468
timestamp 1688980957
transform 1 0 44160 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_89
timestamp 1688980957
transform 1 0 9292 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_122
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_189
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_204
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_216
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_228
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_236
timestamp 1688980957
transform 1 0 22816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_276
timestamp 1688980957
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_296
timestamp 1688980957
transform 1 0 28336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_304
timestamp 1688980957
transform 1 0 29072 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_323
timestamp 1688980957
transform 1 0 30820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_347
timestamp 1688980957
transform 1 0 33028 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_353
timestamp 1688980957
transform 1 0 33580 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_362
timestamp 1688980957
transform 1 0 34408 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_413
timestamp 1688980957
transform 1 0 39100 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_427
timestamp 1688980957
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_439
timestamp 1688980957
transform 1 0 41492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 1688980957
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_460
timestamp 1688980957
transform 1 0 43424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_468
timestamp 1688980957
transform 1 0 44160 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_106
timestamp 1688980957
transform 1 0 10856 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_116
timestamp 1688980957
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_128
timestamp 1688980957
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_144
timestamp 1688980957
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_161
timestamp 1688980957
transform 1 0 15916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_169
timestamp 1688980957
transform 1 0 16652 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_182
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_186
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_227
timestamp 1688980957
transform 1 0 21988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_231
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_257
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_278
timestamp 1688980957
transform 1 0 26680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_282
timestamp 1688980957
transform 1 0 27048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_340
timestamp 1688980957
transform 1 0 32384 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_346
timestamp 1688980957
transform 1 0 32936 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_361
timestamp 1688980957
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_369
timestamp 1688980957
transform 1 0 35052 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_378
timestamp 1688980957
transform 1 0 35880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_410
timestamp 1688980957
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_418
timestamp 1688980957
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 1688980957
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_445
timestamp 1688980957
transform 1 0 42044 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_451
timestamp 1688980957
transform 1 0 42596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_459
timestamp 1688980957
transform 1 0 43332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_467
timestamp 1688980957
transform 1 0 44068 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_131
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_163
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_188
timestamp 1688980957
transform 1 0 18400 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_200
timestamp 1688980957
transform 1 0 19504 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_233
timestamp 1688980957
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_242
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_254
timestamp 1688980957
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 1688980957
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_332
timestamp 1688980957
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_353
timestamp 1688980957
transform 1 0 33580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_370
timestamp 1688980957
transform 1 0 35144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_442
timestamp 1688980957
transform 1 0 41768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_463
timestamp 1688980957
transform 1 0 43700 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_469
timestamp 1688980957
transform 1 0 44252 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_113
timestamp 1688980957
transform 1 0 11500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_134
timestamp 1688980957
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_144
timestamp 1688980957
transform 1 0 14352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_148
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_172
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_225
timestamp 1688980957
transform 1 0 21804 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_237
timestamp 1688980957
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_261
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_273
timestamp 1688980957
transform 1 0 26220 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_285
timestamp 1688980957
transform 1 0 27324 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_297
timestamp 1688980957
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_305
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_313
timestamp 1688980957
transform 1 0 29900 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_328
timestamp 1688980957
transform 1 0 31280 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_340
timestamp 1688980957
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_373
timestamp 1688980957
transform 1 0 35420 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_385
timestamp 1688980957
transform 1 0 36524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_393
timestamp 1688980957
transform 1 0 37260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_397
timestamp 1688980957
transform 1 0 37628 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_409
timestamp 1688980957
transform 1 0 38732 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 1688980957
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_449
timestamp 1688980957
transform 1 0 42412 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_469
timestamp 1688980957
transform 1 0 44252 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_101
timestamp 1688980957
transform 1 0 10396 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_122
timestamp 1688980957
transform 1 0 12328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_134
timestamp 1688980957
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_189
timestamp 1688980957
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_197
timestamp 1688980957
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_209
timestamp 1688980957
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_253
timestamp 1688980957
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_265
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_274
timestamp 1688980957
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_291
timestamp 1688980957
transform 1 0 27876 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_303
timestamp 1688980957
transform 1 0 28980 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_315
timestamp 1688980957
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_327
timestamp 1688980957
transform 1 0 31188 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_357
timestamp 1688980957
transform 1 0 33948 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_369
timestamp 1688980957
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_390
timestamp 1688980957
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_411
timestamp 1688980957
transform 1 0 38916 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_421
timestamp 1688980957
transform 1 0 39836 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_433
timestamp 1688980957
transform 1 0 40940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_445
timestamp 1688980957
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_49
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_76
timestamp 1688980957
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_129
timestamp 1688980957
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1688980957
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_144
timestamp 1688980957
transform 1 0 14352 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_156
timestamp 1688980957
transform 1 0 15456 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_168
timestamp 1688980957
transform 1 0 16560 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_183
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_200
timestamp 1688980957
transform 1 0 19504 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_204
timestamp 1688980957
transform 1 0 19872 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_211
timestamp 1688980957
transform 1 0 20516 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 1688980957
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_261
timestamp 1688980957
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_287
timestamp 1688980957
transform 1 0 27508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_295
timestamp 1688980957
transform 1 0 28244 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_306
timestamp 1688980957
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_312
timestamp 1688980957
transform 1 0 29808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_324
timestamp 1688980957
transform 1 0 30912 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_330
timestamp 1688980957
transform 1 0 31464 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_334
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_343
timestamp 1688980957
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_355
timestamp 1688980957
transform 1 0 33764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_403
timestamp 1688980957
transform 1 0 38180 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_414
timestamp 1688980957
transform 1 0 39192 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_435
timestamp 1688980957
transform 1 0 41124 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_447
timestamp 1688980957
transform 1 0 42228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_60
timestamp 1688980957
transform 1 0 6624 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_134
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_140
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_179
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_191
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_197
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_218
timestamp 1688980957
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_233
timestamp 1688980957
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_265
timestamp 1688980957
transform 1 0 25484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_316
timestamp 1688980957
transform 1 0 30176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_328
timestamp 1688980957
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_347
timestamp 1688980957
transform 1 0 33028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_351
timestamp 1688980957
transform 1 0 33396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_401
timestamp 1688980957
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_430
timestamp 1688980957
transform 1 0 40664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_434
timestamp 1688980957
transform 1 0 41032 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_443
timestamp 1688980957
transform 1 0 41860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_469
timestamp 1688980957
transform 1 0 44252 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_47
timestamp 1688980957
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_59
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_71
timestamp 1688980957
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_89
timestamp 1688980957
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_110
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_118
timestamp 1688980957
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_150
timestamp 1688980957
transform 1 0 14904 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_161
timestamp 1688980957
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_184
timestamp 1688980957
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_222
timestamp 1688980957
transform 1 0 21528 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_234
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_299
timestamp 1688980957
transform 1 0 28612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_323
timestamp 1688980957
transform 1 0 30820 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_399
timestamp 1688980957
transform 1 0 37812 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_408
timestamp 1688980957
transform 1 0 38640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_461
timestamp 1688980957
transform 1 0 43516 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_101
timestamp 1688980957
transform 1 0 10396 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_109
timestamp 1688980957
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_189
timestamp 1688980957
transform 1 0 18492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_201
timestamp 1688980957
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_215
timestamp 1688980957
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_230
timestamp 1688980957
transform 1 0 22264 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_242
timestamp 1688980957
transform 1 0 23368 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_258
timestamp 1688980957
transform 1 0 24840 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_270
timestamp 1688980957
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_312
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_324
timestamp 1688980957
transform 1 0 30912 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_340
timestamp 1688980957
transform 1 0 32384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_352
timestamp 1688980957
transform 1 0 33488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_360
timestamp 1688980957
transform 1 0 34224 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_376
timestamp 1688980957
transform 1 0 35696 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_407
timestamp 1688980957
transform 1 0 38548 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_419
timestamp 1688980957
transform 1 0 39652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_423
timestamp 1688980957
transform 1 0 40020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_6
timestamp 1688980957
transform 1 0 1656 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_18
timestamp 1688980957
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1688980957
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_103
timestamp 1688980957
transform 1 0 10580 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_124
timestamp 1688980957
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_136
timestamp 1688980957
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_154
timestamp 1688980957
transform 1 0 15272 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_256
timestamp 1688980957
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_280
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_292
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_303
timestamp 1688980957
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_341
timestamp 1688980957
transform 1 0 32476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_359
timestamp 1688980957
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_387
timestamp 1688980957
transform 1 0 36708 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_416
timestamp 1688980957
transform 1 0 39376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_429
timestamp 1688980957
transform 1 0 40572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_440
timestamp 1688980957
transform 1 0 41584 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_448
timestamp 1688980957
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_469
timestamp 1688980957
transform 1 0 44252 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_45
timestamp 1688980957
transform 1 0 5244 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_75
timestamp 1688980957
transform 1 0 8004 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_96
timestamp 1688980957
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_108
timestamp 1688980957
transform 1 0 11040 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_122
timestamp 1688980957
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_131
timestamp 1688980957
transform 1 0 13156 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_197
timestamp 1688980957
transform 1 0 19228 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_209
timestamp 1688980957
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_213
timestamp 1688980957
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_245
timestamp 1688980957
transform 1 0 23644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1688980957
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_292
timestamp 1688980957
transform 1 0 27968 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_327
timestamp 1688980957
transform 1 0 31188 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_340
timestamp 1688980957
transform 1 0 32384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_348
timestamp 1688980957
transform 1 0 33120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_433
timestamp 1688980957
transform 1 0 40940 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_443
timestamp 1688980957
transform 1 0 41860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 1688980957
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_449
timestamp 1688980957
transform 1 0 42412 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_57
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_72
timestamp 1688980957
transform 1 0 7728 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_105
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_114
timestamp 1688980957
transform 1 0 11592 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_129
timestamp 1688980957
transform 1 0 12972 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_136
timestamp 1688980957
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_149
timestamp 1688980957
transform 1 0 14812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_173
timestamp 1688980957
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_181
timestamp 1688980957
transform 1 0 17756 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_191
timestamp 1688980957
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_212
timestamp 1688980957
transform 1 0 20608 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_216
timestamp 1688980957
transform 1 0 20976 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_228
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_283
timestamp 1688980957
transform 1 0 27140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_294
timestamp 1688980957
transform 1 0 28152 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_302
timestamp 1688980957
transform 1 0 28888 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_306
timestamp 1688980957
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_350
timestamp 1688980957
transform 1 0 33304 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_359
timestamp 1688980957
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_373
timestamp 1688980957
transform 1 0 35420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_395
timestamp 1688980957
transform 1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_407
timestamp 1688980957
transform 1 0 38548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_411
timestamp 1688980957
transform 1 0 38916 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_36
timestamp 1688980957
transform 1 0 4416 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_52
timestamp 1688980957
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_85
timestamp 1688980957
transform 1 0 8924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1688980957
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_175
timestamp 1688980957
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_187
timestamp 1688980957
transform 1 0 18308 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_199
timestamp 1688980957
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_258
timestamp 1688980957
transform 1 0 24840 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_270
timestamp 1688980957
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_278
timestamp 1688980957
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_294
timestamp 1688980957
transform 1 0 28152 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_306
timestamp 1688980957
transform 1 0 29256 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_314
timestamp 1688980957
transform 1 0 29992 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_322
timestamp 1688980957
transform 1 0 30728 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_331
timestamp 1688980957
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_345
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_354
timestamp 1688980957
transform 1 0 33672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_362
timestamp 1688980957
transform 1 0 34408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_369
timestamp 1688980957
transform 1 0 35052 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_377
timestamp 1688980957
transform 1 0 35788 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_387
timestamp 1688980957
transform 1 0 36708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_409
timestamp 1688980957
transform 1 0 38732 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_431
timestamp 1688980957
transform 1 0 40756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_443
timestamp 1688980957
transform 1 0 41860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_449
timestamp 1688980957
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_453
timestamp 1688980957
transform 1 0 42780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_462
timestamp 1688980957
transform 1 0 43608 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_60
timestamp 1688980957
transform 1 0 6624 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_68
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_78
timestamp 1688980957
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_93
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_105
timestamp 1688980957
transform 1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_131
timestamp 1688980957
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_188
timestamp 1688980957
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_262
timestamp 1688980957
transform 1 0 25208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_274
timestamp 1688980957
transform 1 0 26312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_282
timestamp 1688980957
transform 1 0 27048 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_351
timestamp 1688980957
transform 1 0 33396 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_360
timestamp 1688980957
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_369
timestamp 1688980957
transform 1 0 35052 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_376
timestamp 1688980957
transform 1 0 35696 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_388
timestamp 1688980957
transform 1 0 36800 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_400
timestamp 1688980957
transform 1 0 37904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_404
timestamp 1688980957
transform 1 0 38272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_429
timestamp 1688980957
transform 1 0 40572 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_461
timestamp 1688980957
transform 1 0 43516 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_469
timestamp 1688980957
transform 1 0 44252 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_45
timestamp 1688980957
transform 1 0 5244 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_70
timestamp 1688980957
transform 1 0 7544 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_101
timestamp 1688980957
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_106
timestamp 1688980957
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_120
timestamp 1688980957
transform 1 0 12144 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_141
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_155
timestamp 1688980957
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_192
timestamp 1688980957
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_219
timestamp 1688980957
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_271
timestamp 1688980957
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_289
timestamp 1688980957
transform 1 0 27692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_301
timestamp 1688980957
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_316
timestamp 1688980957
transform 1 0 30176 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_328
timestamp 1688980957
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_346
timestamp 1688980957
transform 1 0 32936 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_355
timestamp 1688980957
transform 1 0 33764 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_366
timestamp 1688980957
transform 1 0 34776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_445
timestamp 1688980957
transform 1 0 42044 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_457
timestamp 1688980957
transform 1 0 43148 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_469
timestamp 1688980957
transform 1 0 44252 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_55
timestamp 1688980957
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_59
timestamp 1688980957
transform 1 0 6532 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_78
timestamp 1688980957
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_107
timestamp 1688980957
transform 1 0 10948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_113
timestamp 1688980957
transform 1 0 11500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_157
timestamp 1688980957
transform 1 0 15548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_169
timestamp 1688980957
transform 1 0 16652 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_181
timestamp 1688980957
transform 1 0 17756 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_185
timestamp 1688980957
transform 1 0 18124 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_222
timestamp 1688980957
transform 1 0 21528 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_261
timestamp 1688980957
transform 1 0 25116 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_372
timestamp 1688980957
transform 1 0 35328 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_394
timestamp 1688980957
transform 1 0 37352 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_398
timestamp 1688980957
transform 1 0 37720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_418
timestamp 1688980957
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_444
timestamp 1688980957
transform 1 0 41952 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_468
timestamp 1688980957
transform 1 0 44160 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_77
timestamp 1688980957
transform 1 0 8188 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_91
timestamp 1688980957
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_103
timestamp 1688980957
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_120
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_132
timestamp 1688980957
transform 1 0 13248 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_196
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_208
timestamp 1688980957
transform 1 0 20240 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_254
timestamp 1688980957
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_262
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_324
timestamp 1688980957
transform 1 0 30912 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_343
timestamp 1688980957
transform 1 0 32660 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_352
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_375
timestamp 1688980957
transform 1 0 35604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_387
timestamp 1688980957
transform 1 0 36708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_446
timestamp 1688980957
transform 1 0 42136 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_458
timestamp 1688980957
transform 1 0 43240 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_67
timestamp 1688980957
transform 1 0 7268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_81
timestamp 1688980957
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_88
timestamp 1688980957
transform 1 0 9200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_113
timestamp 1688980957
transform 1 0 11500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_122
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_134
timestamp 1688980957
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_157
timestamp 1688980957
transform 1 0 15548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_169
timestamp 1688980957
transform 1 0 16652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_179
timestamp 1688980957
transform 1 0 17572 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_191
timestamp 1688980957
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_220
timestamp 1688980957
transform 1 0 21344 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_232
timestamp 1688980957
transform 1 0 22448 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_244
timestamp 1688980957
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_264
timestamp 1688980957
transform 1 0 25392 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_276
timestamp 1688980957
transform 1 0 26496 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_288
timestamp 1688980957
transform 1 0 27600 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_300
timestamp 1688980957
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_339
timestamp 1688980957
transform 1 0 32292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_351
timestamp 1688980957
transform 1 0 33396 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_383
timestamp 1688980957
transform 1 0 36340 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_411
timestamp 1688980957
transform 1 0 38916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_436
timestamp 1688980957
transform 1 0 41216 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_448
timestamp 1688980957
transform 1 0 42320 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_68
timestamp 1688980957
transform 1 0 7360 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_72
timestamp 1688980957
transform 1 0 7728 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_76
timestamp 1688980957
transform 1 0 8096 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_108
timestamp 1688980957
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_202
timestamp 1688980957
transform 1 0 19688 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_214
timestamp 1688980957
transform 1 0 20792 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1688980957
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_231
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_255
timestamp 1688980957
transform 1 0 24564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_278
timestamp 1688980957
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_289
timestamp 1688980957
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_323
timestamp 1688980957
transform 1 0 30820 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_327
timestamp 1688980957
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_360
timestamp 1688980957
transform 1 0 34224 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_376
timestamp 1688980957
transform 1 0 35696 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_388
timestamp 1688980957
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_441
timestamp 1688980957
transform 1 0 41676 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_449
timestamp 1688980957
transform 1 0 42412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_457
timestamp 1688980957
transform 1 0 43148 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_462
timestamp 1688980957
transform 1 0 43608 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_37
timestamp 1688980957
transform 1 0 4508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_50
timestamp 1688980957
transform 1 0 5704 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_62
timestamp 1688980957
transform 1 0 6808 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_129
timestamp 1688980957
transform 1 0 12972 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_149
timestamp 1688980957
transform 1 0 14812 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_157
timestamp 1688980957
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_178
timestamp 1688980957
transform 1 0 17480 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_184
timestamp 1688980957
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_206
timestamp 1688980957
transform 1 0 20056 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_214
timestamp 1688980957
transform 1 0 20792 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_220
timestamp 1688980957
transform 1 0 21344 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_224
timestamp 1688980957
transform 1 0 21712 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_303
timestamp 1688980957
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_332
timestamp 1688980957
transform 1 0 31648 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_344
timestamp 1688980957
transform 1 0 32752 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_352
timestamp 1688980957
transform 1 0 33488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_362
timestamp 1688980957
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_372
timestamp 1688980957
transform 1 0 35328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_384
timestamp 1688980957
transform 1 0 36432 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_402
timestamp 1688980957
transform 1 0 38088 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_414
timestamp 1688980957
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_427
timestamp 1688980957
transform 1 0 40388 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_439
timestamp 1688980957
transform 1 0 41492 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_451
timestamp 1688980957
transform 1 0 42596 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_465
timestamp 1688980957
transform 1 0 43884 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_469
timestamp 1688980957
transform 1 0 44252 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_62
timestamp 1688980957
transform 1 0 6808 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_74
timestamp 1688980957
transform 1 0 7912 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_86
timestamp 1688980957
transform 1 0 9016 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_92
timestamp 1688980957
transform 1 0 9568 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_104
timestamp 1688980957
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_158
timestamp 1688980957
transform 1 0 15640 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_163
timestamp 1688980957
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_186
timestamp 1688980957
transform 1 0 18216 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_203
timestamp 1688980957
transform 1 0 19780 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_222
timestamp 1688980957
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_250
timestamp 1688980957
transform 1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_254
timestamp 1688980957
transform 1 0 24472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_301
timestamp 1688980957
transform 1 0 28796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_334
timestamp 1688980957
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_345
timestamp 1688980957
transform 1 0 32844 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_366
timestamp 1688980957
transform 1 0 34776 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_375
timestamp 1688980957
transform 1 0 35604 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_388
timestamp 1688980957
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_413
timestamp 1688980957
transform 1 0 39100 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_435
timestamp 1688980957
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1688980957
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_469
timestamp 1688980957
transform 1 0 44252 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_47
timestamp 1688980957
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_51
timestamp 1688980957
transform 1 0 5796 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_57
timestamp 1688980957
transform 1 0 6348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_69
timestamp 1688980957
transform 1 0 7452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_89
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_95
timestamp 1688980957
transform 1 0 9844 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_104
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_144
timestamp 1688980957
transform 1 0 14352 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_151
timestamp 1688980957
transform 1 0 14996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_157
timestamp 1688980957
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_184
timestamp 1688980957
transform 1 0 18032 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_205
timestamp 1688980957
transform 1 0 19964 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_211
timestamp 1688980957
transform 1 0 20516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_223
timestamp 1688980957
transform 1 0 21620 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_240
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_250
timestamp 1688980957
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_269
timestamp 1688980957
transform 1 0 25852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_298
timestamp 1688980957
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_313
timestamp 1688980957
transform 1 0 29900 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_328
timestamp 1688980957
transform 1 0 31280 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_349
timestamp 1688980957
transform 1 0 33212 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_372
timestamp 1688980957
transform 1 0 35328 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_384
timestamp 1688980957
transform 1 0 36432 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_388
timestamp 1688980957
transform 1 0 36800 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_397
timestamp 1688980957
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_425
timestamp 1688980957
transform 1 0 40204 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_434
timestamp 1688980957
transform 1 0 41032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_456
timestamp 1688980957
transform 1 0 43056 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_464
timestamp 1688980957
transform 1 0 43792 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_54
timestamp 1688980957
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_63
timestamp 1688980957
transform 1 0 6900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_67
timestamp 1688980957
transform 1 0 7268 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_75
timestamp 1688980957
transform 1 0 8004 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_106
timestamp 1688980957
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_116
timestamp 1688980957
transform 1 0 11776 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_122
timestamp 1688980957
transform 1 0 12328 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_132
timestamp 1688980957
transform 1 0 13248 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_144
timestamp 1688980957
transform 1 0 14352 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_165
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_173
timestamp 1688980957
transform 1 0 17020 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_202
timestamp 1688980957
transform 1 0 19688 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_214
timestamp 1688980957
transform 1 0 20792 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_222
timestamp 1688980957
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_233
timestamp 1688980957
transform 1 0 22540 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_250
timestamp 1688980957
transform 1 0 24104 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_271
timestamp 1688980957
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_288
timestamp 1688980957
transform 1 0 27600 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_292
timestamp 1688980957
transform 1 0 27968 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_302
timestamp 1688980957
transform 1 0 28888 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_314
timestamp 1688980957
transform 1 0 29992 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_325
timestamp 1688980957
transform 1 0 31004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_333
timestamp 1688980957
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_376
timestamp 1688980957
transform 1 0 35696 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_389
timestamp 1688980957
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_433
timestamp 1688980957
transform 1 0 40940 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_441
timestamp 1688980957
transform 1 0 41676 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_113
timestamp 1688980957
transform 1 0 11500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_125
timestamp 1688980957
transform 1 0 12604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_137
timestamp 1688980957
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_147
timestamp 1688980957
transform 1 0 14628 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_167
timestamp 1688980957
transform 1 0 16468 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_217
timestamp 1688980957
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_229
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_244
timestamp 1688980957
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_262
timestamp 1688980957
transform 1 0 25208 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_270
timestamp 1688980957
transform 1 0 25944 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_276
timestamp 1688980957
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_288
timestamp 1688980957
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_300
timestamp 1688980957
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_336
timestamp 1688980957
transform 1 0 32016 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_348
timestamp 1688980957
transform 1 0 33120 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_360
timestamp 1688980957
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_376
timestamp 1688980957
transform 1 0 35696 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_398
timestamp 1688980957
transform 1 0 37720 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_406
timestamp 1688980957
transform 1 0 38456 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_436
timestamp 1688980957
transform 1 0 41216 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_448
timestamp 1688980957
transform 1 0 42320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_462
timestamp 1688980957
transform 1 0 43608 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_20
timestamp 1688980957
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_32
timestamp 1688980957
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_44
timestamp 1688980957
transform 1 0 5152 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_52
timestamp 1688980957
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_72
timestamp 1688980957
transform 1 0 7728 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_84
timestamp 1688980957
transform 1 0 8832 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_96
timestamp 1688980957
transform 1 0 9936 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_108
timestamp 1688980957
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_122
timestamp 1688980957
transform 1 0 12328 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_127
timestamp 1688980957
transform 1 0 12788 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_139
timestamp 1688980957
transform 1 0 13892 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_150
timestamp 1688980957
transform 1 0 14904 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_160
timestamp 1688980957
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_173
timestamp 1688980957
transform 1 0 17020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_178
timestamp 1688980957
transform 1 0 17480 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_186
timestamp 1688980957
transform 1 0 18216 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_197
timestamp 1688980957
transform 1 0 19228 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_211
timestamp 1688980957
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_245
timestamp 1688980957
transform 1 0 23644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_257
timestamp 1688980957
transform 1 0 24748 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_298
timestamp 1688980957
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_319
timestamp 1688980957
transform 1 0 30452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_325
timestamp 1688980957
transform 1 0 31004 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_344
timestamp 1688980957
transform 1 0 32752 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_348
timestamp 1688980957
transform 1 0 33120 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_354
timestamp 1688980957
transform 1 0 33672 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_362
timestamp 1688980957
transform 1 0 34408 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_384
timestamp 1688980957
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_413
timestamp 1688980957
transform 1 0 39100 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_444
timestamp 1688980957
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_469
timestamp 1688980957
transform 1 0 44252 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_49
timestamp 1688980957
transform 1 0 5612 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_55
timestamp 1688980957
transform 1 0 6164 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_103
timestamp 1688980957
transform 1 0 10580 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_115
timestamp 1688980957
transform 1 0 11684 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_136
timestamp 1688980957
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_149
timestamp 1688980957
transform 1 0 14812 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_178
timestamp 1688980957
transform 1 0 17480 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_190
timestamp 1688980957
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_217
timestamp 1688980957
transform 1 0 21068 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_250
timestamp 1688980957
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_261
timestamp 1688980957
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_268
timestamp 1688980957
transform 1 0 25760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_272
timestamp 1688980957
transform 1 0 26128 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_299
timestamp 1688980957
transform 1 0 28612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_361
timestamp 1688980957
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_411
timestamp 1688980957
transform 1 0 38916 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_425
timestamp 1688980957
transform 1 0 40204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_437
timestamp 1688980957
transform 1 0 41308 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_458
timestamp 1688980957
transform 1 0 43240 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_13
timestamp 1688980957
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_25
timestamp 1688980957
transform 1 0 3404 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_33
timestamp 1688980957
transform 1 0 4140 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_83
timestamp 1688980957
transform 1 0 8740 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_91
timestamp 1688980957
transform 1 0 9476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_141
timestamp 1688980957
transform 1 0 14076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_153
timestamp 1688980957
transform 1 0 15180 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_157
timestamp 1688980957
transform 1 0 15548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_209
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_221
timestamp 1688980957
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_238
timestamp 1688980957
transform 1 0 23000 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_267
timestamp 1688980957
transform 1 0 25668 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_275
timestamp 1688980957
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_284
timestamp 1688980957
transform 1 0 27232 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_298
timestamp 1688980957
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_310
timestamp 1688980957
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_318
timestamp 1688980957
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_330
timestamp 1688980957
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_379
timestamp 1688980957
transform 1 0 35972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_397
timestamp 1688980957
transform 1 0 37628 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_404
timestamp 1688980957
transform 1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_415
timestamp 1688980957
transform 1 0 39284 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_423
timestamp 1688980957
transform 1 0 40020 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_432
timestamp 1688980957
transform 1 0 40848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_469
timestamp 1688980957
transform 1 0 44252 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_6
timestamp 1688980957
transform 1 0 1656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_18
timestamp 1688980957
transform 1 0 2760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_26
timestamp 1688980957
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_68
timestamp 1688980957
transform 1 0 7360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_80
timestamp 1688980957
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_90
timestamp 1688980957
transform 1 0 9384 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_102
timestamp 1688980957
transform 1 0 10488 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_113
timestamp 1688980957
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_154
timestamp 1688980957
transform 1 0 15272 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_164
timestamp 1688980957
transform 1 0 16192 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_170
timestamp 1688980957
transform 1 0 16744 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_217
timestamp 1688980957
transform 1 0 21068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_229
timestamp 1688980957
transform 1 0 22172 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_248
timestamp 1688980957
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_270
timestamp 1688980957
transform 1 0 25944 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_291
timestamp 1688980957
transform 1 0 27876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_303
timestamp 1688980957
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_352
timestamp 1688980957
transform 1 0 33488 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_397
timestamp 1688980957
transform 1 0 37628 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_404
timestamp 1688980957
transform 1 0 38272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_416
timestamp 1688980957
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_441
timestamp 1688980957
transform 1 0 41676 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_87
timestamp 1688980957
transform 1 0 9108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_110
timestamp 1688980957
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_135
timestamp 1688980957
transform 1 0 13524 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_163
timestamp 1688980957
transform 1 0 16100 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_221
timestamp 1688980957
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_234
timestamp 1688980957
transform 1 0 22632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_246
timestamp 1688980957
transform 1 0 23736 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_252
timestamp 1688980957
transform 1 0 24288 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_265
timestamp 1688980957
transform 1 0 25484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_277
timestamp 1688980957
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_308
timestamp 1688980957
transform 1 0 29440 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_328
timestamp 1688980957
transform 1 0 31280 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_345
timestamp 1688980957
transform 1 0 32844 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_353
timestamp 1688980957
transform 1 0 33580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_365
timestamp 1688980957
transform 1 0 34684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_411
timestamp 1688980957
transform 1 0 38916 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_419
timestamp 1688980957
transform 1 0 39652 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_426
timestamp 1688980957
transform 1 0 40296 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_438
timestamp 1688980957
transform 1 0 41400 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_446
timestamp 1688980957
transform 1 0 42136 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_449
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_459
timestamp 1688980957
transform 1 0 43332 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_469
timestamp 1688980957
transform 1 0 44252 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_57
timestamp 1688980957
transform 1 0 6348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_78
timestamp 1688980957
transform 1 0 8280 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_104
timestamp 1688980957
transform 1 0 10672 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_114
timestamp 1688980957
transform 1 0 11592 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_126
timestamp 1688980957
transform 1 0 12696 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_137
timestamp 1688980957
transform 1 0 13708 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_157
timestamp 1688980957
transform 1 0 15548 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_261
timestamp 1688980957
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_284
timestamp 1688980957
transform 1 0 27232 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_338
timestamp 1688980957
transform 1 0 32200 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_342
timestamp 1688980957
transform 1 0 32568 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_356
timestamp 1688980957
transform 1 0 33856 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_388
timestamp 1688980957
transform 1 0 36800 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_396
timestamp 1688980957
transform 1 0 37536 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_409
timestamp 1688980957
transform 1 0 38732 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_417
timestamp 1688980957
transform 1 0 39468 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_441
timestamp 1688980957
transform 1 0 41676 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_461
timestamp 1688980957
transform 1 0 43516 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_469
timestamp 1688980957
transform 1 0 44252 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_68
timestamp 1688980957
transform 1 0 7360 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_94
timestamp 1688980957
transform 1 0 9752 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_100
timestamp 1688980957
transform 1 0 10304 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_186
timestamp 1688980957
transform 1 0 18216 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_198
timestamp 1688980957
transform 1 0 19320 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_213
timestamp 1688980957
transform 1 0 20700 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_221
timestamp 1688980957
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_235
timestamp 1688980957
transform 1 0 22724 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_290
timestamp 1688980957
transform 1 0 27784 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_320
timestamp 1688980957
transform 1 0 30544 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_332
timestamp 1688980957
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_353
timestamp 1688980957
transform 1 0 33580 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_362
timestamp 1688980957
transform 1 0 34408 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_374
timestamp 1688980957
transform 1 0 35512 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_413
timestamp 1688980957
transform 1 0 39100 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_421
timestamp 1688980957
transform 1 0 39836 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_432
timestamp 1688980957
transform 1 0 40848 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_444
timestamp 1688980957
transform 1 0 41952 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_71
timestamp 1688980957
transform 1 0 7636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_91
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_112
timestamp 1688980957
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_163
timestamp 1688980957
transform 1 0 16100 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_187
timestamp 1688980957
transform 1 0 18308 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_217
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_225
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_234
timestamp 1688980957
transform 1 0 22632 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_246
timestamp 1688980957
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_273
timestamp 1688980957
transform 1 0 26220 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_295
timestamp 1688980957
transform 1 0 28244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_304
timestamp 1688980957
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_372
timestamp 1688980957
transform 1 0 35328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_384
timestamp 1688980957
transform 1 0 36432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_396
timestamp 1688980957
transform 1 0 37536 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_400
timestamp 1688980957
transform 1 0 37904 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_404
timestamp 1688980957
transform 1 0 38272 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_412
timestamp 1688980957
transform 1 0 39008 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_417
timestamp 1688980957
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_431
timestamp 1688980957
transform 1 0 40756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_443
timestamp 1688980957
transform 1 0 41860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_469
timestamp 1688980957
transform 1 0 44252 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_61
timestamp 1688980957
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_91
timestamp 1688980957
transform 1 0 9476 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_117
timestamp 1688980957
transform 1 0 11868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_134
timestamp 1688980957
transform 1 0 13432 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_138
timestamp 1688980957
transform 1 0 13800 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_209
timestamp 1688980957
transform 1 0 20332 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_220
timestamp 1688980957
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_234
timestamp 1688980957
transform 1 0 22632 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_242
timestamp 1688980957
transform 1 0 23368 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_251
timestamp 1688980957
transform 1 0 24196 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_271
timestamp 1688980957
transform 1 0 26036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_284
timestamp 1688980957
transform 1 0 27232 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_296
timestamp 1688980957
transform 1 0 28336 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_308
timestamp 1688980957
transform 1 0 29440 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_320
timestamp 1688980957
transform 1 0 30544 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_332
timestamp 1688980957
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_348
timestamp 1688980957
transform 1 0 33120 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_380
timestamp 1688980957
transform 1 0 36064 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_426
timestamp 1688980957
transform 1 0 40296 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_439
timestamp 1688980957
transform 1 0 41492 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 1688980957
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_463
timestamp 1688980957
transform 1 0 43700 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_469
timestamp 1688980957
transform 1 0 44252 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_73
timestamp 1688980957
transform 1 0 7820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_107
timestamp 1688980957
transform 1 0 10948 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_117
timestamp 1688980957
transform 1 0 11868 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_137
timestamp 1688980957
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_185
timestamp 1688980957
transform 1 0 18124 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_194
timestamp 1688980957
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_205
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_249
timestamp 1688980957
transform 1 0 24012 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_261
timestamp 1688980957
transform 1 0 25116 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_273
timestamp 1688980957
transform 1 0 26220 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_285
timestamp 1688980957
transform 1 0 27324 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_297
timestamp 1688980957
transform 1 0 28428 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_305
timestamp 1688980957
transform 1 0 29164 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_391
timestamp 1688980957
transform 1 0 37076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_399
timestamp 1688980957
transform 1 0 37812 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_404
timestamp 1688980957
transform 1 0 38272 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_416
timestamp 1688980957
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_432
timestamp 1688980957
transform 1 0 40848 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_444
timestamp 1688980957
transform 1 0 41952 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_456
timestamp 1688980957
transform 1 0 43056 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_468
timestamp 1688980957
transform 1 0 44160 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_110
timestamp 1688980957
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_145
timestamp 1688980957
transform 1 0 14444 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_153
timestamp 1688980957
transform 1 0 15180 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_166
timestamp 1688980957
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_177
timestamp 1688980957
transform 1 0 17388 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_188
timestamp 1688980957
transform 1 0 18400 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_202
timestamp 1688980957
transform 1 0 19688 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_212
timestamp 1688980957
transform 1 0 20608 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_239
timestamp 1688980957
transform 1 0 23092 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1688980957
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1688980957
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1688980957
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1688980957
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_355
timestamp 1688980957
transform 1 0 33764 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_359
timestamp 1688980957
transform 1 0 34132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_371
timestamp 1688980957
transform 1 0 35236 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_418
timestamp 1688980957
transform 1 0 39560 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_422
timestamp 1688980957
transform 1 0 39928 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_71
timestamp 1688980957
transform 1 0 7636 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_89
timestamp 1688980957
transform 1 0 9292 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_119
timestamp 1688980957
transform 1 0 12052 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_137
timestamp 1688980957
transform 1 0 13708 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_149
timestamp 1688980957
transform 1 0 14812 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_161
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_184
timestamp 1688980957
transform 1 0 18032 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_205
timestamp 1688980957
transform 1 0 19964 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_213
timestamp 1688980957
transform 1 0 20700 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_222
timestamp 1688980957
transform 1 0 21528 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_234
timestamp 1688980957
transform 1 0 22632 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_246
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_261
timestamp 1688980957
transform 1 0 25116 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_273
timestamp 1688980957
transform 1 0 26220 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_285
timestamp 1688980957
transform 1 0 27324 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_297
timestamp 1688980957
transform 1 0 28428 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_305
timestamp 1688980957
transform 1 0 29164 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_369
timestamp 1688980957
transform 1 0 35052 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_404
timestamp 1688980957
transform 1 0 38272 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_412
timestamp 1688980957
transform 1 0 39008 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_418
timestamp 1688980957
transform 1 0 39560 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_437
timestamp 1688980957
transform 1 0 41308 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_448
timestamp 1688980957
transform 1 0 42320 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_163
timestamp 1688980957
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_183
timestamp 1688980957
transform 1 0 17940 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_245
timestamp 1688980957
transform 1 0 23644 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_257
timestamp 1688980957
transform 1 0 24748 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_289
timestamp 1688980957
transform 1 0 27692 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_301
timestamp 1688980957
transform 1 0 28796 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_313
timestamp 1688980957
transform 1 0 29900 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_325
timestamp 1688980957
transform 1 0 31004 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_333
timestamp 1688980957
transform 1 0 31740 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_358
timestamp 1688980957
transform 1 0 34040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_390
timestamp 1688980957
transform 1 0 36984 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_409
timestamp 1688980957
transform 1 0 38732 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_413
timestamp 1688980957
transform 1 0 39100 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_441
timestamp 1688980957
transform 1 0 41676 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_469
timestamp 1688980957
transform 1 0 44252 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_49
timestamp 1688980957
transform 1 0 5612 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_62
timestamp 1688980957
transform 1 0 6808 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_74
timestamp 1688980957
transform 1 0 7912 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_82
timestamp 1688980957
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_96
timestamp 1688980957
transform 1 0 9936 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_108
timestamp 1688980957
transform 1 0 11040 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_114
timestamp 1688980957
transform 1 0 11592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_149
timestamp 1688980957
transform 1 0 14812 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_170
timestamp 1688980957
transform 1 0 16744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_191
timestamp 1688980957
transform 1 0 18676 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_225
timestamp 1688980957
transform 1 0 21804 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_237
timestamp 1688980957
transform 1 0 22908 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_249
timestamp 1688980957
transform 1 0 24012 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_262
timestamp 1688980957
transform 1 0 25208 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_274
timestamp 1688980957
transform 1 0 26312 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_286
timestamp 1688980957
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_298
timestamp 1688980957
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_306
timestamp 1688980957
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1688980957
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1688980957
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1688980957
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1688980957
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1688980957
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1688980957
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_385
timestamp 1688980957
transform 1 0 36524 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_397
timestamp 1688980957
transform 1 0 37628 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_405
timestamp 1688980957
transform 1 0 38364 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_414
timestamp 1688980957
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_432
timestamp 1688980957
transform 1 0 40848 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_444
timestamp 1688980957
transform 1 0 41952 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_456
timestamp 1688980957
transform 1 0 43056 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_468
timestamp 1688980957
transform 1 0 44160 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_121
timestamp 1688980957
transform 1 0 12236 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_146
timestamp 1688980957
transform 1 0 14536 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_150
timestamp 1688980957
transform 1 0 14904 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_184
timestamp 1688980957
transform 1 0 18032 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1688980957
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_255
timestamp 1688980957
transform 1 0 24564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_267
timestamp 1688980957
transform 1 0 25668 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1688980957
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1688980957
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_293
timestamp 1688980957
transform 1 0 28060 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_301
timestamp 1688980957
transform 1 0 28796 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_323
timestamp 1688980957
transform 1 0 30820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1688980957
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1688980957
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_349
timestamp 1688980957
transform 1 0 33212 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_359
timestamp 1688980957
transform 1 0 34132 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_371
timestamp 1688980957
transform 1 0 35236 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_382
timestamp 1688980957
transform 1 0 36248 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_390
timestamp 1688980957
transform 1 0 36984 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1688980957
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_405
timestamp 1688980957
transform 1 0 38364 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_431
timestamp 1688980957
transform 1 0 40756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_443
timestamp 1688980957
transform 1 0 41860 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 1688980957
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1688980957
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_461
timestamp 1688980957
transform 1 0 43516 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_469
timestamp 1688980957
transform 1 0 44252 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_81
timestamp 1688980957
transform 1 0 8556 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_123
timestamp 1688980957
transform 1 0 12420 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_153
timestamp 1688980957
transform 1 0 15180 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_182
timestamp 1688980957
transform 1 0 17848 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_225
timestamp 1688980957
transform 1 0 21804 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_237
timestamp 1688980957
transform 1 0 22908 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_249
timestamp 1688980957
transform 1 0 24012 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_261
timestamp 1688980957
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_272
timestamp 1688980957
transform 1 0 26128 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_284
timestamp 1688980957
transform 1 0 27232 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_296
timestamp 1688980957
transform 1 0 28336 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1688980957
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_321
timestamp 1688980957
transform 1 0 30636 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_327
timestamp 1688980957
transform 1 0 31188 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_348
timestamp 1688980957
transform 1 0 33120 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_360
timestamp 1688980957
transform 1 0 34224 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1688980957
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_377
timestamp 1688980957
transform 1 0 35788 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_400
timestamp 1688980957
transform 1 0 37904 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_412
timestamp 1688980957
transform 1 0 39008 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1688980957
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1688980957
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1688980957
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_457
timestamp 1688980957
transform 1 0 43148 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_60
timestamp 1688980957
transform 1 0 6624 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_72
timestamp 1688980957
transform 1 0 7728 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_86
timestamp 1688980957
transform 1 0 9016 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_98
timestamp 1688980957
transform 1 0 10120 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_104
timestamp 1688980957
transform 1 0 10672 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_108
timestamp 1688980957
transform 1 0 11040 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_158
timestamp 1688980957
transform 1 0 15640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_166
timestamp 1688980957
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_178
timestamp 1688980957
transform 1 0 17480 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_196
timestamp 1688980957
transform 1 0 19136 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_202
timestamp 1688980957
transform 1 0 19688 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1688980957
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1688980957
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1688980957
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1688980957
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1688980957
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1688980957
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1688980957
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1688980957
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1688980957
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1688980957
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_329
timestamp 1688980957
transform 1 0 31372 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1688980957
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1688980957
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1688980957
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1688980957
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_373
timestamp 1688980957
transform 1 0 35420 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_381
timestamp 1688980957
transform 1 0 36156 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1688980957
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1688980957
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1688980957
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1688980957
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1688980957
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1688980957
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 1688980957
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 1688980957
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1688980957
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_461
timestamp 1688980957
transform 1 0 43516 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_469
timestamp 1688980957
transform 1 0 44252 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_55
timestamp 1688980957
transform 1 0 6164 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_67
timestamp 1688980957
transform 1 0 7268 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_79
timestamp 1688980957
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_127
timestamp 1688980957
transform 1 0 12788 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_137
timestamp 1688980957
transform 1 0 13708 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_147
timestamp 1688980957
transform 1 0 14628 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_159
timestamp 1688980957
transform 1 0 15732 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_183
timestamp 1688980957
transform 1 0 17940 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_187
timestamp 1688980957
transform 1 0 18308 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_194
timestamp 1688980957
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_197
timestamp 1688980957
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_203
timestamp 1688980957
transform 1 0 19780 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_215
timestamp 1688980957
transform 1 0 20884 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_227
timestamp 1688980957
transform 1 0 21988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_239
timestamp 1688980957
transform 1 0 23092 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 1688980957
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1688980957
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1688980957
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1688980957
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1688980957
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1688980957
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1688980957
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1688980957
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_321
timestamp 1688980957
transform 1 0 30636 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_329
timestamp 1688980957
transform 1 0 31372 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_337
timestamp 1688980957
transform 1 0 32108 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_349
timestamp 1688980957
transform 1 0 33212 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_361
timestamp 1688980957
transform 1 0 34316 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1688980957
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_377
timestamp 1688980957
transform 1 0 35788 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_383
timestamp 1688980957
transform 1 0 36340 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_390
timestamp 1688980957
transform 1 0 36984 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_402
timestamp 1688980957
transform 1 0 38088 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_414
timestamp 1688980957
transform 1 0 39192 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1688980957
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1688980957
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1688980957
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1688980957
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_469
timestamp 1688980957
transform 1 0 44252 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_6
timestamp 1688980957
transform 1 0 1656 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_18
timestamp 1688980957
transform 1 0 2760 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_26
timestamp 1688980957
transform 1 0 3496 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_29
timestamp 1688980957
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_41
timestamp 1688980957
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_53
timestamp 1688980957
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_63
timestamp 1688980957
transform 1 0 6900 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_75
timestamp 1688980957
transform 1 0 8004 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_83
timestamp 1688980957
transform 1 0 8740 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_85
timestamp 1688980957
transform 1 0 8924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_97
timestamp 1688980957
transform 1 0 10028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_109
timestamp 1688980957
transform 1 0 11132 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_141
timestamp 1688980957
transform 1 0 14076 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_149
timestamp 1688980957
transform 1 0 14812 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_153
timestamp 1688980957
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_165
timestamp 1688980957
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1688980957
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_193
timestamp 1688980957
transform 1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_197
timestamp 1688980957
transform 1 0 19228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_209
timestamp 1688980957
transform 1 0 20332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_221
timestamp 1688980957
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1688980957
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_237
timestamp 1688980957
transform 1 0 22908 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_245
timestamp 1688980957
transform 1 0 23644 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_251
timestamp 1688980957
transform 1 0 24196 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_253
timestamp 1688980957
transform 1 0 24380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_265
timestamp 1688980957
transform 1 0 25484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_277
timestamp 1688980957
transform 1 0 26588 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1688980957
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1688980957
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_305
timestamp 1688980957
transform 1 0 29164 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_309
timestamp 1688980957
transform 1 0 29532 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_321
timestamp 1688980957
transform 1 0 30636 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_333
timestamp 1688980957
transform 1 0 31740 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_337
timestamp 1688980957
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_342
timestamp 1688980957
transform 1 0 32568 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_354
timestamp 1688980957
transform 1 0 33672 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_362
timestamp 1688980957
transform 1 0 34408 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_365
timestamp 1688980957
transform 1 0 34684 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_377
timestamp 1688980957
transform 1 0 35788 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_389
timestamp 1688980957
transform 1 0 36892 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1688980957
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1688980957
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_417
timestamp 1688980957
transform 1 0 39468 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_421
timestamp 1688980957
transform 1 0 39836 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_433
timestamp 1688980957
transform 1 0 40940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_440
timestamp 1688980957
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1688980957
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_461
timestamp 1688980957
transform 1 0 43516 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_469
timestamp 1688980957
transform 1 0 44252 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 33396 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 38732 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 41584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 7636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 34500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 43148 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 29072 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 25392 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 9660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 8740 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 8096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 4784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 39836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 5336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 38732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 27232 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 25116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 25852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 25208 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold38 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 44252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 18492 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 18308 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 13984 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 13248 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 17296 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 21804 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 19136 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 22816 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 24104 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 23000 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 23736 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 13064 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 12236 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 17112 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 16468 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 11592 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 10672 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 43332 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 43516 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 18768 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 18032 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 23368 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 22448 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 23828 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 18676 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 23092 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 23276 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 11868 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 10948 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold71
timestamp 1688980957
transform -1 0 37352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  hold72
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 20608 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 19964 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 12696 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 12696 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 37260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 17480 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 17204 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 13708 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 14444 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 35604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 38088 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 37352 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 39652 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 15548 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 15364 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 44344 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 42044 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 37444 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 37996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 36892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 27692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 43608 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 41860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 39928 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 39192 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 42320 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 41308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 31188 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 23920 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 21160 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold107
timestamp 1688980957
transform -1 0 35420 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 43976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 41492 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 35420 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 41860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 40848 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 28428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 38732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 21804 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 32108 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 35052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 43884 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 44160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 15732 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 31096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 30728 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 29532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 14812 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 28244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 19044 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 17848 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 38640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 37996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 36616 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 21620 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 36156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 35788 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 26036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 24564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform -1 0 40940 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 10672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 26220 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 35880 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform -1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 36524 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 40480 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 36248 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 31372 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 36156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform 1 0 41952 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 37076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 36892 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform -1 0 40572 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform -1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 35696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform 1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 32660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 42596 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 42688 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform -1 0 34132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 23368 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform -1 0 36708 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 39744 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform -1 0 41308 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 28888 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 34408 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 39284 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform 1 0 32384 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 25116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 44344 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform -1 0 43516 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 32200 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 40572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 43148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform -1 0 30544 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 9844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 41308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 39744 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 34960 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 39744 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 40572 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 38548 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform -1 0 36708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform -1 0 40572 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 43240 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 37076 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 34960 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 18216 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 13892 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 37628 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 19228 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform 1 0 27600 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 9108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 16468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform -1 0 32844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 9200 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 13064 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 8096 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform -1 0 16192 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 16560 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 21804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 15916 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform -1 0 17388 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 13984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 17388 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 18308 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 11684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 11040 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform -1 0 17480 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 17848 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 24380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 41952 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 37076 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 27508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 12788 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 15640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 19228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 14812 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 37168 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 21160 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 21988 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform -1 0 9660 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 7084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 38824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 20792 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 18768 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 16100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform -1 0 25116 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 18952 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 11684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  input1
timestamp 1688980957
transform -1 0 44344 0 1 43520
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 24196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 44068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 1656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 44068 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 15180 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 44068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 1656 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 32292 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1688980957
transform 1 0 6532 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1688980957
transform 1 0 43976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 44620 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 44620 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 44620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 44620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 44620 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 44620 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 44620 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 44620 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 44620 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 44620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 44620 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 44620 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 44620 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 44620 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 44620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 44620 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 44620 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 44620 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 44620 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 44620 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 44620 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 44620 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 44620 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 44620 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 44620 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 44620 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 44620 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 44620 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 44620 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 44620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 44620 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 44620 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 44620 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 44620 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 44620 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 44620 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 44620 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 44620 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 44620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 44620 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 44620 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 44620 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 44620 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 44620 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 44620 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 44620 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 44620 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 44620 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 44620 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 44620 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 44620 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1688980957
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1688980957
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1688980957
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1688980957
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1688980957
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1688980957
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1688980957
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1688980957
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1688980957
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1688980957
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1688980957
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1688980957
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1688980957
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1688980957
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1688980957
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1688980957
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1688980957
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1688980957
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1688980957
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1688980957
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1688980957
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1688980957
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1688980957
transform 1 0 3680 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1688980957
transform 1 0 8832 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1688980957
transform 1 0 13984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1688980957
transform 1 0 19136 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1688980957
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1688980957
transform 1 0 24288 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1688980957
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1688980957
transform 1 0 29440 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1688980957
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1688980957
transform 1 0 34592 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1688980957
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1688980957
transform 1 0 39744 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1688980957
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  wire21
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
<< labels >>
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 44933 43528 45733 43648 0 FreeSans 480 0 0 0 cs
port 1 nsew signal input
flabel metal2 s 41234 47077 41290 47877 0 FreeSans 224 90 0 0 gpio[0]
port 2 nsew signal input
flabel metal2 s 23846 47077 23902 47877 0 FreeSans 224 90 0 0 gpio[10]
port 3 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpio[11]
port 4 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpio[12]
port 5 nsew signal input
flabel metal3 s 44933 6808 45733 6928 0 FreeSans 480 0 0 0 gpio[13]
port 6 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 gpio[14]
port 7 nsew signal input
flabel metal3 s 44933 34008 45733 34128 0 FreeSans 480 0 0 0 gpio[15]
port 8 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio[16]
port 9 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio[1]
port 10 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 gpio[2]
port 11 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio[3]
port 12 nsew signal input
flabel metal2 s 14830 47077 14886 47877 0 FreeSans 224 90 0 0 gpio[4]
port 13 nsew signal input
flabel metal3 s 44933 25168 45733 25288 0 FreeSans 480 0 0 0 gpio[5]
port 14 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 gpio[6]
port 15 nsew signal input
flabel metal2 s 32218 47077 32274 47877 0 FreeSans 224 90 0 0 gpio[7]
port 16 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 gpio[8]
port 17 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gpio[9]
port 18 nsew signal input
flabel metal2 s 6458 47077 6514 47877 0 FreeSans 224 90 0 0 nrst
port 19 nsew signal input
flabel metal3 s 44933 15648 45733 15768 0 FreeSans 480 0 0 0 pwm
port 20 nsew signal tristate
flabel metal4 s 4208 2128 4528 45744 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 34928 2128 35248 45744 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 19568 2128 19888 45744 0 FreeSans 1920 90 0 0 vssd1
port 22 nsew ground bidirectional
rlabel metal1 22862 45152 22862 45152 0 vccd1
rlabel metal1 22862 45696 22862 45696 0 vssd1
rlabel metal1 23782 2924 23782 2924 0 _0000_
rlabel metal1 21528 3570 21528 3570 0 _0001_
rlabel metal1 24334 4522 24334 4522 0 _0002_
rlabel metal1 33396 23834 33396 23834 0 _0003_
rlabel metal1 35282 21896 35282 21896 0 _0004_
rlabel metal1 34960 20502 34960 20502 0 _0005_
rlabel metal1 35788 18190 35788 18190 0 _0006_
rlabel metal1 33350 14926 33350 14926 0 _0007_
rlabel metal1 32798 15538 32798 15538 0 _0008_
rlabel metal1 28612 15538 28612 15538 0 _0009_
rlabel metal2 31142 18972 31142 18972 0 _0010_
rlabel metal1 27508 19278 27508 19278 0 _0011_
rlabel metal1 28336 21658 28336 21658 0 _0012_
rlabel metal1 29624 22746 29624 22746 0 _0013_
rlabel metal1 32798 24718 32798 24718 0 _0014_
rlabel metal1 28658 27030 28658 27030 0 _0015_
rlabel metal1 33166 26010 33166 26010 0 _0016_
rlabel metal1 28934 28152 28934 28152 0 _0017_
rlabel metal1 33488 27642 33488 27642 0 _0018_
rlabel metal1 32246 30328 32246 30328 0 _0019_
rlabel metal1 35696 30362 35696 30362 0 _0020_
rlabel metal1 37766 33422 37766 33422 0 _0021_
rlabel metal2 36110 35156 36110 35156 0 _0022_
rlabel metal1 32706 38794 32706 38794 0 _0023_
rlabel metal1 31970 39066 31970 39066 0 _0024_
rlabel metal1 30268 37978 30268 37978 0 _0025_
rlabel metal1 28934 35768 28934 35768 0 _0026_
rlabel metal1 30360 33422 30360 33422 0 _0027_
rlabel metal2 29578 31450 29578 31450 0 _0028_
rlabel metal1 37204 31994 37204 31994 0 _0029_
rlabel metal1 38870 30906 38870 30906 0 _0030_
rlabel metal1 39054 30328 39054 30328 0 _0031_
rlabel metal1 40066 29818 40066 29818 0 _0032_
rlabel metal1 39606 27574 39606 27574 0 _0033_
rlabel metal1 37766 27098 37766 27098 0 _0034_
rlabel metal1 36156 28186 36156 28186 0 _0035_
rlabel metal1 35006 26860 35006 26860 0 _0036_
rlabel metal1 27738 30362 27738 30362 0 _0037_
rlabel metal1 26634 30770 26634 30770 0 _0038_
rlabel metal1 25254 31994 25254 31994 0 _0039_
rlabel metal1 25898 32980 25898 32980 0 _0040_
rlabel metal2 25070 34612 25070 34612 0 _0041_
rlabel metal2 24426 36788 24426 36788 0 _0042_
rlabel metal1 20240 36890 20240 36890 0 _0043_
rlabel metal1 17894 37740 17894 37740 0 _0044_
rlabel metal1 14214 38522 14214 38522 0 _0045_
rlabel metal2 12098 39508 12098 39508 0 _0046_
rlabel metal1 13616 40698 13616 40698 0 _0047_
rlabel metal1 14168 41650 14168 41650 0 _0048_
rlabel metal1 15410 42330 15410 42330 0 _0049_
rlabel metal2 17342 41956 17342 41956 0 _0050_
rlabel metal1 19136 41650 19136 41650 0 _0051_
rlabel metal2 22126 41956 22126 41956 0 _0052_
rlabel metal2 24150 40324 24150 40324 0 _0053_
rlabel metal1 24518 39066 24518 39066 0 _0054_
rlabel metal1 34914 26350 34914 26350 0 _0055_
rlabel metal1 26772 39474 26772 39474 0 _0056_
rlabel metal1 28336 38522 28336 38522 0 _0057_
rlabel metal1 26680 37298 26680 37298 0 _0058_
rlabel metal1 26772 36210 26772 36210 0 _0059_
rlabel metal1 27048 34034 27048 34034 0 _0060_
rlabel metal2 42228 30906 42228 30906 0 _0061_
rlabel metal1 42504 28458 42504 28458 0 _0062_
rlabel metal2 44022 27098 44022 27098 0 _0063_
rlabel metal1 43700 25330 43700 25330 0 _0064_
rlabel metal1 40618 24106 40618 24106 0 _0065_
rlabel metal1 39422 23800 39422 23800 0 _0066_
rlabel metal1 37352 23154 37352 23154 0 _0067_
rlabel metal1 36524 19890 36524 19890 0 _0068_
rlabel metal1 40894 31654 40894 31654 0 _0069_
rlabel metal2 41906 30396 41906 30396 0 _0070_
rlabel metal2 41722 27778 41722 27778 0 _0071_
rlabel metal1 41492 26894 41492 26894 0 _0072_
rlabel metal1 40618 25466 40618 25466 0 _0073_
rlabel metal1 39514 25330 39514 25330 0 _0074_
rlabel metal1 37628 25874 37628 25874 0 _0075_
rlabel metal1 36616 26418 36616 26418 0 _0076_
rlabel metal1 18308 19414 18308 19414 0 _0077_
rlabel metal1 22632 19278 22632 19278 0 _0078_
rlabel metal1 16284 17578 16284 17578 0 _0079_
rlabel metal2 20838 19992 20838 19992 0 _0080_
rlabel metal2 18722 16932 18722 16932 0 _0081_
rlabel metal1 23828 16014 23828 16014 0 _0082_
rlabel metal1 27416 14314 27416 14314 0 _0083_
rlabel metal2 14398 17306 14398 17306 0 _0084_
rlabel metal1 24748 18326 24748 18326 0 _0085_
rlabel metal1 10350 18394 10350 18394 0 _0086_
rlabel metal1 12788 18326 12788 18326 0 _0087_
rlabel metal1 10527 20026 10527 20026 0 _0088_
rlabel metal1 13478 21454 13478 21454 0 _0089_
rlabel via1 15495 20026 15495 20026 0 _0090_
rlabel metal1 22586 24718 22586 24718 0 _0091_
rlabel metal1 24794 27302 24794 27302 0 _0092_
rlabel metal1 24968 27642 24968 27642 0 _0093_
rlabel metal1 23644 25466 23644 25466 0 _0094_
rlabel metal1 17986 18394 17986 18394 0 _0095_
rlabel metal2 20746 18020 20746 18020 0 _0096_
rlabel metal1 16652 16218 16652 16218 0 _0097_
rlabel metal1 20470 15130 20470 15130 0 _0098_
rlabel metal1 18354 14926 18354 14926 0 _0099_
rlabel metal1 22678 15402 22678 15402 0 _0100_
rlabel metal2 25254 14756 25254 14756 0 _0101_
rlabel metal1 13662 15674 13662 15674 0 _0102_
rlabel metal2 22218 16932 22218 16932 0 _0103_
rlabel metal1 10534 17306 10534 17306 0 _0104_
rlabel metal1 11822 16218 11822 16218 0 _0105_
rlabel metal1 10718 15130 10718 15130 0 _0106_
rlabel metal1 12788 19890 12788 19890 0 _0107_
rlabel metal1 15180 18938 15180 18938 0 _0108_
rlabel metal1 21567 22202 21567 22202 0 _0109_
rlabel metal1 22954 20978 22954 20978 0 _0110_
rlabel metal1 22908 22746 22908 22746 0 _0111_
rlabel metal2 22034 25500 22034 25500 0 _0112_
rlabel metal1 13984 23290 13984 23290 0 _0113_
rlabel metal1 20194 23800 20194 23800 0 _0114_
rlabel metal1 15778 21658 15778 21658 0 _0115_
rlabel metal1 20194 21114 20194 21114 0 _0116_
rlabel metal1 18308 20502 18308 20502 0 _0117_
rlabel metal1 16744 22678 16744 22678 0 _0118_
rlabel metal1 17894 23834 17894 23834 0 _0119_
rlabel metal2 12466 21794 12466 21794 0 _0120_
rlabel metal1 19918 22406 19918 22406 0 _0121_
rlabel metal1 10389 22202 10389 22202 0 _0122_
rlabel metal1 12006 23834 12006 23834 0 _0123_
rlabel metal1 9798 22712 9798 22712 0 _0124_
rlabel metal1 11132 24650 11132 24650 0 _0125_
rlabel metal1 14306 24378 14306 24378 0 _0126_
rlabel metal1 16928 24378 16928 24378 0 _0127_
rlabel metal1 22724 30906 22724 30906 0 _0128_
rlabel metal1 24334 29818 24334 29818 0 _0129_
rlabel metal2 22494 30362 22494 30362 0 _0130_
rlabel metal1 19826 25466 19826 25466 0 _0131_
rlabel metal1 16974 27064 16974 27064 0 _0132_
rlabel metal1 23552 28118 23552 28118 0 _0133_
rlabel metal1 23782 34034 23782 34034 0 _0134_
rlabel metal1 16376 29274 16376 29274 0 _0135_
rlabel metal1 23644 36346 23644 36346 0 _0136_
rlabel metal1 18308 34510 18308 34510 0 _0137_
rlabel metal1 17572 36686 17572 36686 0 _0138_
rlabel metal1 12834 37298 12834 37298 0 _0139_
rlabel metal1 9982 38386 9982 38386 0 _0140_
rlabel metal1 10488 39950 10488 39950 0 _0141_
rlabel metal1 11730 43214 11730 43214 0 _0142_
rlabel metal1 13340 42874 13340 42874 0 _0143_
rlabel metal1 16422 43180 16422 43180 0 _0144_
rlabel metal1 18814 43826 18814 43826 0 _0145_
rlabel metal1 19504 40562 19504 40562 0 _0146_
rlabel metal1 22816 41106 22816 41106 0 _0147_
rlabel metal2 22126 38828 22126 38828 0 _0148_
rlabel metal1 12006 25942 12006 25942 0 _0149_
rlabel metal1 14352 25466 14352 25466 0 _0150_
rlabel metal1 14122 28118 14122 28118 0 _0151_
rlabel metal1 16744 32470 16744 32470 0 _0152_
rlabel metal1 11079 27642 11079 27642 0 _0153_
rlabel metal2 14766 34340 14766 34340 0 _0154_
rlabel metal2 15962 33048 15962 33048 0 _0155_
rlabel metal2 15318 37332 15318 37332 0 _0156_
rlabel metal1 7038 37434 7038 37434 0 _0157_
rlabel metal1 6900 38250 6900 38250 0 _0158_
rlabel metal1 7268 39610 7268 39610 0 _0159_
rlabel metal1 10764 41242 10764 41242 0 _0160_
rlabel metal1 9384 42262 9384 42262 0 _0161_
rlabel metal1 7590 41786 7590 41786 0 _0162_
rlabel metal1 15870 40562 15870 40562 0 _0163_
rlabel metal1 17112 40086 17112 40086 0 _0164_
rlabel metal1 14260 39338 14260 39338 0 _0165_
rlabel metal1 15042 35802 15042 35802 0 _0166_
rlabel metal1 21022 26418 21022 26418 0 _0167_
rlabel metal1 17434 27336 17434 27336 0 _0168_
rlabel metal1 21988 27098 21988 27098 0 _0169_
rlabel metal1 23598 32946 23598 32946 0 _0170_
rlabel metal2 18078 29682 18078 29682 0 _0171_
rlabel metal2 22126 35938 22126 35938 0 _0172_
rlabel metal1 19320 34986 19320 34986 0 _0173_
rlabel metal1 20985 36346 20985 36346 0 _0174_
rlabel metal1 12512 35802 12512 35802 0 _0175_
rlabel metal1 10120 36278 10120 36278 0 _0176_
rlabel metal1 9982 39066 9982 39066 0 _0177_
rlabel metal1 10672 44506 10672 44506 0 _0178_
rlabel metal1 13386 44472 13386 44472 0 _0179_
rlabel metal1 16238 44914 16238 44914 0 _0180_
rlabel metal1 18952 43690 18952 43690 0 _0181_
rlabel metal1 19320 39338 19320 39338 0 _0182_
rlabel metal2 21114 40426 21114 40426 0 _0183_
rlabel metal1 20746 37978 20746 37978 0 _0184_
rlabel metal1 6670 5134 6670 5134 0 _0185_
rlabel metal2 7682 6426 7682 6426 0 _0186_
rlabel metal1 7314 4046 7314 4046 0 _0187_
rlabel metal1 7912 8466 7912 8466 0 _0188_
rlabel metal1 7728 11322 7728 11322 0 _0189_
rlabel metal1 8464 12750 8464 12750 0 _0190_
rlabel metal1 33718 20978 33718 20978 0 _0191_
rlabel metal1 33580 20774 33580 20774 0 _0192_
rlabel metal1 33212 20910 33212 20910 0 _0193_
rlabel metal1 34086 20842 34086 20842 0 _0194_
rlabel metal1 35006 20944 35006 20944 0 _0195_
rlabel metal1 34730 20910 34730 20910 0 _0196_
rlabel metal1 34730 19380 34730 19380 0 _0197_
rlabel metal2 32982 20570 32982 20570 0 _0198_
rlabel metal1 33442 20366 33442 20366 0 _0199_
rlabel metal1 34270 19380 34270 19380 0 _0200_
rlabel metal1 34270 17204 34270 17204 0 _0201_
rlabel metal1 34270 19210 34270 19210 0 _0202_
rlabel metal2 35834 18938 35834 18938 0 _0203_
rlabel metal1 36018 18768 36018 18768 0 _0204_
rlabel metal1 33166 16184 33166 16184 0 _0205_
rlabel metal1 33902 20468 33902 20468 0 _0206_
rlabel metal1 34408 17170 34408 17170 0 _0207_
rlabel metal1 34362 16626 34362 16626 0 _0208_
rlabel metal1 27186 17748 27186 17748 0 _0209_
rlabel metal1 27791 17170 27791 17170 0 _0210_
rlabel metal1 32338 17782 32338 17782 0 _0211_
rlabel metal1 34960 16490 34960 16490 0 _0212_
rlabel metal2 33902 16252 33902 16252 0 _0213_
rlabel metal1 33810 16116 33810 16116 0 _0214_
rlabel metal1 33672 17170 33672 17170 0 _0215_
rlabel metal1 33718 15402 33718 15402 0 _0216_
rlabel metal1 32752 16558 32752 16558 0 _0217_
rlabel metal2 26082 17578 26082 17578 0 _0218_
rlabel metal1 26818 17068 26818 17068 0 _0219_
rlabel metal1 32890 16762 32890 16762 0 _0220_
rlabel metal1 33074 15674 33074 15674 0 _0221_
rlabel metal2 33350 15878 33350 15878 0 _0222_
rlabel metal1 30958 16116 30958 16116 0 _0223_
rlabel metal1 26082 17816 26082 17816 0 _0224_
rlabel metal1 27508 16626 27508 16626 0 _0225_
rlabel viali 31132 16082 31132 16082 0 _0226_
rlabel metal1 30636 16558 30636 16558 0 _0227_
rlabel metal1 31648 16218 31648 16218 0 _0228_
rlabel metal1 31096 16422 31096 16422 0 _0229_
rlabel metal1 33718 16762 33718 16762 0 _0230_
rlabel metal1 33626 17034 33626 17034 0 _0231_
rlabel metal2 32430 17340 32430 17340 0 _0232_
rlabel metal1 32982 17136 32982 17136 0 _0233_
rlabel metal1 32246 17000 32246 17000 0 _0234_
rlabel metal2 29578 16320 29578 16320 0 _0235_
rlabel metal1 29486 15980 29486 15980 0 _0236_
rlabel metal1 30084 17102 30084 17102 0 _0237_
rlabel metal1 26542 17714 26542 17714 0 _0238_
rlabel metal1 29210 17612 29210 17612 0 _0239_
rlabel metal1 30498 17646 30498 17646 0 _0240_
rlabel metal1 29578 17714 29578 17714 0 _0241_
rlabel metal1 29854 17782 29854 17782 0 _0242_
rlabel metal1 30176 17306 30176 17306 0 _0243_
rlabel metal1 31096 18190 31096 18190 0 _0244_
rlabel metal2 29578 17476 29578 17476 0 _0245_
rlabel metal1 29394 19788 29394 19788 0 _0246_
rlabel metal1 30728 20910 30728 20910 0 _0247_
rlabel metal1 26082 21590 26082 21590 0 _0248_
rlabel metal1 25944 19822 25944 19822 0 _0249_
rlabel metal1 25944 20978 25944 20978 0 _0250_
rlabel metal1 28750 20468 28750 20468 0 _0251_
rlabel metal1 29762 20808 29762 20808 0 _0252_
rlabel metal1 29992 20842 29992 20842 0 _0253_
rlabel metal2 29578 20638 29578 20638 0 _0254_
rlabel metal1 28566 19958 28566 19958 0 _0255_
rlabel metal1 28244 19822 28244 19822 0 _0256_
rlabel metal1 25438 19822 25438 19822 0 _0257_
rlabel metal1 28428 20434 28428 20434 0 _0258_
rlabel metal2 28934 20162 28934 20162 0 _0259_
rlabel metal2 29946 20128 29946 20128 0 _0260_
rlabel metal1 28888 20978 28888 20978 0 _0261_
rlabel metal1 28934 21114 28934 21114 0 _0262_
rlabel metal1 28658 21046 28658 21046 0 _0263_
rlabel metal1 25392 21998 25392 21998 0 _0264_
rlabel metal1 25162 22746 25162 22746 0 _0265_
rlabel metal1 27232 23154 27232 23154 0 _0266_
rlabel metal1 32154 23120 32154 23120 0 _0267_
rlabel metal1 30176 20026 30176 20026 0 _0268_
rlabel metal1 30498 20434 30498 20434 0 _0269_
rlabel metal1 32338 23154 32338 23154 0 _0270_
rlabel metal2 30314 23834 30314 23834 0 _0271_
rlabel metal1 29578 22644 29578 22644 0 _0272_
rlabel metal1 25714 22542 25714 22542 0 _0273_
rlabel metal1 26312 22746 26312 22746 0 _0274_
rlabel metal1 29486 22066 29486 22066 0 _0275_
rlabel metal1 29900 24174 29900 24174 0 _0276_
rlabel metal1 30544 24174 30544 24174 0 _0277_
rlabel metal1 31050 23732 31050 23732 0 _0278_
rlabel metal1 31142 23834 31142 23834 0 _0279_
rlabel metal1 28612 22746 28612 22746 0 _0280_
rlabel metal1 29486 24038 29486 24038 0 _0281_
rlabel metal1 30498 24242 30498 24242 0 _0282_
rlabel metal1 31280 24378 31280 24378 0 _0283_
rlabel metal1 30360 25194 30360 25194 0 _0284_
rlabel metal2 26082 23392 26082 23392 0 _0285_
rlabel metal2 27738 25092 27738 25092 0 _0286_
rlabel metal1 28566 25296 28566 25296 0 _0287_
rlabel metal2 29210 25874 29210 25874 0 _0288_
rlabel metal1 29348 25262 29348 25262 0 _0289_
rlabel metal1 29946 26384 29946 26384 0 _0290_
rlabel metal1 29578 23766 29578 23766 0 _0291_
rlabel metal1 29854 25670 29854 25670 0 _0292_
rlabel metal1 29440 26010 29440 26010 0 _0293_
rlabel metal1 29026 26928 29026 26928 0 _0294_
rlabel metal1 28566 25874 28566 25874 0 _0295_
rlabel metal1 26542 25364 26542 25364 0 _0296_
rlabel metal1 27554 25874 27554 25874 0 _0297_
rlabel metal1 28520 26010 28520 26010 0 _0298_
rlabel metal1 28980 25942 28980 25942 0 _0299_
rlabel metal1 29762 26316 29762 26316 0 _0300_
rlabel metal1 30314 26010 30314 26010 0 _0301_
rlabel metal2 32154 26180 32154 26180 0 _0302_
rlabel metal1 32614 26962 32614 26962 0 _0303_
rlabel metal2 25714 25126 25714 25126 0 _0304_
rlabel metal1 31510 27030 31510 27030 0 _0305_
rlabel metal1 32108 28050 32108 28050 0 _0306_
rlabel metal2 32338 27574 32338 27574 0 _0307_
rlabel metal1 32292 28186 32292 28186 0 _0308_
rlabel metal1 28842 26316 28842 26316 0 _0309_
rlabel metal1 29486 26350 29486 26350 0 _0310_
rlabel metal2 31142 27302 31142 27302 0 _0311_
rlabel metal2 30498 28288 30498 28288 0 _0312_
rlabel metal1 30774 28186 30774 28186 0 _0313_
rlabel metal1 27784 28526 27784 28526 0 _0314_
rlabel metal1 27784 28662 27784 28662 0 _0315_
rlabel metal1 29026 28560 29026 28560 0 _0316_
rlabel metal2 31970 28492 31970 28492 0 _0317_
rlabel metal1 31556 29138 31556 29138 0 _0318_
rlabel metal1 31004 29138 31004 29138 0 _0319_
rlabel metal2 32154 28832 32154 28832 0 _0320_
rlabel metal1 32982 28050 32982 28050 0 _0321_
rlabel metal1 32752 27438 32752 27438 0 _0322_
rlabel metal1 33810 29138 33810 29138 0 _0323_
rlabel metal1 27278 29036 27278 29036 0 _0324_
rlabel metal1 33074 29138 33074 29138 0 _0325_
rlabel metal1 34086 30294 34086 30294 0 _0326_
rlabel metal1 33810 29274 33810 29274 0 _0327_
rlabel metal2 34454 29852 34454 29852 0 _0328_
rlabel metal1 31970 28526 31970 28526 0 _0329_
rlabel metal1 33028 28458 33028 28458 0 _0330_
rlabel metal1 32660 30294 32660 30294 0 _0331_
rlabel metal1 32430 30294 32430 30294 0 _0332_
rlabel metal1 32729 38998 32729 38998 0 _0333_
rlabel metal1 38272 26962 38272 26962 0 _0334_
rlabel metal1 34270 30158 34270 30158 0 _0335_
rlabel metal1 27646 30056 27646 30056 0 _0336_
rlabel metal2 29486 30498 29486 30498 0 _0337_
rlabel via1 33166 30243 33166 30243 0 _0338_
rlabel metal1 34408 30906 34408 30906 0 _0339_
rlabel metal1 34776 30362 34776 30362 0 _0340_
rlabel metal1 35098 30260 35098 30260 0 _0341_
rlabel metal1 33856 36142 33856 36142 0 _0342_
rlabel metal1 34362 32470 34362 32470 0 _0343_
rlabel metal1 35466 32538 35466 32538 0 _0344_
rlabel metal1 34086 34034 34086 34034 0 _0345_
rlabel metal1 33994 32878 33994 32878 0 _0346_
rlabel metal1 33672 30294 33672 30294 0 _0347_
rlabel metal1 34178 32844 34178 32844 0 _0348_
rlabel metal1 34776 32946 34776 32946 0 _0349_
rlabel metal1 36041 33490 36041 33490 0 _0350_
rlabel metal1 34086 33932 34086 33932 0 _0351_
rlabel metal1 34868 33082 34868 33082 0 _0352_
rlabel metal1 35282 34170 35282 34170 0 _0353_
rlabel metal1 34500 33490 34500 33490 0 _0354_
rlabel metal1 32706 35734 32706 35734 0 _0355_
rlabel viali 33442 33490 33442 33490 0 _0356_
rlabel metal1 33718 32538 33718 32538 0 _0357_
rlabel metal1 34132 33490 34132 33490 0 _0358_
rlabel metal1 33534 36720 33534 36720 0 _0359_
rlabel metal1 34086 36720 34086 36720 0 _0360_
rlabel metal1 34040 36278 34040 36278 0 _0361_
rlabel metal1 33672 37230 33672 37230 0 _0362_
rlabel metal1 33166 38930 33166 38930 0 _0363_
rlabel metal1 33672 38522 33672 38522 0 _0364_
rlabel metal1 33442 36890 33442 36890 0 _0365_
rlabel metal1 33948 36346 33948 36346 0 _0366_
rlabel metal1 33672 37162 33672 37162 0 _0367_
rlabel metal1 32568 38522 32568 38522 0 _0368_
rlabel metal1 32338 38828 32338 38828 0 _0369_
rlabel metal1 33350 36686 33350 36686 0 _0370_
rlabel metal1 32890 36788 32890 36788 0 _0371_
rlabel metal2 31786 35428 31786 35428 0 _0372_
rlabel metal1 31970 35156 31970 35156 0 _0373_
rlabel metal2 32706 36516 32706 36516 0 _0374_
rlabel metal1 32246 36244 32246 36244 0 _0375_
rlabel metal2 32982 37128 32982 37128 0 _0376_
rlabel metal2 30038 35938 30038 35938 0 _0377_
rlabel metal1 31970 36108 31970 36108 0 _0378_
rlabel metal1 29946 36210 29946 36210 0 _0379_
rlabel metal1 29854 36074 29854 36074 0 _0380_
rlabel metal1 32660 36006 32660 36006 0 _0381_
rlabel metal2 32614 34850 32614 34850 0 _0382_
rlabel metal1 31050 34170 31050 34170 0 _0383_
rlabel metal1 30590 34170 30590 34170 0 _0384_
rlabel metal2 32338 34238 32338 34238 0 _0385_
rlabel metal1 31326 33388 31326 33388 0 _0386_
rlabel metal1 32384 33490 32384 33490 0 _0387_
rlabel metal1 31970 33456 31970 33456 0 _0388_
rlabel metal1 31280 32402 31280 32402 0 _0389_
rlabel metal2 30958 32572 30958 32572 0 _0390_
rlabel metal1 31234 31824 31234 31824 0 _0391_
rlabel metal1 29854 31858 29854 31858 0 _0392_
rlabel via1 29762 31800 29762 31800 0 _0393_
rlabel metal1 31096 31110 31096 31110 0 _0394_
rlabel metal1 34408 31790 34408 31790 0 _0395_
rlabel metal2 13754 26384 13754 26384 0 _0396_
rlabel metal1 19780 25262 19780 25262 0 _0397_
rlabel metal1 16468 37230 16468 37230 0 _0398_
rlabel metal1 17434 28050 17434 28050 0 _0399_
rlabel metal1 19366 36788 19366 36788 0 _0400_
rlabel metal1 19412 27914 19412 27914 0 _0401_
rlabel metal1 24058 32878 24058 32878 0 _0402_
rlabel metal1 16928 29138 16928 29138 0 _0403_
rlabel metal1 17756 35258 17756 35258 0 _0404_
rlabel metal1 12512 38998 12512 38998 0 _0405_
rlabel metal1 18538 34646 18538 34646 0 _0406_
rlabel metal1 16882 37434 16882 37434 0 _0407_
rlabel metal1 13064 37842 13064 37842 0 _0408_
rlabel metal2 12742 38692 12742 38692 0 _0409_
rlabel metal1 11822 40154 11822 40154 0 _0410_
rlabel metal1 16422 18666 16422 18666 0 _0411_
rlabel metal1 12742 42874 12742 42874 0 _0412_
rlabel metal1 13662 42636 13662 42636 0 _0413_
rlabel metal1 16882 42330 16882 42330 0 _0414_
rlabel metal1 18354 42228 18354 42228 0 _0415_
rlabel metal1 19366 41174 19366 41174 0 _0416_
rlabel metal2 20746 39780 20746 39780 0 _0417_
rlabel metal1 19504 38998 19504 38998 0 _0418_
rlabel metal2 27002 39372 27002 39372 0 _0419_
rlabel metal1 28750 38216 28750 38216 0 _0420_
rlabel metal2 28566 38794 28566 38794 0 _0421_
rlabel metal1 28474 36788 28474 36788 0 _0422_
rlabel metal1 27830 36754 27830 36754 0 _0423_
rlabel metal1 27968 36686 27968 36686 0 _0424_
rlabel metal1 27462 35462 27462 35462 0 _0425_
rlabel metal1 27730 35802 27730 35802 0 _0426_
rlabel metal1 27140 35802 27140 35802 0 _0427_
rlabel metal1 27646 34646 27646 34646 0 _0428_
rlabel metal1 42274 32402 42274 32402 0 _0429_
rlabel metal1 42412 29138 42412 29138 0 _0430_
rlabel metal1 44206 27472 44206 27472 0 _0431_
rlabel metal1 43240 25874 43240 25874 0 _0432_
rlabel metal1 40618 23834 40618 23834 0 _0433_
rlabel metal1 38962 24174 38962 24174 0 _0434_
rlabel metal2 37582 23460 37582 23460 0 _0435_
rlabel metal2 17250 16932 17250 16932 0 _0436_
rlabel metal1 37122 20434 37122 20434 0 _0437_
rlabel metal1 37766 34578 37766 34578 0 _0438_
rlabel metal1 37996 34714 37996 34714 0 _0439_
rlabel metal1 37490 30158 37490 30158 0 _0440_
rlabel metal1 37674 29274 37674 29274 0 _0441_
rlabel metal1 38272 30362 38272 30362 0 _0442_
rlabel metal1 38272 30906 38272 30906 0 _0443_
rlabel metal1 18952 18938 18952 18938 0 _0444_
rlabel metal1 22310 18938 22310 18938 0 _0445_
rlabel metal1 16652 17306 16652 17306 0 _0446_
rlabel metal1 20976 19482 20976 19482 0 _0447_
rlabel metal1 19090 16558 19090 16558 0 _0448_
rlabel metal1 24150 16558 24150 16558 0 _0449_
rlabel metal1 26864 15674 26864 15674 0 _0450_
rlabel metal2 14582 17204 14582 17204 0 _0451_
rlabel metal2 23138 18564 23138 18564 0 _0452_
rlabel metal1 19458 18224 19458 18224 0 _0453_
rlabel metal1 10810 18258 10810 18258 0 _0454_
rlabel metal1 12834 17850 12834 17850 0 _0455_
rlabel metal1 11224 20434 11224 20434 0 _0456_
rlabel metal1 13616 21114 13616 21114 0 _0457_
rlabel metal1 15456 20434 15456 20434 0 _0458_
rlabel metal1 22172 24378 22172 24378 0 _0459_
rlabel metal1 24610 27098 24610 27098 0 _0460_
rlabel metal1 24334 27642 24334 27642 0 _0461_
rlabel metal1 23920 25262 23920 25262 0 _0462_
rlabel metal1 22724 11730 22724 11730 0 _0463_
rlabel metal1 22034 7922 22034 7922 0 _0464_
rlabel metal1 14306 6120 14306 6120 0 _0465_
rlabel metal2 15502 4505 15502 4505 0 _0466_
rlabel metal1 6670 9010 6670 9010 0 _0467_
rlabel metal1 9430 3400 9430 3400 0 _0468_
rlabel metal1 11546 4114 11546 4114 0 _0469_
rlabel metal1 10626 7412 10626 7412 0 _0470_
rlabel via1 11096 4522 11096 4522 0 _0471_
rlabel metal1 14812 12886 14812 12886 0 _0472_
rlabel metal1 7406 6698 7406 6698 0 _0473_
rlabel metal1 15180 7378 15180 7378 0 _0474_
rlabel metal1 19044 7854 19044 7854 0 _0475_
rlabel metal1 11546 6290 11546 6290 0 _0476_
rlabel via1 13754 8466 13754 8466 0 _0477_
rlabel metal2 11270 4998 11270 4998 0 _0478_
rlabel metal1 13432 8942 13432 8942 0 _0479_
rlabel metal2 19550 11305 19550 11305 0 _0480_
rlabel metal2 16054 8432 16054 8432 0 _0481_
rlabel metal1 19964 7922 19964 7922 0 _0482_
rlabel metal1 19090 8058 19090 8058 0 _0483_
rlabel via2 11546 8772 11546 8772 0 _0484_
rlabel metal1 18124 13294 18124 13294 0 _0485_
rlabel metal1 7314 7446 7314 7446 0 _0486_
rlabel metal1 17526 7922 17526 7922 0 _0487_
rlabel metal1 15318 5338 15318 5338 0 _0488_
rlabel metal2 18722 6596 18722 6596 0 _0489_
rlabel metal1 18492 8058 18492 8058 0 _0490_
rlabel metal2 17204 4114 17204 4114 0 _0491_
rlabel metal1 17710 8806 17710 8806 0 _0492_
rlabel metal2 14950 3876 14950 3876 0 _0493_
rlabel metal1 17250 8500 17250 8500 0 _0494_
rlabel metal1 17572 6630 17572 6630 0 _0495_
rlabel metal1 17802 8942 17802 8942 0 _0496_
rlabel metal1 12650 6392 12650 6392 0 _0497_
rlabel metal1 14582 4182 14582 4182 0 _0498_
rlabel metal1 13708 8942 13708 8942 0 _0499_
rlabel metal1 17986 8976 17986 8976 0 _0500_
rlabel metal1 19757 8398 19757 8398 0 _0501_
rlabel metal2 14582 10013 14582 10013 0 _0502_
rlabel metal2 17066 5916 17066 5916 0 _0503_
rlabel metal1 19182 8398 19182 8398 0 _0504_
rlabel metal2 15778 6443 15778 6443 0 _0505_
rlabel metal1 10948 6766 10948 6766 0 _0506_
rlabel metal2 17618 3825 17618 3825 0 _0507_
rlabel metal1 14122 4148 14122 4148 0 _0508_
rlabel metal1 20286 8602 20286 8602 0 _0509_
rlabel metal1 31326 5236 31326 5236 0 _0510_
rlabel metal3 31349 12852 31349 12852 0 _0511_
rlabel metal2 31050 13668 31050 13668 0 _0512_
rlabel metal1 30038 13328 30038 13328 0 _0513_
rlabel metal1 29624 12818 29624 12818 0 _0514_
rlabel metal1 30912 12614 30912 12614 0 _0515_
rlabel metal1 32108 10642 32108 10642 0 _0516_
rlabel metal2 29486 10880 29486 10880 0 _0517_
rlabel metal1 29900 12410 29900 12410 0 _0518_
rlabel metal1 31050 12852 31050 12852 0 _0519_
rlabel metal1 30774 12954 30774 12954 0 _0520_
rlabel metal1 30682 13158 30682 13158 0 _0521_
rlabel metal2 31970 10812 31970 10812 0 _0522_
rlabel viali 31786 7859 31786 7859 0 _0523_
rlabel metal2 28934 6528 28934 6528 0 _0524_
rlabel metal2 31326 11356 31326 11356 0 _0525_
rlabel metal1 32338 10676 32338 10676 0 _0526_
rlabel metal1 28704 10642 28704 10642 0 _0527_
rlabel metal1 28750 9520 28750 9520 0 _0528_
rlabel metal1 28428 6766 28428 6766 0 _0529_
rlabel metal2 30682 9350 30682 9350 0 _0530_
rlabel metal1 27968 8398 27968 8398 0 _0531_
rlabel metal1 27876 6834 27876 6834 0 _0532_
rlabel metal1 18998 12852 18998 12852 0 _0533_
rlabel metal1 28612 10574 28612 10574 0 _0534_
rlabel metal1 30360 10030 30360 10030 0 _0535_
rlabel metal1 29716 10234 29716 10234 0 _0536_
rlabel metal1 29394 7242 29394 7242 0 _0537_
rlabel metal1 30452 8466 30452 8466 0 _0538_
rlabel metal2 27922 10030 27922 10030 0 _0539_
rlabel metal1 27554 7378 27554 7378 0 _0540_
rlabel metal1 27508 7310 27508 7310 0 _0541_
rlabel metal1 25346 8874 25346 8874 0 _0542_
rlabel metal1 29210 9520 29210 9520 0 _0543_
rlabel metal1 28566 8058 28566 8058 0 _0544_
rlabel metal2 26910 8704 26910 8704 0 _0545_
rlabel metal1 28842 8500 28842 8500 0 _0546_
rlabel metal1 27784 10642 27784 10642 0 _0547_
rlabel metal1 27186 10778 27186 10778 0 _0548_
rlabel metal1 28980 10166 28980 10166 0 _0549_
rlabel metal2 28474 9690 28474 9690 0 _0550_
rlabel metal2 27002 9452 27002 9452 0 _0551_
rlabel metal1 24886 9044 24886 9044 0 _0552_
rlabel metal1 24794 7378 24794 7378 0 _0553_
rlabel metal1 25346 12750 25346 12750 0 _0554_
rlabel metal2 21758 9146 21758 9146 0 _0555_
rlabel metal1 26036 12614 26036 12614 0 _0556_
rlabel metal1 30176 10642 30176 10642 0 _0557_
rlabel metal1 30452 9894 30452 9894 0 _0558_
rlabel metal1 27784 6766 27784 6766 0 _0559_
rlabel metal1 30774 7208 30774 7208 0 _0560_
rlabel metal1 31418 6834 31418 6834 0 _0561_
rlabel metal1 31004 7378 31004 7378 0 _0562_
rlabel via1 26713 6834 26713 6834 0 _0563_
rlabel metal1 24932 8466 24932 8466 0 _0564_
rlabel metal1 28566 8534 28566 8534 0 _0565_
rlabel metal1 31050 8500 31050 8500 0 _0566_
rlabel metal1 28842 8262 28842 8262 0 _0567_
rlabel metal1 26450 7412 26450 7412 0 _0568_
rlabel viali 26713 7378 26713 7378 0 _0569_
rlabel metal1 25714 7446 25714 7446 0 _0570_
rlabel metal2 22034 8772 22034 8772 0 _0571_
rlabel metal2 20746 13702 20746 13702 0 _0572_
rlabel metal1 21068 9010 21068 9010 0 _0573_
rlabel metal1 19228 18190 19228 18190 0 _0574_
rlabel metal1 18722 18258 18722 18258 0 _0575_
rlabel metal1 18814 4556 18814 4556 0 _0576_
rlabel metal1 15778 10064 15778 10064 0 _0577_
rlabel metal1 18446 5882 18446 5882 0 _0578_
rlabel metal3 15295 12580 15295 12580 0 _0579_
rlabel metal1 15778 3570 15778 3570 0 _0580_
rlabel metal1 12052 8398 12052 8398 0 _0581_
rlabel metal1 17250 4080 17250 4080 0 _0582_
rlabel metal1 17342 6426 17342 6426 0 _0583_
rlabel metal1 18354 6324 18354 6324 0 _0584_
rlabel metal1 17066 11662 17066 11662 0 _0585_
rlabel metal2 19366 6800 19366 6800 0 _0586_
rlabel metal1 17940 6290 17940 6290 0 _0587_
rlabel metal1 12834 5644 12834 5644 0 _0588_
rlabel metal1 18078 10676 18078 10676 0 _0589_
rlabel metal1 19102 6222 19102 6222 0 _0590_
rlabel metal1 10028 10030 10028 10030 0 _0591_
rlabel metal2 16054 3230 16054 3230 0 _0592_
rlabel metal1 18124 6766 18124 6766 0 _0593_
rlabel metal2 19274 6562 19274 6562 0 _0594_
rlabel metal1 21068 6426 21068 6426 0 _0595_
rlabel metal1 29578 7514 29578 7514 0 _0596_
rlabel metal1 26174 8364 26174 8364 0 _0597_
rlabel metal1 25254 7854 25254 7854 0 _0598_
rlabel metal1 24334 7310 24334 7310 0 _0599_
rlabel metal1 23184 8942 23184 8942 0 _0600_
rlabel metal1 21666 7820 21666 7820 0 _0601_
rlabel metal1 24702 6766 24702 6766 0 _0602_
rlabel metal1 15778 14416 15778 14416 0 _0603_
rlabel metal1 21804 7854 21804 7854 0 _0604_
rlabel metal2 21574 15028 21574 15028 0 _0605_
rlabel metal1 13524 17510 13524 17510 0 _0606_
rlabel metal1 20976 17646 20976 17646 0 _0607_
rlabel metal1 26910 8942 26910 8942 0 _0608_
rlabel metal1 24748 9690 24748 9690 0 _0609_
rlabel via1 23966 9690 23966 9690 0 _0610_
rlabel metal1 23874 8602 23874 8602 0 _0611_
rlabel metal1 22586 9690 22586 9690 0 _0612_
rlabel metal1 19550 7990 19550 7990 0 _0613_
rlabel metal1 19228 7514 19228 7514 0 _0614_
rlabel metal1 11516 7854 11516 7854 0 _0615_
rlabel metal1 12972 3978 12972 3978 0 _0616_
rlabel metal1 19458 8976 19458 8976 0 _0617_
rlabel metal1 19964 9146 19964 9146 0 _0618_
rlabel metal1 19274 4658 19274 4658 0 _0619_
rlabel metal1 18262 3978 18262 3978 0 _0620_
rlabel metal2 18262 4539 18262 4539 0 _0621_
rlabel metal1 18814 3978 18814 3978 0 _0622_
rlabel metal1 19228 4794 19228 4794 0 _0623_
rlabel metal1 19412 10166 19412 10166 0 _0624_
rlabel metal1 17802 16150 17802 16150 0 _0625_
rlabel metal1 17020 16082 17020 16082 0 _0626_
rlabel metal2 32890 10030 32890 10030 0 _0627_
rlabel metal2 27370 10030 27370 10030 0 _0628_
rlabel metal1 25346 9350 25346 9350 0 _0629_
rlabel metal1 23552 7786 23552 7786 0 _0630_
rlabel metal2 25070 7208 25070 7208 0 _0631_
rlabel metal1 23368 7514 23368 7514 0 _0632_
rlabel metal2 22310 8194 22310 8194 0 _0633_
rlabel metal1 15870 3910 15870 3910 0 _0634_
rlabel metal1 16744 3162 16744 3162 0 _0635_
rlabel metal1 15824 3502 15824 3502 0 _0636_
rlabel metal1 16330 3434 16330 3434 0 _0637_
rlabel metal1 16376 3638 16376 3638 0 _0638_
rlabel metal2 20102 9554 20102 9554 0 _0639_
rlabel metal1 18193 3570 18193 3570 0 _0640_
rlabel metal2 17342 3740 17342 3740 0 _0641_
rlabel metal1 18446 3366 18446 3366 0 _0642_
rlabel metal2 21390 7956 21390 7956 0 _0643_
rlabel metal2 21390 11764 21390 11764 0 _0644_
rlabel metal1 20838 14994 20838 14994 0 _0645_
rlabel metal2 19458 10880 19458 10880 0 _0646_
rlabel metal1 14444 8942 14444 8942 0 _0647_
rlabel metal2 17526 4811 17526 4811 0 _0648_
rlabel metal1 19596 10438 19596 10438 0 _0649_
rlabel metal1 19826 12818 19826 12818 0 _0650_
rlabel metal1 19918 10574 19918 10574 0 _0651_
rlabel metal1 20286 10506 20286 10506 0 _0652_
rlabel metal2 13570 3706 13570 3706 0 _0653_
rlabel metal1 13984 9146 13984 9146 0 _0654_
rlabel metal1 14260 9622 14260 9622 0 _0655_
rlabel metal1 13777 5610 13777 5610 0 _0656_
rlabel metal1 14306 6970 14306 6970 0 _0657_
rlabel metal1 15502 13974 15502 13974 0 _0658_
rlabel metal2 20562 10030 20562 10030 0 _0659_
rlabel metal1 28382 10676 28382 10676 0 _0660_
rlabel metal1 28382 10234 28382 10234 0 _0661_
rlabel metal1 27002 10710 27002 10710 0 _0662_
rlabel metal1 24794 10540 24794 10540 0 _0663_
rlabel metal1 23690 11118 23690 11118 0 _0664_
rlabel metal1 20838 10676 20838 10676 0 _0665_
rlabel metal1 21850 9656 21850 9656 0 _0666_
rlabel metal1 19964 15334 19964 15334 0 _0667_
rlabel metal1 18722 15436 18722 15436 0 _0668_
rlabel metal1 16146 5882 16146 5882 0 _0669_
rlabel metal1 15870 6324 15870 6324 0 _0670_
rlabel metal1 16514 6426 16514 6426 0 _0671_
rlabel metal1 16422 3978 16422 3978 0 _0672_
rlabel metal1 16652 9078 16652 9078 0 _0673_
rlabel metal1 16376 8806 16376 8806 0 _0674_
rlabel metal1 17020 9146 17020 9146 0 _0675_
rlabel metal1 15042 12784 15042 12784 0 _0676_
rlabel metal1 16238 10132 16238 10132 0 _0677_
rlabel metal1 16790 9554 16790 9554 0 _0678_
rlabel viali 16054 9482 16054 9482 0 _0679_
rlabel metal1 22172 10030 22172 10030 0 _0680_
rlabel metal1 22586 9146 22586 9146 0 _0681_
rlabel metal1 25990 10778 25990 10778 0 _0682_
rlabel metal1 22770 10676 22770 10676 0 _0683_
rlabel metal1 22770 10030 22770 10030 0 _0684_
rlabel metal1 21988 10234 21988 10234 0 _0685_
rlabel metal1 22310 14858 22310 14858 0 _0686_
rlabel metal1 30590 10574 30590 10574 0 _0687_
rlabel metal1 29716 10778 29716 10778 0 _0688_
rlabel metal1 27462 11594 27462 11594 0 _0689_
rlabel metal1 25944 11594 25944 11594 0 _0690_
rlabel metal1 24840 11322 24840 11322 0 _0691_
rlabel metal2 24702 13634 24702 13634 0 _0692_
rlabel metal1 24380 10778 24380 10778 0 _0693_
rlabel metal1 25254 13498 25254 13498 0 _0694_
rlabel metal1 12558 3672 12558 3672 0 _0695_
rlabel metal1 16744 13226 16744 13226 0 _0696_
rlabel metal1 15824 12410 15824 12410 0 _0697_
rlabel metal2 16974 13158 16974 13158 0 _0698_
rlabel metal1 7544 12818 7544 12818 0 _0699_
rlabel metal2 16790 13294 16790 13294 0 _0700_
rlabel metal2 17158 13736 17158 13736 0 _0701_
rlabel metal1 18768 10642 18768 10642 0 _0702_
rlabel metal1 18492 10778 18492 10778 0 _0703_
rlabel metal1 18492 11322 18492 11322 0 _0704_
rlabel metal1 18492 11866 18492 11866 0 _0705_
rlabel metal2 18814 14144 18814 14144 0 _0706_
rlabel metal1 13800 4794 13800 4794 0 _0707_
rlabel metal1 12972 3706 12972 3706 0 _0708_
rlabel metal2 12742 3298 12742 3298 0 _0709_
rlabel metal2 12374 3808 12374 3808 0 _0710_
rlabel metal1 14812 3094 14812 3094 0 _0711_
rlabel metal1 14352 2958 14352 2958 0 _0712_
rlabel metal1 13202 4046 13202 4046 0 _0713_
rlabel metal1 14444 14382 14444 14382 0 _0714_
rlabel metal1 28198 12172 28198 12172 0 _0715_
rlabel metal1 27968 12274 27968 12274 0 _0716_
rlabel metal1 26128 12886 26128 12886 0 _0717_
rlabel metal2 22034 12903 22034 12903 0 _0718_
rlabel metal1 22126 13974 22126 13974 0 _0719_
rlabel metal1 20427 14042 20427 14042 0 _0720_
rlabel metal1 14398 14586 14398 14586 0 _0721_
rlabel metal1 14030 15470 14030 15470 0 _0722_
rlabel metal1 13800 9078 13800 9078 0 _0723_
rlabel metal1 14352 9350 14352 9350 0 _0724_
rlabel metal1 15456 10778 15456 10778 0 _0725_
rlabel metal1 14812 11322 14812 11322 0 _0726_
rlabel metal2 14582 12823 14582 12823 0 _0727_
rlabel metal1 14398 11084 14398 11084 0 _0728_
rlabel metal2 14582 11492 14582 11492 0 _0729_
rlabel metal1 12926 11764 12926 11764 0 _0730_
rlabel metal1 14007 7446 14007 7446 0 _0731_
rlabel metal1 14122 11662 14122 11662 0 _0732_
rlabel metal2 22034 11322 22034 11322 0 _0733_
rlabel metal1 21850 11152 21850 11152 0 _0734_
rlabel metal2 27416 12614 27416 12614 0 _0735_
rlabel metal1 25806 12070 25806 12070 0 _0736_
rlabel metal1 23322 12342 23322 12342 0 _0737_
rlabel metal1 21712 11118 21712 11118 0 _0738_
rlabel metal2 22264 13124 22264 13124 0 _0739_
rlabel metal1 21712 16558 21712 16558 0 _0740_
rlabel metal1 11730 12716 11730 12716 0 _0741_
rlabel metal1 10994 7378 10994 7378 0 _0742_
rlabel metal1 10718 11594 10718 11594 0 _0743_
rlabel metal1 10350 12648 10350 12648 0 _0744_
rlabel metal1 11269 11798 11269 11798 0 _0745_
rlabel metal1 10550 12886 10550 12886 0 _0746_
rlabel metal1 10994 12954 10994 12954 0 _0747_
rlabel metal1 12052 9146 12052 9146 0 _0748_
rlabel metal1 10718 10132 10718 10132 0 _0749_
rlabel metal1 12236 10778 12236 10778 0 _0750_
rlabel metal1 12144 11186 12144 11186 0 _0751_
rlabel metal2 12098 11492 12098 11492 0 _0752_
rlabel metal1 11822 13294 11822 13294 0 _0753_
rlabel metal1 25438 6086 25438 6086 0 _0754_
rlabel metal1 27324 12614 27324 12614 0 _0755_
rlabel metal1 22586 13294 22586 13294 0 _0756_
rlabel metal2 22034 13209 22034 13209 0 _0757_
rlabel metal1 11822 13498 11822 13498 0 _0758_
rlabel metal1 11224 17170 11224 17170 0 _0759_
rlabel metal1 24150 12954 24150 12954 0 _0760_
rlabel metal1 23414 13906 23414 13906 0 _0761_
rlabel metal1 17066 14552 17066 14552 0 _0762_
rlabel metal1 10258 7378 10258 7378 0 _0763_
rlabel metal1 10994 7480 10994 7480 0 _0764_
rlabel metal1 12006 7854 12006 7854 0 _0765_
rlabel metal1 12374 7922 12374 7922 0 _0766_
rlabel metal1 11914 7514 11914 7514 0 _0767_
rlabel metal1 13110 5610 13110 5610 0 _0768_
rlabel metal2 12926 6596 12926 6596 0 _0769_
rlabel metal1 12604 7514 12604 7514 0 _0770_
rlabel metal2 12558 14110 12558 14110 0 _0771_
rlabel metal2 12742 15300 12742 15300 0 _0772_
rlabel metal1 12190 16082 12190 16082 0 _0773_
rlabel metal2 11178 8500 11178 8500 0 _0774_
rlabel metal1 11224 8942 11224 8942 0 _0775_
rlabel metal2 11270 9316 11270 9316 0 _0776_
rlabel metal1 10350 9996 10350 9996 0 _0777_
rlabel via1 10337 9554 10337 9554 0 _0778_
rlabel metal2 10442 9316 10442 9316 0 _0779_
rlabel metal1 11638 13702 11638 13702 0 _0780_
rlabel metal1 26910 12750 26910 12750 0 _0781_
rlabel metal1 23368 13294 23368 13294 0 _0782_
rlabel metal1 22264 12818 22264 12818 0 _0783_
rlabel metal1 20516 12682 20516 12682 0 _0784_
rlabel metal2 12466 14688 12466 14688 0 _0785_
rlabel metal1 11592 14994 11592 14994 0 _0786_
rlabel metal1 12880 10778 12880 10778 0 _0787_
rlabel metal2 13294 12857 13294 12857 0 _0788_
rlabel metal1 17526 13396 17526 13396 0 _0789_
rlabel metal1 13846 13294 13846 13294 0 _0790_
rlabel metal1 13708 13498 13708 13498 0 _0791_
rlabel metal1 16882 13770 16882 13770 0 _0792_
rlabel metal1 14904 12410 14904 12410 0 _0793_
rlabel metal1 14352 13498 14352 13498 0 _0794_
rlabel metal1 22264 10778 22264 10778 0 _0795_
rlabel metal3 16031 13804 16031 13804 0 _0796_
rlabel metal1 14536 14042 14536 14042 0 _0797_
rlabel metal1 14904 19890 14904 19890 0 _0798_
rlabel metal1 13938 19958 13938 19958 0 _0799_
rlabel metal1 20286 13158 20286 13158 0 _0800_
rlabel metal1 16422 14042 16422 14042 0 _0801_
rlabel metal2 12926 13362 12926 13362 0 _0802_
rlabel metal1 15824 12750 15824 12750 0 _0803_
rlabel metal1 15548 12954 15548 12954 0 _0804_
rlabel metal1 15728 14042 15728 14042 0 _0805_
rlabel metal1 16376 14450 16376 14450 0 _0806_
rlabel metal1 16284 14586 16284 14586 0 _0807_
rlabel metal1 15548 18734 15548 18734 0 _0808_
rlabel metal1 17112 12886 17112 12886 0 _0809_
rlabel metal1 17342 12274 17342 12274 0 _0810_
rlabel metal2 17158 12410 17158 12410 0 _0811_
rlabel metal1 17388 12410 17388 12410 0 _0812_
rlabel metal2 17434 13005 17434 13005 0 _0813_
rlabel metal2 22310 13668 22310 13668 0 _0814_
rlabel metal2 22770 17782 22770 17782 0 _0815_
rlabel metal1 21988 21658 21988 21658 0 _0816_
rlabel metal1 18998 12410 18998 12410 0 _0817_
rlabel metal2 17342 12240 17342 12240 0 _0818_
rlabel metal1 18262 12682 18262 12682 0 _0819_
rlabel metal1 20102 12886 20102 12886 0 _0820_
rlabel metal1 23552 13498 23552 13498 0 _0821_
rlabel metal1 23230 20570 23230 20570 0 _0822_
rlabel metal1 19780 12410 19780 12410 0 _0823_
rlabel metal1 19136 12750 19136 12750 0 _0824_
rlabel metal1 20470 12954 20470 12954 0 _0825_
rlabel metal1 23736 13294 23736 13294 0 _0826_
rlabel metal1 23644 13226 23644 13226 0 _0827_
rlabel metal1 23276 22610 23276 22610 0 _0828_
rlabel metal1 16790 36788 16790 36788 0 _0829_
rlabel metal1 21574 15130 21574 15130 0 _0830_
rlabel metal1 18630 14042 18630 14042 0 _0831_
rlabel metal1 21114 14994 21114 14994 0 _0832_
rlabel metal1 21574 14450 21574 14450 0 _0833_
rlabel metal1 14444 23086 14444 23086 0 _0834_
rlabel metal1 21114 23290 21114 23290 0 _0835_
rlabel metal1 16376 21114 16376 21114 0 _0836_
rlabel metal1 20700 20910 20700 20910 0 _0837_
rlabel metal1 18906 20026 18906 20026 0 _0838_
rlabel metal2 20010 23188 20010 23188 0 _0839_
rlabel metal2 17618 22304 17618 22304 0 _0840_
rlabel metal1 18814 23698 18814 23698 0 _0841_
rlabel metal1 12788 21522 12788 21522 0 _0842_
rlabel metal2 19826 22423 19826 22423 0 _0843_
rlabel metal1 10902 23086 10902 23086 0 _0844_
rlabel metal1 12328 23698 12328 23698 0 _0845_
rlabel metal1 11040 22746 11040 22746 0 _0846_
rlabel metal1 11132 24786 11132 24786 0 _0847_
rlabel metal1 14674 24208 14674 24208 0 _0848_
rlabel metal1 16928 24174 16928 24174 0 _0849_
rlabel metal1 17250 33388 17250 33388 0 _0850_
rlabel metal1 22586 30702 22586 30702 0 _0851_
rlabel metal1 24242 29614 24242 29614 0 _0852_
rlabel metal1 22126 30736 22126 30736 0 _0853_
rlabel metal1 12328 26350 12328 26350 0 _0854_
rlabel metal2 14122 25738 14122 25738 0 _0855_
rlabel metal1 14490 27608 14490 27608 0 _0856_
rlabel metal1 16560 31994 16560 31994 0 _0857_
rlabel metal1 11454 28050 11454 28050 0 _0858_
rlabel metal1 14904 33626 14904 33626 0 _0859_
rlabel metal1 16376 33490 16376 33490 0 _0860_
rlabel metal1 15180 37298 15180 37298 0 _0861_
rlabel metal1 15364 36754 15364 36754 0 _0862_
rlabel metal1 7498 37230 7498 37230 0 _0863_
rlabel metal1 7498 38930 7498 38930 0 _0864_
rlabel metal1 8142 39406 8142 39406 0 _0865_
rlabel metal1 11362 41106 11362 41106 0 _0866_
rlabel metal2 10166 42228 10166 42228 0 _0867_
rlabel metal1 8004 41582 8004 41582 0 _0868_
rlabel metal1 16192 41106 16192 41106 0 _0869_
rlabel metal1 17526 39610 17526 39610 0 _0870_
rlabel metal1 13754 39508 13754 39508 0 _0871_
rlabel metal1 15548 35598 15548 35598 0 _0872_
rlabel metal1 14674 35598 14674 35598 0 _0873_
rlabel metal1 21390 26350 21390 26350 0 _0874_
rlabel metal1 16882 27472 16882 27472 0 _0875_
rlabel metal1 22172 26962 22172 26962 0 _0876_
rlabel metal1 24058 33524 24058 33524 0 _0877_
rlabel metal1 18308 29138 18308 29138 0 _0878_
rlabel metal1 21482 36176 21482 36176 0 _0879_
rlabel metal2 18906 34884 18906 34884 0 _0880_
rlabel metal1 21390 36686 21390 36686 0 _0881_
rlabel metal1 12926 35666 12926 35666 0 _0882_
rlabel metal1 10626 36142 10626 36142 0 _0883_
rlabel metal1 10396 38930 10396 38930 0 _0884_
rlabel metal1 11270 44370 11270 44370 0 _0885_
rlabel metal2 14122 44404 14122 44404 0 _0886_
rlabel metal1 16284 44506 16284 44506 0 _0887_
rlabel metal1 19734 43146 19734 43146 0 _0888_
rlabel metal1 19228 39066 19228 39066 0 _0889_
rlabel metal1 21298 40052 21298 40052 0 _0890_
rlabel metal1 21620 37842 21620 37842 0 _0891_
rlabel metal1 8050 10574 8050 10574 0 _0892_
rlabel metal2 7498 10948 7498 10948 0 _0893_
rlabel metal1 7544 7514 7544 7514 0 _0894_
rlabel metal1 7360 9010 7360 9010 0 _0895_
rlabel metal1 6762 5712 6762 5712 0 _0896_
rlabel metal1 7268 6766 7268 6766 0 _0897_
rlabel metal1 6900 6766 6900 6766 0 _0898_
rlabel metal2 8234 7004 8234 7004 0 _0899_
rlabel metal1 7452 4590 7452 4590 0 _0900_
rlabel metal1 7268 8942 7268 8942 0 _0901_
rlabel metal1 8004 8942 8004 8942 0 _0902_
rlabel metal1 7774 11186 7774 11186 0 _0903_
rlabel metal1 7958 12750 7958 12750 0 _0904_
rlabel metal1 8648 13294 8648 13294 0 _0905_
rlabel metal1 37904 8942 37904 8942 0 _0906_
rlabel metal1 35466 8432 35466 8432 0 _0907_
rlabel metal1 34776 13906 34776 13906 0 _0908_
rlabel metal1 35512 12818 35512 12818 0 _0909_
rlabel metal1 36478 34374 36478 34374 0 _0910_
rlabel metal1 27370 37808 27370 37808 0 _0911_
rlabel metal1 28244 35598 28244 35598 0 _0912_
rlabel metal2 36570 34782 36570 34782 0 _0913_
rlabel metal1 25806 36142 25806 36142 0 _0914_
rlabel metal1 34776 32402 34776 32402 0 _0915_
rlabel metal1 35236 21998 35236 21998 0 _0916_
rlabel metal1 25254 2414 25254 2414 0 _0917_
rlabel metal1 36708 44370 36708 44370 0 _0918_
rlabel metal1 8050 2992 8050 2992 0 _0919_
rlabel metal2 36570 3332 36570 3332 0 _0920_
rlabel metal1 19228 3162 19228 3162 0 _0921_
rlabel metal1 19550 44880 19550 44880 0 _0922_
rlabel metal1 36708 24786 36708 24786 0 _0923_
rlabel metal1 6256 44370 6256 44370 0 _0924_
rlabel metal1 31970 44370 31970 44370 0 _0925_
rlabel metal1 26404 2618 26404 2618 0 _0926_
rlabel metal1 6164 25874 6164 25874 0 _0927_
rlabel metal1 24932 42670 24932 42670 0 _0928_
rlabel metal1 2392 9146 2392 9146 0 _0929_
rlabel metal1 2438 18258 2438 18258 0 _0930_
rlabel metal1 2599 6834 2599 6834 0 _0931_
rlabel metal2 43378 7684 43378 7684 0 _0932_
rlabel metal1 2484 35666 2484 35666 0 _0933_
rlabel metal1 43700 32402 43700 32402 0 _0934_
rlabel metal2 43286 14790 43286 14790 0 _0935_
rlabel metal1 35558 40528 35558 40528 0 _0936_
rlabel metal1 35420 40698 35420 40698 0 _0937_
rlabel metal1 35420 39406 35420 39406 0 _0938_
rlabel metal1 34868 39406 34868 39406 0 _0939_
rlabel metal1 35742 36822 35742 36822 0 _0940_
rlabel metal1 35972 37638 35972 37638 0 _0941_
rlabel metal1 37996 37978 37996 37978 0 _0942_
rlabel metal1 37582 38318 37582 38318 0 _0943_
rlabel metal1 40112 37230 40112 37230 0 _0944_
rlabel metal1 41676 40018 41676 40018 0 _0945_
rlabel metal1 41032 40018 41032 40018 0 _0946_
rlabel metal2 41262 38454 41262 38454 0 _0947_
rlabel metal1 41262 37162 41262 37162 0 _0948_
rlabel metal2 41446 36720 41446 36720 0 _0949_
rlabel metal1 40710 36856 40710 36856 0 _0950_
rlabel metal1 38180 36618 38180 36618 0 _0951_
rlabel metal1 38456 37230 38456 37230 0 _0952_
rlabel metal1 37766 36788 37766 36788 0 _0953_
rlabel metal1 38042 39372 38042 39372 0 _0954_
rlabel metal1 41906 41548 41906 41548 0 _0955_
rlabel metal1 38824 37978 38824 37978 0 _0956_
rlabel metal1 40250 37774 40250 37774 0 _0957_
rlabel metal1 40388 38726 40388 38726 0 _0958_
rlabel metal1 39468 41174 39468 41174 0 _0959_
rlabel metal1 39422 39440 39422 39440 0 _0960_
rlabel metal2 38870 42534 38870 42534 0 _0961_
rlabel metal1 39238 41242 39238 41242 0 _0962_
rlabel metal1 38686 40494 38686 40494 0 _0963_
rlabel metal1 40710 41106 40710 41106 0 _0964_
rlabel metal1 40756 40970 40756 40970 0 _0965_
rlabel metal1 40664 41242 40664 41242 0 _0966_
rlabel metal1 41952 41786 41952 41786 0 _0967_
rlabel via1 42098 41446 42098 41446 0 _0968_
rlabel metal2 42274 41990 42274 41990 0 _0969_
rlabel metal1 43654 40052 43654 40052 0 _0970_
rlabel metal1 44022 40460 44022 40460 0 _0971_
rlabel metal1 39422 35020 39422 35020 0 _0972_
rlabel metal1 42366 39474 42366 39474 0 _0973_
rlabel metal1 39836 35258 39836 35258 0 _0974_
rlabel metal1 39744 36142 39744 36142 0 _0975_
rlabel metal1 40342 33014 40342 33014 0 _0976_
rlabel metal2 40618 33354 40618 33354 0 _0977_
rlabel metal1 42826 35054 42826 35054 0 _0978_
rlabel metal1 43516 35054 43516 35054 0 _0979_
rlabel metal1 42090 36890 42090 36890 0 _0980_
rlabel metal1 42474 37162 42474 37162 0 _0981_
rlabel metal1 41630 36788 41630 36788 0 _0982_
rlabel metal1 34454 8466 34454 8466 0 _0983_
rlabel metal1 42090 17204 42090 17204 0 _0984_
rlabel metal2 43378 18598 43378 18598 0 _0985_
rlabel metal1 39744 17170 39744 17170 0 _0986_
rlabel metal1 42044 15470 42044 15470 0 _0987_
rlabel metal1 39330 17204 39330 17204 0 _0988_
rlabel metal1 39471 17306 39471 17306 0 _0989_
rlabel metal1 38778 18802 38778 18802 0 _0990_
rlabel metal1 37996 18734 37996 18734 0 _0991_
rlabel metal1 36846 18292 36846 18292 0 _0992_
rlabel metal1 35880 14042 35880 14042 0 _0993_
rlabel metal1 18400 19754 18400 19754 0 _0994_
rlabel metal1 25070 37842 25070 37842 0 _0995_
rlabel metal1 32798 33422 32798 33422 0 _0996_
rlabel metal1 37950 8364 37950 8364 0 _0997_
rlabel metal1 35650 8500 35650 8500 0 _0998_
rlabel metal1 35926 10438 35926 10438 0 _0999_
rlabel metal1 34868 12818 34868 12818 0 _1000_
rlabel metal1 36846 15334 36846 15334 0 _1001_
rlabel metal1 35144 14586 35144 14586 0 _1002_
rlabel metal2 21206 29716 21206 29716 0 _1003_
rlabel metal1 13616 31246 13616 31246 0 _1004_
rlabel metal1 13156 29614 13156 29614 0 _1005_
rlabel metal2 12558 33405 12558 33405 0 _1006_
rlabel metal1 21160 32742 21160 32742 0 _1007_
rlabel metal1 11638 31858 11638 31858 0 _1008_
rlabel metal1 12604 29818 12604 29818 0 _1009_
rlabel metal1 11684 29750 11684 29750 0 _1010_
rlabel metal1 11178 30022 11178 30022 0 _1011_
rlabel metal2 11546 29172 11546 29172 0 _1012_
rlabel metal1 12581 29682 12581 29682 0 _1013_
rlabel metal1 12834 30260 12834 30260 0 _1014_
rlabel metal2 12650 29852 12650 29852 0 _1015_
rlabel metal1 13708 29478 13708 29478 0 _1016_
rlabel metal1 15180 31858 15180 31858 0 _1017_
rlabel metal1 15226 31348 15226 31348 0 _1018_
rlabel metal1 18722 30260 18722 30260 0 _1019_
rlabel metal1 15732 31110 15732 31110 0 _1020_
rlabel metal1 14628 31654 14628 31654 0 _1021_
rlabel metal1 18262 32946 18262 32946 0 _1022_
rlabel metal1 9338 35088 9338 35088 0 _1023_
rlabel metal1 14858 28730 14858 28730 0 _1024_
rlabel via1 14296 30906 14296 30906 0 _1025_
rlabel metal1 12052 30362 12052 30362 0 _1026_
rlabel metal1 9154 31858 9154 31858 0 _1027_
rlabel metal1 11270 30702 11270 30702 0 _1028_
rlabel metal1 12282 30634 12282 30634 0 _1029_
rlabel metal1 19044 24786 19044 24786 0 _1030_
rlabel metal1 14582 30702 14582 30702 0 _1031_
rlabel metal1 13340 30906 13340 30906 0 _1032_
rlabel metal2 13110 25874 13110 25874 0 _1033_
rlabel metal2 12098 28254 12098 28254 0 _1034_
rlabel metal1 13018 27642 13018 27642 0 _1035_
rlabel metal2 12466 29410 12466 29410 0 _1036_
rlabel metal1 19918 31314 19918 31314 0 _1037_
rlabel metal2 13570 30770 13570 30770 0 _1038_
rlabel metal1 12880 30634 12880 30634 0 _1039_
rlabel via2 14122 30651 14122 30651 0 _1040_
rlabel metal1 6256 32810 6256 32810 0 _1041_
rlabel metal2 8970 34901 8970 34901 0 _1042_
rlabel metal1 10074 25704 10074 25704 0 _1043_
rlabel metal1 9944 26010 9944 26010 0 _1044_
rlabel metal1 10994 25908 10994 25908 0 _1045_
rlabel metal1 8924 27846 8924 27846 0 _1046_
rlabel metal1 9614 28458 9614 28458 0 _1047_
rlabel metal1 8464 28050 8464 28050 0 _1048_
rlabel metal1 8326 28594 8326 28594 0 _1049_
rlabel metal1 8786 28730 8786 28730 0 _1050_
rlabel metal1 9354 28458 9354 28458 0 _1051_
rlabel metal1 9292 28730 9292 28730 0 _1052_
rlabel metal2 6118 28220 6118 28220 0 _1053_
rlabel via1 5848 28050 5848 28050 0 _1054_
rlabel metal1 6946 28628 6946 28628 0 _1055_
rlabel metal1 5382 28118 5382 28118 0 _1056_
rlabel metal1 5796 28934 5796 28934 0 _1057_
rlabel metal1 5612 29818 5612 29818 0 _1058_
rlabel metal1 5558 29274 5558 29274 0 _1059_
rlabel metal1 4784 29138 4784 29138 0 _1060_
rlabel metal2 6118 30532 6118 30532 0 _1061_
rlabel metal2 5658 30532 5658 30532 0 _1062_
rlabel metal1 6762 30906 6762 30906 0 _1063_
rlabel metal1 7590 30770 7590 30770 0 _1064_
rlabel metal2 7406 30872 7406 30872 0 _1065_
rlabel metal2 6210 32071 6210 32071 0 _1066_
rlabel metal1 7774 29648 7774 29648 0 _1067_
rlabel metal1 8326 31246 8326 31246 0 _1068_
rlabel metal1 8004 31994 8004 31994 0 _1069_
rlabel metal2 8556 31790 8556 31790 0 _1070_
rlabel metal2 8050 32164 8050 32164 0 _1071_
rlabel metal1 8970 31348 8970 31348 0 _1072_
rlabel metal1 7314 33490 7314 33490 0 _1073_
rlabel metal1 5658 33082 5658 33082 0 _1074_
rlabel metal2 6394 34102 6394 34102 0 _1075_
rlabel metal1 5512 32810 5512 32810 0 _1076_
rlabel metal1 5060 32878 5060 32878 0 _1077_
rlabel metal2 5658 35088 5658 35088 0 _1078_
rlabel metal1 5382 35156 5382 35156 0 _1079_
rlabel metal1 5980 35802 5980 35802 0 _1080_
rlabel metal1 6854 34612 6854 34612 0 _1081_
rlabel metal1 5888 34170 5888 34170 0 _1082_
rlabel metal1 8004 35054 8004 35054 0 _1083_
rlabel metal1 8004 35258 8004 35258 0 _1084_
rlabel metal1 9016 34918 9016 34918 0 _1085_
rlabel metal2 7682 35462 7682 35462 0 _1086_
rlabel metal2 8326 34918 8326 34918 0 _1087_
rlabel metal1 8740 34442 8740 34442 0 _1088_
rlabel metal1 9154 33966 9154 33966 0 _1089_
rlabel metal2 39146 14450 39146 14450 0 _1090_
rlabel metal1 39468 12750 39468 12750 0 _1091_
rlabel metal1 39560 12818 39560 12818 0 _1092_
rlabel metal1 6808 14042 6808 14042 0 _1093_
rlabel metal1 5382 13940 5382 13940 0 _1094_
rlabel metal2 5658 15402 5658 15402 0 _1095_
rlabel metal1 38180 11730 38180 11730 0 _1096_
rlabel metal1 33626 6766 33626 6766 0 _1097_
rlabel metal1 33902 8432 33902 8432 0 _1098_
rlabel metal2 41722 22202 41722 22202 0 _1099_
rlabel metal2 18538 33252 18538 33252 0 _1100_
rlabel metal1 20976 33966 20976 33966 0 _1101_
rlabel metal1 20056 32946 20056 32946 0 _1102_
rlabel metal1 20562 32912 20562 32912 0 _1103_
rlabel metal1 20560 33490 20560 33490 0 _1104_
rlabel metal1 20010 32810 20010 32810 0 _1105_
rlabel metal1 19274 33456 19274 33456 0 _1106_
rlabel metal1 12926 34578 12926 34578 0 _1107_
rlabel metal2 12742 34374 12742 34374 0 _1108_
rlabel metal1 13432 32878 13432 32878 0 _1109_
rlabel metal1 14260 33966 14260 33966 0 _1110_
rlabel metal1 13800 33082 13800 33082 0 _1111_
rlabel metal2 12512 41718 12512 41718 0 _1112_
rlabel metal2 11638 34170 11638 34170 0 _1113_
rlabel metal2 12466 33031 12466 33031 0 _1114_
rlabel metal2 13018 33932 13018 33932 0 _1115_
rlabel metal2 12466 33745 12466 33745 0 _1116_
rlabel via2 11914 33507 11914 33507 0 _1117_
rlabel metal1 13386 34136 13386 34136 0 _1118_
rlabel metal1 13064 32878 13064 32878 0 _1119_
rlabel metal1 16054 32742 16054 32742 0 _1120_
rlabel metal2 19504 32844 19504 32844 0 _1121_
rlabel metal1 20700 31790 20700 31790 0 _1122_
rlabel metal1 20654 31994 20654 31994 0 _1123_
rlabel metal1 21804 29206 21804 29206 0 _1124_
rlabel metal1 20700 28526 20700 28526 0 _1125_
rlabel metal1 20470 29274 20470 29274 0 _1126_
rlabel metal1 19872 27982 19872 27982 0 _1127_
rlabel metal1 20378 27846 20378 27846 0 _1128_
rlabel metal1 20194 27642 20194 27642 0 _1129_
rlabel metal1 19964 28526 19964 28526 0 _1130_
rlabel metal1 20148 28458 20148 28458 0 _1131_
rlabel metal1 19964 29138 19964 29138 0 _1132_
rlabel metal2 20286 29444 20286 29444 0 _1133_
rlabel metal1 20746 30226 20746 30226 0 _1134_
rlabel metal1 20884 31858 20884 31858 0 _1135_
rlabel metal1 20470 30872 20470 30872 0 _1136_
rlabel metal2 19458 30090 19458 30090 0 _1137_
rlabel metal1 19688 30158 19688 30158 0 _1138_
rlabel metal1 19550 30226 19550 30226 0 _1139_
rlabel metal2 19366 30668 19366 30668 0 _1140_
rlabel metal1 19918 30090 19918 30090 0 _1141_
rlabel metal1 20516 31926 20516 31926 0 _1142_
rlabel metal1 12098 33524 12098 33524 0 _1143_
rlabel metal1 12742 34000 12742 34000 0 _1144_
rlabel metal2 13846 33150 13846 33150 0 _1145_
rlabel metal2 19366 33796 19366 33796 0 _1146_
rlabel metal1 19918 33490 19918 33490 0 _1147_
rlabel metal1 19964 33286 19964 33286 0 _1148_
rlabel metal2 21344 32436 21344 32436 0 _1149_
rlabel metal2 19734 30804 19734 30804 0 _1150_
rlabel metal1 20746 30906 20746 30906 0 _1151_
rlabel metal1 20516 30362 20516 30362 0 _1152_
rlabel metal1 19872 30634 19872 30634 0 _1153_
rlabel metal2 20102 31008 20102 31008 0 _1154_
rlabel metal2 21574 30821 21574 30821 0 _1155_
rlabel metal1 41032 21454 41032 21454 0 _1156_
rlabel metal2 40158 20672 40158 20672 0 _1157_
rlabel metal1 40158 21114 40158 21114 0 _1158_
rlabel metal1 40848 21522 40848 21522 0 _1159_
rlabel metal1 39514 19414 39514 19414 0 _1160_
rlabel metal1 39698 21522 39698 21522 0 _1161_
rlabel metal1 38916 20026 38916 20026 0 _1162_
rlabel metal1 40388 20910 40388 20910 0 _1163_
rlabel metal1 39836 20774 39836 20774 0 _1164_
rlabel metal1 39422 20910 39422 20910 0 _1165_
rlabel metal2 40572 22100 40572 22100 0 _1166_
rlabel metal1 40802 18802 40802 18802 0 _1167_
rlabel metal2 43194 23596 43194 23596 0 _1168_
rlabel metal1 42780 22950 42780 22950 0 _1169_
rlabel metal1 42458 18802 42458 18802 0 _1170_
rlabel metal1 43332 20978 43332 20978 0 _1171_
rlabel metal2 43194 21216 43194 21216 0 _1172_
rlabel metal1 43010 20978 43010 20978 0 _1173_
rlabel metal1 42872 19346 42872 19346 0 _1174_
rlabel metal1 42964 19822 42964 19822 0 _1175_
rlabel metal1 42642 19448 42642 19448 0 _1176_
rlabel metal1 43562 19380 43562 19380 0 _1177_
rlabel metal1 42550 19346 42550 19346 0 _1178_
rlabel metal1 42964 18734 42964 18734 0 _1179_
rlabel metal1 41354 18768 41354 18768 0 _1180_
rlabel metal1 43010 23630 43010 23630 0 _1181_
rlabel metal1 42044 21522 42044 21522 0 _1182_
rlabel metal2 41998 20060 41998 20060 0 _1183_
rlabel metal1 41308 18394 41308 18394 0 _1184_
rlabel metal1 41584 18734 41584 18734 0 _1185_
rlabel metal1 39330 18224 39330 18224 0 _1186_
rlabel metal1 39698 22576 39698 22576 0 _1187_
rlabel metal2 39974 22032 39974 22032 0 _1188_
rlabel metal2 39330 20094 39330 20094 0 _1189_
rlabel metal1 39146 18292 39146 18292 0 _1190_
rlabel metal1 39376 20366 39376 20366 0 _1191_
rlabel metal1 39192 20434 39192 20434 0 _1192_
rlabel metal2 39054 20740 39054 20740 0 _1193_
rlabel metal1 38916 18258 38916 18258 0 _1194_
rlabel metal1 38732 18258 38732 18258 0 _1195_
rlabel metal1 39008 13362 39008 13362 0 _1196_
rlabel metal1 39100 13158 39100 13158 0 _1197_
rlabel metal2 38732 12954 38732 12954 0 _1198_
rlabel metal1 30728 10710 30728 10710 0 _1199_
rlabel metal1 32246 12818 32246 12818 0 _1200_
rlabel metal2 32890 12852 32890 12852 0 _1201_
rlabel metal2 32706 13294 32706 13294 0 _1202_
rlabel metal1 35880 12614 35880 12614 0 _1203_
rlabel metal1 41078 13362 41078 13362 0 _1204_
rlabel metal1 22816 4998 22816 4998 0 _1205_
rlabel metal1 22586 9044 22586 9044 0 _1206_
rlabel metal1 21942 9588 21942 9588 0 _1207_
rlabel metal1 23138 13260 23138 13260 0 _1208_
rlabel metal1 22724 3026 22724 3026 0 _1209_
rlabel metal1 33166 4726 33166 4726 0 _1210_
rlabel metal1 23690 4624 23690 4624 0 _1211_
rlabel metal2 23598 3808 23598 3808 0 _1212_
rlabel metal1 22770 2890 22770 2890 0 _1213_
rlabel metal1 26584 5202 26584 5202 0 _1214_
rlabel metal1 25300 12682 25300 12682 0 _1215_
rlabel metal1 24426 4114 24426 4114 0 _1216_
rlabel metal1 23874 4114 23874 4114 0 _1217_
rlabel metal2 23506 3009 23506 3009 0 _1218_
rlabel metal1 22770 3366 22770 3366 0 _1219_
rlabel metal1 23230 4556 23230 4556 0 _1220_
rlabel metal1 22816 4250 22816 4250 0 _1221_
rlabel metal1 22586 3536 22586 3536 0 _1222_
rlabel metal1 22540 5678 22540 5678 0 _1223_
rlabel metal2 22586 13532 22586 13532 0 _1224_
rlabel metal1 34270 21386 34270 21386 0 _1225_
rlabel metal1 33994 23630 33994 23630 0 _1226_
rlabel metal1 33902 23766 33902 23766 0 _1227_
rlabel metal1 34592 29002 34592 29002 0 _1228_
rlabel metal1 26358 22032 26358 22032 0 _1229_
rlabel metal1 32936 23290 32936 23290 0 _1230_
rlabel metal1 33128 22950 33128 22950 0 _1231_
rlabel metal1 34086 23188 34086 23188 0 _1232_
rlabel metal2 33902 22848 33902 22848 0 _1233_
rlabel metal1 34638 22542 34638 22542 0 _1234_
rlabel metal2 34730 22202 34730 22202 0 _1235_
rlabel metal1 34454 21556 34454 21556 0 _1236_
rlabel metal1 34040 20910 34040 20910 0 _1237_
rlabel metal1 32476 20978 32476 20978 0 _1238_
rlabel metal2 33074 4828 33074 4828 0 clk
rlabel via2 14766 12835 14766 12835 0 clknet_0_clk
rlabel metal2 21758 8262 21758 8262 0 clknet_2_0__leaf_clk
rlabel metal2 42550 10880 42550 10880 0 clknet_2_1__leaf_clk
rlabel metal1 19228 37230 19228 37230 0 clknet_2_2__leaf_clk
rlabel metal1 38410 39032 38410 39032 0 clknet_2_3__leaf_clk
rlabel metal2 12466 18428 12466 18428 0 clknet_leaf_0_clk
rlabel metal1 15824 34170 15824 34170 0 clknet_leaf_10_clk
rlabel metal1 21436 26418 21436 26418 0 clknet_leaf_11_clk
rlabel metal2 28658 34340 28658 34340 0 clknet_leaf_12_clk
rlabel metal1 24748 42126 24748 42126 0 clknet_leaf_13_clk
rlabel metal1 31280 43758 31280 43758 0 clknet_leaf_14_clk
rlabel metal1 34914 38318 34914 38318 0 clknet_leaf_15_clk
rlabel metal1 42504 41650 42504 41650 0 clknet_leaf_16_clk
rlabel metal1 39468 38862 39468 38862 0 clknet_leaf_17_clk
rlabel metal1 40848 29614 40848 29614 0 clknet_leaf_18_clk
rlabel metal1 39882 26316 39882 26316 0 clknet_leaf_19_clk
rlabel metal1 17112 21658 17112 21658 0 clknet_leaf_1_clk
rlabel metal2 31970 27064 31970 27064 0 clknet_leaf_20_clk
rlabel metal1 30774 21318 30774 21318 0 clknet_leaf_21_clk
rlabel metal1 32568 15470 32568 15470 0 clknet_leaf_22_clk
rlabel metal1 37766 23596 37766 23596 0 clknet_leaf_23_clk
rlabel metal2 39974 16082 39974 16082 0 clknet_leaf_24_clk
rlabel metal1 38686 13260 38686 13260 0 clknet_leaf_25_clk
rlabel metal1 44298 8500 44298 8500 0 clknet_leaf_26_clk
rlabel metal1 36432 7718 36432 7718 0 clknet_leaf_27_clk
rlabel via1 33166 9010 33166 9010 0 clknet_leaf_28_clk
rlabel metal1 24472 3026 24472 3026 0 clknet_leaf_29_clk
rlabel metal1 13984 25806 13984 25806 0 clknet_leaf_2_clk
rlabel metal1 32246 13226 32246 13226 0 clknet_leaf_30_clk
rlabel metal1 19918 18122 19918 18122 0 clknet_leaf_31_clk
rlabel metal1 18400 17102 18400 17102 0 clknet_leaf_32_clk
rlabel metal1 20148 4114 20148 4114 0 clknet_leaf_33_clk
rlabel metal1 7268 4114 7268 4114 0 clknet_leaf_34_clk
rlabel metal1 4738 13362 4738 13362 0 clknet_leaf_35_clk
rlabel metal1 3404 14994 3404 14994 0 clknet_leaf_36_clk
rlabel metal1 6900 21318 6900 21318 0 clknet_leaf_37_clk
rlabel metal1 6532 25806 6532 25806 0 clknet_leaf_3_clk
rlabel metal1 9292 31790 9292 31790 0 clknet_leaf_4_clk
rlabel metal1 9062 34612 9062 34612 0 clknet_leaf_5_clk
rlabel metal1 8832 40494 8832 40494 0 clknet_leaf_6_clk
rlabel metal2 14030 36482 14030 36482 0 clknet_leaf_7_clk
rlabel metal1 18906 39474 18906 39474 0 clknet_leaf_8_clk
rlabel metal1 17020 35122 17020 35122 0 clknet_leaf_9_clk
rlabel metal1 44482 43690 44482 43690 0 cs
rlabel metal2 41262 46284 41262 46284 0 gpio[0]
rlabel metal2 23966 45499 23966 45499 0 gpio[10]
rlabel metal3 820 8908 820 8908 0 gpio[11]
rlabel metal3 820 18428 820 18428 0 gpio[12]
rlabel metal3 44536 6868 44536 6868 0 gpio[13]
rlabel metal3 820 36788 820 36788 0 gpio[14]
rlabel metal1 44482 33966 44482 33966 0 gpio[15]
rlabel metal2 46 1588 46 1588 0 gpio[16]
rlabel metal2 8418 1027 8418 1027 0 gpio[1]
rlabel metal2 43194 1588 43194 1588 0 gpio[2]
rlabel metal2 17434 1027 17434 1027 0 gpio[3]
rlabel metal1 14904 45458 14904 45458 0 gpio[4]
rlabel metal1 44482 24786 44482 24786 0 gpio[5]
rlabel metal3 1050 45628 1050 45628 0 gpio[6]
rlabel metal1 32384 45458 32384 45458 0 gpio[7]
rlabel metal2 25806 823 25806 823 0 gpio[8]
rlabel metal3 820 27268 820 27268 0 gpio[9]
rlabel metal1 33948 4590 33948 4590 0 inputs.down.det_edge
rlabel metal1 32791 5882 32791 5882 0 inputs.down.ff_in
rlabel metal2 33442 7276 33442 7276 0 inputs.down.ff_out
rlabel metal1 34316 7786 34316 7786 0 inputs.down.in
rlabel metal1 9062 5304 9062 5304 0 inputs.frequency_lut.rng\[0\]
rlabel via1 9890 6290 9890 6290 0 inputs.frequency_lut.rng\[1\]
rlabel metal1 9430 4080 9430 4080 0 inputs.frequency_lut.rng\[2\]
rlabel metal1 9775 8466 9775 8466 0 inputs.frequency_lut.rng\[3\]
rlabel metal2 9706 11424 9706 11424 0 inputs.frequency_lut.rng\[4\]
rlabel metal1 10465 12750 10465 12750 0 inputs.frequency_lut.rng\[5\]
rlabel metal1 38272 11186 38272 11186 0 inputs.key_encoder.mode_key
rlabel metal1 41998 11254 41998 11254 0 inputs.key_encoder.octave_key_up
rlabel metal1 32522 12750 32522 12750 0 inputs.key_encoder.sync_keys\[0\]
rlabel metal2 29210 12988 29210 12988 0 inputs.key_encoder.sync_keys\[10\]
rlabel metal1 30222 12818 30222 12818 0 inputs.key_encoder.sync_keys\[11\]
rlabel metal1 17434 18836 17434 18836 0 inputs.key_encoder.sync_keys\[12\]
rlabel metal1 33074 12750 33074 12750 0 inputs.key_encoder.sync_keys\[13\]
rlabel metal1 37904 10234 37904 10234 0 inputs.key_encoder.sync_keys\[14\]
rlabel metal1 34730 12274 34730 12274 0 inputs.key_encoder.sync_keys\[15\]
rlabel metal2 32154 8840 32154 8840 0 inputs.key_encoder.sync_keys\[1\]
rlabel metal1 31510 5100 31510 5100 0 inputs.key_encoder.sync_keys\[2\]
rlabel metal1 31004 5202 31004 5202 0 inputs.key_encoder.sync_keys\[3\]
rlabel metal1 31004 43078 31004 43078 0 inputs.key_encoder.sync_keys\[4\]
rlabel metal1 34546 15606 34546 15606 0 inputs.key_encoder.sync_keys\[5\]
rlabel metal1 17250 14858 17250 14858 0 inputs.key_encoder.sync_keys\[6\]
rlabel metal1 31602 41990 31602 41990 0 inputs.key_encoder.sync_keys\[7\]
rlabel metal1 30176 13294 30176 13294 0 inputs.key_encoder.sync_keys\[8\]
rlabel metal2 13662 15742 13662 15742 0 inputs.key_encoder.sync_keys\[9\]
rlabel metal2 36386 43996 36386 43996 0 inputs.keypad\[0\]
rlabel metal1 25346 42296 25346 42296 0 inputs.keypad\[10\]
rlabel metal1 2714 9656 2714 9656 0 inputs.keypad\[11\]
rlabel metal1 2990 18394 2990 18394 0 inputs.keypad\[12\]
rlabel metal1 3496 6358 3496 6358 0 inputs.keypad\[13\]
rlabel metal1 43792 8058 43792 8058 0 inputs.keypad\[14\]
rlabel metal1 3496 35802 3496 35802 0 inputs.keypad\[15\]
rlabel metal1 43102 31858 43102 31858 0 inputs.keypad\[16\]
rlabel metal1 9246 3128 9246 3128 0 inputs.keypad\[1\]
rlabel metal1 36570 3706 36570 3706 0 inputs.keypad\[2\]
rlabel metal1 19734 2958 19734 2958 0 inputs.keypad\[3\]
rlabel metal1 20194 44472 20194 44472 0 inputs.keypad\[4\]
rlabel metal1 36846 23800 36846 23800 0 inputs.keypad\[5\]
rlabel metal1 6992 43690 6992 43690 0 inputs.keypad\[6\]
rlabel metal1 31648 43826 31648 43826 0 inputs.keypad\[7\]
rlabel metal1 27094 3434 27094 3434 0 inputs.keypad\[8\]
rlabel metal1 6164 25330 6164 25330 0 inputs.keypad\[9\]
rlabel metal2 37996 38692 37996 38692 0 inputs.keypad_synchronizer.half_sync\[0\]
rlabel metal1 26956 41990 26956 41990 0 inputs.keypad_synchronizer.half_sync\[10\]
rlabel metal1 4876 9690 4876 9690 0 inputs.keypad_synchronizer.half_sync\[11\]
rlabel metal1 6670 19312 6670 19312 0 inputs.keypad_synchronizer.half_sync\[12\]
rlabel metal1 11914 6324 11914 6324 0 inputs.keypad_synchronizer.half_sync\[13\]
rlabel metal1 42044 8602 42044 8602 0 inputs.keypad_synchronizer.half_sync\[14\]
rlabel metal2 14720 31484 14720 31484 0 inputs.keypad_synchronizer.half_sync\[15\]
rlabel metal1 44252 22066 44252 22066 0 inputs.keypad_synchronizer.half_sync\[16\]
rlabel metal1 15272 2482 15272 2482 0 inputs.keypad_synchronizer.half_sync\[1\]
rlabel metal1 35006 4250 35006 4250 0 inputs.keypad_synchronizer.half_sync\[2\]
rlabel metal1 22770 3128 22770 3128 0 inputs.keypad_synchronizer.half_sync\[3\]
rlabel metal2 25438 43996 25438 43996 0 inputs.keypad_synchronizer.half_sync\[4\]
rlabel metal1 37122 20978 37122 20978 0 inputs.keypad_synchronizer.half_sync\[5\]
rlabel metal2 8740 39916 8740 39916 0 inputs.keypad_synchronizer.half_sync\[6\]
rlabel metal1 33442 43350 33442 43350 0 inputs.keypad_synchronizer.half_sync\[7\]
rlabel metal1 28888 3706 28888 3706 0 inputs.keypad_synchronizer.half_sync\[8\]
rlabel metal1 8648 20978 8648 20978 0 inputs.keypad_synchronizer.half_sync\[9\]
rlabel metal1 39146 12920 39146 12920 0 inputs.mode_edge.det_edge
rlabel metal1 37720 11866 37720 11866 0 inputs.mode_edge.ff_in
rlabel metal1 39284 10778 39284 10778 0 inputs.mode_edge.ff_out
rlabel metal1 34822 4760 34822 4760 0 inputs.octave_fsm.octave_key_up
rlabel metal1 25944 5066 25944 5066 0 inputs.octave_fsm.state\[0\]
rlabel metal1 24242 5678 24242 5678 0 inputs.octave_fsm.state\[1\]
rlabel metal1 23138 3468 23138 3468 0 inputs.octave_fsm.state\[2\]
rlabel metal1 6348 15130 6348 15130 0 inputs.random_note_generator.feedback
rlabel via1 5405 15674 5405 15674 0 inputs.random_note_generator.out\[0\]
rlabel metal1 6555 16014 6555 16014 0 inputs.random_note_generator.out\[10\]
rlabel metal1 4002 15538 4002 15538 0 inputs.random_note_generator.out\[11\]
rlabel metal1 5290 14450 5290 14450 0 inputs.random_note_generator.out\[12\]
rlabel metal2 4646 13396 4646 13396 0 inputs.random_note_generator.out\[13\]
rlabel metal2 6946 12988 6946 12988 0 inputs.random_note_generator.out\[14\]
rlabel metal1 7567 13498 7567 13498 0 inputs.random_note_generator.out\[15\]
rlabel metal2 2806 16932 2806 16932 0 inputs.random_note_generator.out\[1\]
rlabel metal1 5359 18190 5359 18190 0 inputs.random_note_generator.out\[2\]
rlabel metal1 4554 17170 4554 17170 0 inputs.random_note_generator.out\[3\]
rlabel metal1 7245 18938 7245 18938 0 inputs.random_note_generator.out\[4\]
rlabel metal1 8694 18394 8694 18394 0 inputs.random_note_generator.out\[5\]
rlabel metal1 8142 17646 8142 17646 0 inputs.random_note_generator.out\[6\]
rlabel metal1 9706 17102 9706 17102 0 inputs.random_note_generator.out\[7\]
rlabel metal2 8970 16932 8970 16932 0 inputs.random_note_generator.out\[8\]
rlabel metal1 8740 17714 8740 17714 0 inputs.random_note_generator.out\[9\]
rlabel metal1 35006 40460 35006 40460 0 inputs.random_update_clock.count\[0\]
rlabel metal1 38962 41242 38962 41242 0 inputs.random_update_clock.count\[10\]
rlabel metal1 40618 42738 40618 42738 0 inputs.random_update_clock.count\[11\]
rlabel metal1 41998 41990 41998 41990 0 inputs.random_update_clock.count\[12\]
rlabel metal1 41722 41514 41722 41514 0 inputs.random_update_clock.count\[13\]
rlabel metal1 44206 41446 44206 41446 0 inputs.random_update_clock.count\[14\]
rlabel metal1 42642 39610 42642 39610 0 inputs.random_update_clock.count\[15\]
rlabel metal2 39514 34544 39514 34544 0 inputs.random_update_clock.count\[16\]
rlabel metal1 40986 35190 40986 35190 0 inputs.random_update_clock.count\[17\]
rlabel metal1 40940 34034 40940 34034 0 inputs.random_update_clock.count\[18\]
rlabel metal2 42090 33796 42090 33796 0 inputs.random_update_clock.count\[19\]
rlabel metal1 36846 40426 36846 40426 0 inputs.random_update_clock.count\[1\]
rlabel metal2 42734 35632 42734 35632 0 inputs.random_update_clock.count\[20\]
rlabel metal1 43056 36142 43056 36142 0 inputs.random_update_clock.count\[21\]
rlabel metal1 42872 37094 42872 37094 0 inputs.random_update_clock.count\[22\]
rlabel metal1 36662 41038 36662 41038 0 inputs.random_update_clock.count\[2\]
rlabel metal1 36202 40494 36202 40494 0 inputs.random_update_clock.count\[3\]
rlabel metal2 36754 38046 36754 38046 0 inputs.random_update_clock.count\[4\]
rlabel metal1 37260 37842 37260 37842 0 inputs.random_update_clock.count\[5\]
rlabel metal1 39008 36686 39008 36686 0 inputs.random_update_clock.count\[6\]
rlabel metal1 37352 37774 37352 37774 0 inputs.random_update_clock.count\[7\]
rlabel metal1 40848 38930 40848 38930 0 inputs.random_update_clock.count\[8\]
rlabel metal2 40618 40256 40618 40256 0 inputs.random_update_clock.count\[9\]
rlabel metal1 33580 41242 33580 41242 0 inputs.random_update_clock.next_count\[0\]
rlabel metal1 37812 40698 37812 40698 0 inputs.random_update_clock.next_count\[10\]
rlabel metal1 39146 42874 39146 42874 0 inputs.random_update_clock.next_count\[11\]
rlabel metal1 40158 42296 40158 42296 0 inputs.random_update_clock.next_count\[12\]
rlabel metal1 42504 42262 42504 42262 0 inputs.random_update_clock.next_count\[13\]
rlabel metal1 43102 41650 43102 41650 0 inputs.random_update_clock.next_count\[14\]
rlabel metal1 42458 39338 42458 39338 0 inputs.random_update_clock.next_count\[15\]
rlabel metal1 38134 33864 38134 33864 0 inputs.random_update_clock.next_count\[16\]
rlabel metal1 39836 36006 39836 36006 0 inputs.random_update_clock.next_count\[17\]
rlabel metal2 40158 33252 40158 33252 0 inputs.random_update_clock.next_count\[18\]
rlabel metal1 42918 34034 42918 34034 0 inputs.random_update_clock.next_count\[19\]
rlabel metal2 35006 42364 35006 42364 0 inputs.random_update_clock.next_count\[1\]
rlabel metal1 43884 34646 43884 34646 0 inputs.random_update_clock.next_count\[20\]
rlabel metal1 42274 36686 42274 36686 0 inputs.random_update_clock.next_count\[21\]
rlabel metal1 43286 37842 43286 37842 0 inputs.random_update_clock.next_count\[22\]
rlabel metal1 36087 41242 36087 41242 0 inputs.random_update_clock.next_count\[2\]
rlabel metal1 34822 39610 34822 39610 0 inputs.random_update_clock.next_count\[3\]
rlabel metal1 35328 37774 35328 37774 0 inputs.random_update_clock.next_count\[4\]
rlabel metal2 35374 37026 35374 37026 0 inputs.random_update_clock.next_count\[5\]
rlabel metal1 37582 36210 37582 36210 0 inputs.random_update_clock.next_count\[6\]
rlabel metal1 38456 38862 38456 38862 0 inputs.random_update_clock.next_count\[7\]
rlabel metal1 40204 37978 40204 37978 0 inputs.random_update_clock.next_count\[8\]
rlabel metal1 39100 39610 39100 39610 0 inputs.random_update_clock.next_count\[9\]
rlabel metal1 33212 5270 33212 5270 0 inputs.up.ff_in
rlabel metal1 34500 8534 34500 8534 0 inputs.up.ff_out
rlabel metal1 39974 12954 39974 12954 0 inputs.wavetype_fsm.next_state\[0\]
rlabel metal1 38916 15470 38916 15470 0 inputs.wavetype_fsm.next_state\[1\]
rlabel metal1 39330 12750 39330 12750 0 inputs.wavetype_fsm.state\[0\]
rlabel metal1 39468 15470 39468 15470 0 inputs.wavetype_fsm.state\[1\]
rlabel metal2 1794 36958 1794 36958 0 net1
rlabel metal1 8602 2890 8602 2890 0 net10
rlabel metal2 43102 16830 43102 16830 0 net100
rlabel metal1 19320 34714 19320 34714 0 net101
rlabel metal1 17480 34714 17480 34714 0 net102
rlabel metal1 13938 43622 13938 43622 0 net103
rlabel metal1 12788 43350 12788 43350 0 net104
rlabel metal1 17940 29274 17940 29274 0 net105
rlabel metal1 20286 43214 20286 43214 0 net106
rlabel metal2 18446 43418 18446 43418 0 net107
rlabel metal2 23506 34204 23506 34204 0 net108
rlabel metal1 23460 33558 23460 33558 0 net109
rlabel metal2 43286 2754 43286 2754 0 net11
rlabel metal1 23184 28390 23184 28390 0 net110
rlabel metal1 22402 39270 22402 39270 0 net111
rlabel metal2 12006 43826 12006 43826 0 net112
rlabel metal1 11224 43418 11224 43418 0 net113
rlabel metal1 17480 43962 17480 43962 0 net114
rlabel metal1 15686 43418 15686 43418 0 net115
rlabel metal1 10350 38250 10350 38250 0 net116
rlabel metal1 9706 37944 9706 37944 0 net117
rlabel metal2 42642 38148 42642 38148 0 net118
rlabel metal1 44344 37298 44344 37298 0 net119
rlabel metal1 18354 2618 18354 2618 0 net12
rlabel metal1 18952 36618 18952 36618 0 net120
rlabel metal2 17342 37026 17342 37026 0 net121
rlabel metal1 23138 26010 23138 26010 0 net122
rlabel metal1 23552 37162 23552 37162 0 net123
rlabel metal1 23184 36210 23184 36210 0 net124
rlabel metal1 18078 28186 18078 28186 0 net125
rlabel metal1 22264 40154 22264 40154 0 net126
rlabel metal1 23782 40562 23782 40562 0 net127
rlabel metal1 20332 25262 20332 25262 0 net128
rlabel metal1 13662 37230 13662 37230 0 net129
rlabel metal1 18722 45016 18722 45016 0 net13
rlabel metal1 13754 36856 13754 36856 0 net130
rlabel metal2 10994 39712 10994 39712 0 net131
rlabel metal1 9844 40154 9844 40154 0 net132
rlabel metal1 36616 6222 36616 6222 0 net133
rlabel metal2 32522 18462 32522 18462 0 net134
rlabel metal1 20010 40902 20010 40902 0 net135
rlabel metal1 18952 40086 18952 40086 0 net136
rlabel via1 13386 39066 13386 39066 0 net137
rlabel metal1 11868 39474 11868 39474 0 net138
rlabel metal1 36110 10710 36110 10710 0 net139
rlabel metal1 40342 24650 40342 24650 0 net14
rlabel metal1 35374 11866 35374 11866 0 net140
rlabel via1 16790 41582 16790 41582 0 net141
rlabel metal1 18124 42330 18124 42330 0 net142
rlabel metal1 12540 40494 12540 40494 0 net143
rlabel metal1 13570 41174 13570 41174 0 net144
rlabel metal1 34362 11186 34362 11186 0 net145
rlabel metal1 36478 10642 36478 10642 0 net146
rlabel metal1 37490 10710 37490 10710 0 net147
rlabel metal1 38134 6834 38134 6834 0 net148
rlabel metal1 38870 11526 38870 11526 0 net149
rlabel metal2 5934 45118 5934 45118 0 net15
rlabel metal1 16100 38182 16100 38182 0 net150
rlabel metal1 14490 38862 14490 38862 0 net151
rlabel metal1 37628 8942 37628 8942 0 net152
rlabel metal1 43010 15028 43010 15028 0 net153
rlabel metal2 43102 30464 43102 30464 0 net154
rlabel metal1 41216 29682 41216 29682 0 net155
rlabel metal1 38088 8058 38088 8058 0 net156
rlabel metal1 37214 8466 37214 8466 0 net157
rlabel metal1 35926 7310 35926 7310 0 net158
rlabel via1 26266 14858 26266 14858 0 net159
rlabel metal1 32154 44982 32154 44982 0 net16
rlabel metal1 42780 27506 42780 27506 0 net160
rlabel metal1 40940 28186 40940 28186 0 net161
rlabel metal1 40526 25262 40526 25262 0 net162
rlabel metal1 38456 25466 38456 25466 0 net163
rlabel metal1 41285 31790 41285 31790 0 net164
rlabel metal2 40618 31076 40618 31076 0 net165
rlabel metal1 30452 28526 30452 28526 0 net166
rlabel metal2 18998 36924 18998 36924 0 net167
rlabel metal1 20286 37774 20286 37774 0 net168
rlabel metal1 34362 41106 34362 41106 0 net169
rlabel metal1 26082 2550 26082 2550 0 net17
rlabel metal1 40894 26894 40894 26894 0 net170
rlabel metal1 42083 26554 42083 26554 0 net171
rlabel metal1 32890 30260 32890 30260 0 net172
rlabel metal1 34362 23732 34362 23732 0 net173
rlabel metal2 41078 24548 41078 24548 0 net174
rlabel metal2 40158 26588 40158 26588 0 net175
rlabel metal1 27692 37774 27692 37774 0 net176
rlabel metal1 37858 18258 37858 18258 0 net177
rlabel metal1 18520 42194 18520 42194 0 net178
rlabel metal1 19642 41786 19642 41786 0 net179
rlabel metal2 1610 26928 1610 26928 0 net18
rlabel metal1 30130 22610 30130 22610 0 net180
rlabel metal2 29486 27132 29486 27132 0 net181
rlabel metal1 34316 16014 34316 16014 0 net182
rlabel metal1 25070 32742 25070 32742 0 net183
rlabel metal2 26542 33320 26542 33320 0 net184
rlabel metal1 43010 40528 43010 40528 0 net185
rlabel metal1 43424 40494 43424 40494 0 net186
rlabel via1 15042 42194 15042 42194 0 net187
rlabel metal1 30360 36142 30360 36142 0 net188
rlabel via1 24868 31790 24868 31790 0 net189
rlabel metal2 27370 43248 27370 43248 0 net19
rlabel metal1 29992 16014 29992 16014 0 net190
rlabel metal1 32844 16014 32844 16014 0 net191
rlabel metal2 28842 19618 28842 19618 0 net192
rlabel viali 13110 41582 13110 41582 0 net193
rlabel metal1 13754 41786 13754 41786 0 net194
rlabel metal1 27094 31246 27094 31246 0 net195
rlabel metal1 17232 37842 17232 37842 0 net196
rlabel metal1 18262 37978 18262 37978 0 net197
rlabel metal1 37904 26554 37904 26554 0 net198
rlabel metal1 36977 25466 36977 25466 0 net199
rlabel metal1 39100 44982 39100 44982 0 net2
rlabel metal1 43792 15130 43792 15130 0 net20
rlabel metal2 35926 38250 35926 38250 0 net200
rlabel viali 20930 41582 20930 41582 0 net201
rlabel metal2 35374 40426 35374 40426 0 net202
rlabel metal1 36432 41582 36432 41582 0 net203
rlabel metal1 23948 38930 23948 38930 0 net204
rlabel metal1 25024 38862 25024 38862 0 net205
rlabel metal1 39698 34714 39698 34714 0 net206
rlabel metal1 9016 33830 9016 33830 0 net207
rlabel metal1 25254 35802 25254 35802 0 net208
rlabel metal1 25208 36822 25208 36822 0 net209
rlabel metal1 35742 22168 35742 22168 0 net21
rlabel metal1 34914 21998 34914 21998 0 net210
rlabel metal1 31786 19414 31786 19414 0 net211
rlabel metal1 34730 40562 34730 40562 0 net212
rlabel metal1 40940 39406 40940 39406 0 net213
rlabel metal1 34776 42194 34776 42194 0 net214
rlabel metal1 31924 33558 31924 33558 0 net215
rlabel metal1 34270 26384 34270 26384 0 net216
rlabel metal1 33810 25976 33810 25976 0 net217
rlabel metal1 42090 33898 42090 33898 0 net218
rlabel metal1 37720 20570 37720 20570 0 net219
rlabel metal2 6762 13464 6762 13464 0 net22
rlabel metal1 35788 25942 35788 25942 0 net220
rlabel metal1 39330 42670 39330 42670 0 net221
rlabel metal1 17342 17170 17342 17170 0 net222
rlabel metal1 34960 13906 34960 13906 0 net223
rlabel metal1 32246 25942 32246 25942 0 net224
rlabel metal2 31970 24990 31970 24990 0 net225
rlabel metal1 43148 33966 43148 33966 0 net226
rlabel metal1 43424 40018 43424 40018 0 net227
rlabel metal1 33258 27370 33258 27370 0 net228
rlabel metal1 35374 30192 35374 30192 0 net229
rlabel metal1 20739 5610 20739 5610 0 net23
rlabel metal1 22494 23494 22494 23494 0 net230
rlabel metal1 35696 20910 35696 20910 0 net231
rlabel metal1 24058 25126 24058 25126 0 net232
rlabel metal1 38502 29614 38502 29614 0 net233
rlabel metal1 40434 29240 40434 29240 0 net234
rlabel metal1 28060 34578 28060 34578 0 net235
rlabel metal1 33626 38862 33626 38862 0 net236
rlabel metal1 38410 36754 38410 36754 0 net237
rlabel metal2 32798 39338 32798 39338 0 net238
rlabel metal1 23966 24038 23966 24038 0 net239
rlabel metal1 4777 14994 4777 14994 0 net24
rlabel metal1 21482 17714 21482 17714 0 net240
rlabel metal2 43654 18530 43654 18530 0 net241
rlabel metal1 42458 17748 42458 17748 0 net242
rlabel metal1 31372 37842 31372 37842 0 net243
rlabel metal1 39238 30600 39238 30600 0 net244
rlabel metal1 39882 16116 39882 16116 0 net245
rlabel metal1 29026 38420 29026 38420 0 net246
rlabel metal1 38640 37842 38640 37842 0 net247
rlabel metal1 8602 25262 8602 25262 0 net248
rlabel metal1 39422 17136 39422 17136 0 net249
rlabel metal1 13846 18149 13846 18149 0 net25
rlabel metal1 39330 16592 39330 16592 0 net250
rlabel metal2 35374 34782 35374 34782 0 net251
rlabel metal1 38824 27438 38824 27438 0 net252
rlabel metal1 40572 28118 40572 28118 0 net253
rlabel metal1 40802 13328 40802 13328 0 net254
rlabel metal1 38180 15062 38180 15062 0 net255
rlabel metal1 14766 20570 14766 20570 0 net256
rlabel metal1 38686 31994 38686 31994 0 net257
rlabel metal1 38042 28390 38042 28390 0 net258
rlabel metal1 35972 28594 35972 28594 0 net259
rlabel metal1 12558 19720 12558 19720 0 net26
rlabel metal1 39192 26962 39192 26962 0 net260
rlabel metal1 42412 17170 42412 17170 0 net261
rlabel metal1 34362 26928 34362 26928 0 net262
rlabel metal1 35420 27098 35420 27098 0 net263
rlabel metal1 17296 33490 17296 33490 0 net264
rlabel metal1 12972 26282 12972 26282 0 net265
rlabel metal1 36708 33558 36708 33558 0 net266
rlabel metal2 18538 31994 18538 31994 0 net267
rlabel metal1 28658 21488 28658 21488 0 net268
rlabel metal1 8234 37230 8234 37230 0 net269
rlabel metal1 18867 18666 18867 18666 0 net27
rlabel metal1 15502 33626 15502 33626 0 net270
rlabel metal2 29026 29716 29026 29716 0 net271
rlabel metal1 8280 38930 8280 38930 0 net272
rlabel metal2 20010 16320 20010 16320 0 net273
rlabel metal1 12098 28186 12098 28186 0 net274
rlabel metal1 12144 42194 12144 42194 0 net275
rlabel metal1 8924 40154 8924 40154 0 net276
rlabel metal1 15180 37162 15180 37162 0 net277
rlabel metal1 35558 18666 35558 18666 0 net278
rlabel metal1 15364 27438 15364 27438 0 net279
rlabel metal1 19649 19346 19649 19346 0 net28
rlabel metal2 21942 18224 21942 18224 0 net280
rlabel metal1 14858 26350 14858 26350 0 net281
rlabel metal2 15134 15674 15134 15674 0 net282
rlabel metal1 19918 18598 19918 18598 0 net283
rlabel metal1 16192 41174 16192 41174 0 net284
rlabel metal1 13202 16762 13202 16762 0 net285
rlabel metal1 16376 19482 16376 19482 0 net286
rlabel metal1 17158 39338 17158 39338 0 net287
rlabel metal2 12374 19414 12374 19414 0 net288
rlabel metal1 9936 41446 9936 41446 0 net289
rlabel metal2 20378 21046 20378 21046 0 net29
rlabel metal1 16100 35802 16100 35802 0 net290
rlabel metal1 16514 40086 16514 40086 0 net291
rlabel metal1 23276 16966 23276 16966 0 net292
rlabel viali 39699 35054 39699 35054 0 net293
rlabel metal1 24656 15334 24656 15334 0 net294
rlabel metal2 11914 18258 11914 18258 0 net295
rlabel metal1 36110 37842 36110 37842 0 net296
rlabel metal1 20746 24072 20746 24072 0 net297
rlabel metal1 12006 44506 12006 44506 0 net298
rlabel metal2 14490 43962 14490 43962 0 net299
rlabel metal1 24242 45254 24242 45254 0 net3
rlabel metal1 38877 12818 38877 12818 0 net30
rlabel metal1 18308 28050 18308 28050 0 net300
rlabel metal1 13800 35802 13800 35802 0 net301
rlabel metal1 30268 31858 30268 31858 0 net302
rlabel metal1 34730 14348 34730 14348 0 net303
rlabel metal1 20194 36754 20194 36754 0 net304
rlabel metal1 22448 37978 22448 37978 0 net305
rlabel metal1 8418 41684 8418 41684 0 net306
rlabel metal1 6302 28050 6302 28050 0 net307
rlabel metal1 37904 20434 37904 20434 0 net308
rlabel metal1 19872 24106 19872 24106 0 net309
rlabel metal1 42865 8466 42865 8466 0 net31
rlabel metal1 17802 25194 17802 25194 0 net310
rlabel metal1 15180 23086 15180 23086 0 net311
rlabel metal1 23736 30634 23736 30634 0 net312
rlabel metal1 18124 40698 18124 40698 0 net313
rlabel metal1 12650 42738 12650 42738 0 net314
rlabel metal1 16790 28118 16790 28118 0 net315
rlabel metal1 35144 13498 35144 13498 0 net32
rlabel metal1 29118 21862 29118 21862 0 net33
rlabel metal1 36570 14987 36570 14987 0 net34
rlabel metal1 40710 16762 40710 16762 0 net35
rlabel metal1 36294 18224 36294 18224 0 net36
rlabel metal1 36662 24174 36662 24174 0 net37
rlabel metal1 34178 13396 34178 13396 0 net38
rlabel metal2 12466 24684 12466 24684 0 net39
rlabel metal1 1840 9078 1840 9078 0 net4
rlabel metal1 8885 32810 8885 32810 0 net40
rlabel metal1 15824 27574 15824 27574 0 net41
rlabel metal2 21574 33830 21574 33830 0 net42
rlabel metal1 17434 32198 17434 32198 0 net43
rlabel metal2 9614 39168 9614 39168 0 net44
rlabel metal1 11599 36754 11599 36754 0 net45
rlabel metal1 14720 39066 14720 39066 0 net46
rlabel metal2 20654 35258 20654 35258 0 net47
rlabel metal2 16054 39882 16054 39882 0 net48
rlabel metal1 22487 42262 22487 42262 0 net49
rlabel metal1 1840 18870 1840 18870 0 net5
rlabel metal1 8510 42119 8510 42119 0 net50
rlabel metal2 32614 25568 32614 25568 0 net51
rlabel metal2 26266 33014 26266 33014 0 net52
rlabel metal1 34861 25874 34861 25874 0 net53
rlabel metal1 41209 26350 41209 26350 0 net54
rlabel metal1 40296 33286 40296 33286 0 net55
rlabel metal2 37674 33626 37674 33626 0 net56
rlabel metal1 32338 39304 32338 39304 0 net57
rlabel metal1 30314 43241 30314 43241 0 net58
rlabel metal2 38318 38692 38318 38692 0 net59
rlabel metal1 43838 7242 43838 7242 0 net6
rlabel metal1 42550 42092 42550 42092 0 net60
rlabel metal1 36340 38998 36340 38998 0 net61
rlabel metal1 37490 34510 37490 34510 0 net62
rlabel metal1 8556 18326 8556 18326 0 net63
rlabel metal1 33718 42296 33718 42296 0 net64
rlabel metal1 37858 15538 37858 15538 0 net65
rlabel metal1 27232 3706 27232 3706 0 net66
rlabel metal2 40894 9826 40894 9826 0 net67
rlabel metal1 10534 16626 10534 16626 0 net68
rlabel metal1 8556 18734 8556 18734 0 net69
rlabel metal2 2162 36856 2162 36856 0 net7
rlabel metal1 6716 17306 6716 17306 0 net70
rlabel metal1 9246 16184 9246 16184 0 net71
rlabel metal1 32982 4522 32982 4522 0 net72
rlabel metal1 4692 10234 4692 10234 0 net73
rlabel metal1 6210 12954 6210 12954 0 net74
rlabel metal1 42044 14042 42044 14042 0 net75
rlabel metal1 28152 4658 28152 4658 0 net76
rlabel metal1 3772 15062 3772 15062 0 net77
rlabel metal2 29210 43486 29210 43486 0 net78
rlabel metal1 5244 17306 5244 17306 0 net79
rlabel metal1 43930 33014 43930 33014 0 net8
rlabel metal1 8602 16014 8602 16014 0 net80
rlabel metal1 3680 17850 3680 17850 0 net81
rlabel metal1 24656 2482 24656 2482 0 net82
rlabel metal1 8004 17238 8004 17238 0 net83
rlabel metal1 6670 18360 6670 18360 0 net84
rlabel metal1 6026 17578 6026 17578 0 net85
rlabel metal1 19918 5746 19918 5746 0 net86
rlabel metal1 4462 16150 4462 16150 0 net87
rlabel metal1 5888 14246 5888 14246 0 net88
rlabel metal2 43976 11186 43976 11186 0 net89
rlabel metal1 1840 2618 1840 2618 0 net9
rlabel metal2 8970 16660 8970 16660 0 net90
rlabel metal2 4094 13464 4094 13464 0 net91
rlabel metal1 34999 9146 34999 9146 0 net92
rlabel metal1 2162 15368 2162 15368 0 net93
rlabel metal1 38226 13226 38226 13226 0 net94
rlabel metal1 27876 13226 27876 13226 0 net95
rlabel metal1 22816 41514 22816 41514 0 net96
rlabel metal1 24840 39338 24840 39338 0 net97
rlabel metal1 24638 33966 24638 33966 0 net98
rlabel metal2 24518 34782 24518 34782 0 net99
rlabel metal1 6532 45458 6532 45458 0 nrst
rlabel metal1 34914 24242 34914 24242 0 outputs.div.a\[0\]
rlabel metal1 30222 21998 30222 21998 0 outputs.div.a\[10\]
rlabel via1 32154 25262 32154 25262 0 outputs.div.a\[11\]
rlabel metal1 28382 26452 28382 26452 0 outputs.div.a\[12\]
rlabel metal1 32476 26214 32476 26214 0 outputs.div.a\[13\]
rlabel metal1 30498 29104 30498 29104 0 outputs.div.a\[14\]
rlabel metal1 34224 28526 34224 28526 0 outputs.div.a\[15\]
rlabel metal1 33396 30770 33396 30770 0 outputs.div.a\[16\]
rlabel metal1 36041 32334 36041 32334 0 outputs.div.a\[17\]
rlabel metal1 37490 34068 37490 34068 0 outputs.div.a\[18\]
rlabel metal1 34546 35462 34546 35462 0 outputs.div.a\[19\]
rlabel metal2 35558 22039 35558 22039 0 outputs.div.a\[1\]
rlabel metal1 34086 38930 34086 38930 0 outputs.div.a\[20\]
rlabel metal1 32384 39950 32384 39950 0 outputs.div.a\[21\]
rlabel metal1 32154 35700 32154 35700 0 outputs.div.a\[22\]
rlabel metal1 30498 35802 30498 35802 0 outputs.div.a\[23\]
rlabel metal1 31234 33626 31234 33626 0 outputs.div.a\[24\]
rlabel metal1 31188 20978 31188 20978 0 outputs.div.a\[25\]
rlabel metal2 36662 20740 36662 20740 0 outputs.div.a\[2\]
rlabel metal1 34546 18054 34546 18054 0 outputs.div.a\[3\]
rlabel metal1 34362 15504 34362 15504 0 outputs.div.a\[4\]
rlabel metal1 32062 16082 32062 16082 0 outputs.div.a\[5\]
rlabel metal1 30360 16014 30360 16014 0 outputs.div.a\[6\]
rlabel metal1 32246 19346 32246 19346 0 outputs.div.a\[7\]
rlabel metal1 28750 19448 28750 19448 0 outputs.div.a\[8\]
rlabel via1 28106 22609 28106 22609 0 outputs.div.a\[9\]
rlabel metal1 29026 39440 29026 39440 0 outputs.div.count\[0\]
rlabel metal1 30084 38862 30084 38862 0 outputs.div.count\[1\]
rlabel metal1 28060 37774 28060 37774 0 outputs.div.count\[2\]
rlabel metal1 28106 36346 28106 36346 0 outputs.div.count\[3\]
rlabel metal1 28750 34612 28750 34612 0 outputs.div.count\[4\]
rlabel metal1 36478 34680 36478 34680 0 outputs.div.div
rlabel metal1 19918 18734 19918 18734 0 outputs.div.divisor\[0\]
rlabel metal1 13846 16592 13846 16592 0 outputs.div.divisor\[10\]
rlabel metal1 11914 15674 11914 15674 0 outputs.div.divisor\[11\]
rlabel metal1 14122 20026 14122 20026 0 outputs.div.divisor\[12\]
rlabel metal1 16882 19278 16882 19278 0 outputs.div.divisor\[13\]
rlabel metal1 22908 22066 22908 22066 0 outputs.div.divisor\[14\]
rlabel metal1 24426 21114 24426 21114 0 outputs.div.divisor\[15\]
rlabel metal2 24242 24276 24242 24276 0 outputs.div.divisor\[16\]
rlabel metal1 23368 25466 23368 25466 0 outputs.div.divisor\[17\]
rlabel metal1 21758 17714 21758 17714 0 outputs.div.divisor\[1\]
rlabel metal1 17894 16762 17894 16762 0 outputs.div.divisor\[2\]
rlabel metal1 22586 15640 22586 15640 0 outputs.div.divisor\[3\]
rlabel metal1 19872 15130 19872 15130 0 outputs.div.divisor\[4\]
rlabel metal1 24334 15538 24334 15538 0 outputs.div.divisor\[5\]
rlabel metal1 27140 14926 27140 14926 0 outputs.div.divisor\[6\]
rlabel metal1 15364 16014 15364 16014 0 outputs.div.divisor\[7\]
rlabel metal1 23920 17102 23920 17102 0 outputs.div.divisor\[8\]
rlabel metal1 11822 17578 11822 17578 0 outputs.div.divisor\[9\]
rlabel metal1 19550 18666 19550 18666 0 outputs.div.m\[0\]
rlabel metal1 14444 18326 14444 18326 0 outputs.div.m\[10\]
rlabel metal1 16422 22610 16422 22610 0 outputs.div.m\[11\]
rlabel metal1 15962 21454 15962 21454 0 outputs.div.m\[12\]
rlabel metal1 16100 20570 16100 20570 0 outputs.div.m\[13\]
rlabel metal2 19274 24854 19274 24854 0 outputs.div.m\[14\]
rlabel metal1 26358 28186 26358 28186 0 outputs.div.m\[15\]
rlabel metal1 25992 27506 25992 27506 0 outputs.div.m\[16\]
rlabel metal2 25438 26112 25438 26112 0 outputs.div.m\[17\]
rlabel metal1 21988 18734 21988 18734 0 outputs.div.m\[1\]
rlabel metal1 17940 17714 17940 17714 0 outputs.div.m\[2\]
rlabel metal1 21252 19482 21252 19482 0 outputs.div.m\[3\]
rlabel metal2 20470 18462 20470 18462 0 outputs.div.m\[4\]
rlabel metal1 21114 22134 21114 22134 0 outputs.div.m\[5\]
rlabel metal1 26312 17646 26312 17646 0 outputs.div.m\[6\]
rlabel metal1 15410 17102 15410 17102 0 outputs.div.m\[7\]
rlabel metal1 23368 18394 23368 18394 0 outputs.div.m\[8\]
rlabel metal1 17066 20264 17066 20264 0 outputs.div.m\[9\]
rlabel metal1 36616 31790 36616 31790 0 outputs.div.next_div
rlabel metal2 27922 33082 27922 33082 0 outputs.div.next_start
rlabel metal1 13570 25942 13570 25942 0 outputs.div.oscillator_out\[0\]
rlabel metal1 8602 40120 8602 40120 0 outputs.div.oscillator_out\[10\]
rlabel metal1 12673 42126 12673 42126 0 outputs.div.oscillator_out\[11\]
rlabel metal1 11362 42670 11362 42670 0 outputs.div.oscillator_out\[12\]
rlabel metal1 12926 42568 12926 42568 0 outputs.div.oscillator_out\[13\]
rlabel metal1 17480 41106 17480 41106 0 outputs.div.oscillator_out\[14\]
rlabel metal1 18492 39882 18492 39882 0 outputs.div.oscillator_out\[15\]
rlabel metal1 17434 39474 17434 39474 0 outputs.div.oscillator_out\[16\]
rlabel metal1 17480 36210 17480 36210 0 outputs.div.oscillator_out\[17\]
rlabel metal1 16146 26418 16146 26418 0 outputs.div.oscillator_out\[1\]
rlabel metal1 16422 28118 16422 28118 0 outputs.div.oscillator_out\[2\]
rlabel metal1 18768 32334 18768 32334 0 outputs.div.oscillator_out\[3\]
rlabel metal2 12834 28084 12834 28084 0 outputs.div.oscillator_out\[4\]
rlabel metal1 16284 35054 16284 35054 0 outputs.div.oscillator_out\[5\]
rlabel metal1 17342 33082 17342 33082 0 outputs.div.oscillator_out\[6\]
rlabel metal2 16054 37468 16054 37468 0 outputs.div.oscillator_out\[7\]
rlabel metal1 8648 37774 8648 37774 0 outputs.div.oscillator_out\[8\]
rlabel metal1 9016 38386 9016 38386 0 outputs.div.oscillator_out\[9\]
rlabel metal2 38134 30838 38134 30838 0 outputs.div.q\[0\]
rlabel metal1 26542 32334 26542 32334 0 outputs.div.q\[10\]
rlabel metal1 24702 33354 24702 33354 0 outputs.div.q\[11\]
rlabel metal1 26036 34714 26036 34714 0 outputs.div.q\[12\]
rlabel metal2 23874 37060 23874 37060 0 outputs.div.q\[13\]
rlabel metal1 18768 37638 18768 37638 0 outputs.div.q\[14\]
rlabel metal1 16008 38386 16008 38386 0 outputs.div.q\[15\]
rlabel metal2 12834 39508 12834 39508 0 outputs.div.q\[16\]
rlabel metal1 13432 39610 13432 39610 0 outputs.div.q\[17\]
rlabel metal1 12650 40392 12650 40392 0 outputs.div.q\[18\]
rlabel metal2 14858 42772 14858 42772 0 outputs.div.q\[19\]
rlabel metal1 40112 30702 40112 30702 0 outputs.div.q\[1\]
rlabel metal1 17020 42874 17020 42874 0 outputs.div.q\[20\]
rlabel metal1 17756 42534 17756 42534 0 outputs.div.q\[21\]
rlabel metal1 20010 41990 20010 41990 0 outputs.div.q\[22\]
rlabel metal1 24288 41650 24288 41650 0 outputs.div.q\[23\]
rlabel metal1 25898 40052 25898 40052 0 outputs.div.q\[24\]
rlabel metal2 33948 28628 33948 28628 0 outputs.div.q\[25\]
rlabel metal1 35374 26010 35374 26010 0 outputs.div.q\[26\]
rlabel metal1 40802 30090 40802 30090 0 outputs.div.q\[2\]
rlabel metal1 39836 28526 39836 28526 0 outputs.div.q\[3\]
rlabel metal1 40664 27438 40664 27438 0 outputs.div.q\[4\]
rlabel metal1 39652 27982 39652 27982 0 outputs.div.q\[5\]
rlabel metal1 37168 28730 37168 28730 0 outputs.div.q\[6\]
rlabel metal2 34638 28084 34638 28084 0 outputs.div.q\[7\]
rlabel metal1 32982 30804 32982 30804 0 outputs.div.q\[8\]
rlabel metal1 25806 30906 25806 30906 0 outputs.div.q\[9\]
rlabel metal1 42136 31450 42136 31450 0 outputs.div.q_out\[0\]
rlabel metal1 42596 29818 42596 29818 0 outputs.div.q_out\[1\]
rlabel metal1 42550 28730 42550 28730 0 outputs.div.q_out\[2\]
rlabel metal1 43654 26554 43654 26554 0 outputs.div.q_out\[3\]
rlabel metal1 41676 25874 41676 25874 0 outputs.div.q_out\[4\]
rlabel metal1 39928 25806 39928 25806 0 outputs.div.q_out\[5\]
rlabel metal1 38088 25126 38088 25126 0 outputs.div.q_out\[6\]
rlabel metal2 37122 26180 37122 26180 0 outputs.div.q_out\[7\]
rlabel metal1 28520 35666 28520 35666 0 outputs.div.start
rlabel metal1 14950 23834 14950 23834 0 outputs.divider_buffer\[0\]
rlabel metal1 13064 33898 13064 33898 0 outputs.divider_buffer\[10\]
rlabel metal1 11776 33966 11776 33966 0 outputs.divider_buffer\[11\]
rlabel metal1 11822 33524 11822 33524 0 outputs.divider_buffer\[12\]
rlabel metal1 15870 24922 15870 24922 0 outputs.divider_buffer\[13\]
rlabel metal1 18538 25262 18538 25262 0 outputs.divider_buffer\[14\]
rlabel metal1 21390 33388 21390 33388 0 outputs.divider_buffer\[15\]
rlabel metal2 20056 32980 20056 32980 0 outputs.divider_buffer\[16\]
rlabel metal2 22034 30532 22034 30532 0 outputs.divider_buffer\[17\]
rlabel metal1 21620 23494 21620 23494 0 outputs.divider_buffer\[1\]
rlabel metal1 18170 21862 18170 21862 0 outputs.divider_buffer\[2\]
rlabel metal1 20976 29138 20976 29138 0 outputs.divider_buffer\[3\]
rlabel metal1 20194 20570 20194 20570 0 outputs.divider_buffer\[4\]
rlabel metal1 18216 22406 18216 22406 0 outputs.divider_buffer\[5\]
rlabel metal1 19872 24310 19872 24310 0 outputs.divider_buffer\[6\]
rlabel metal1 13386 22610 13386 22610 0 outputs.divider_buffer\[7\]
rlabel metal1 20102 31246 20102 31246 0 outputs.divider_buffer\[8\]
rlabel metal2 11822 30464 11822 30464 0 outputs.divider_buffer\[9\]
rlabel metal1 43508 17306 43508 17306 0 outputs.output_gen.count\[0\]
rlabel metal2 44298 15164 44298 15164 0 outputs.output_gen.count\[1\]
rlabel metal1 42642 18836 42642 18836 0 outputs.output_gen.count\[2\]
rlabel metal1 42918 17102 42918 17102 0 outputs.output_gen.count\[3\]
rlabel metal1 40503 17306 40503 17306 0 outputs.output_gen.count\[4\]
rlabel metal1 40986 18700 40986 18700 0 outputs.output_gen.count\[5\]
rlabel metal1 38410 18666 38410 18666 0 outputs.output_gen.count\[6\]
rlabel metal1 39054 18156 39054 18156 0 outputs.output_gen.count\[7\]
rlabel metal1 42964 13362 42964 13362 0 outputs.output_gen.next_count\[0\]
rlabel metal1 42734 14926 42734 14926 0 outputs.output_gen.next_count\[1\]
rlabel metal1 42596 17578 42596 17578 0 outputs.output_gen.next_count\[2\]
rlabel metal1 41768 15674 41768 15674 0 outputs.output_gen.next_count\[3\]
rlabel metal2 40250 15708 40250 15708 0 outputs.output_gen.next_count\[4\]
rlabel metal1 39744 16762 39744 16762 0 outputs.output_gen.next_count\[5\]
rlabel metal2 37306 17884 37306 17884 0 outputs.output_gen.next_count\[6\]
rlabel metal1 37490 17238 37490 17238 0 outputs.output_gen.next_count\[7\]
rlabel metal1 42642 13838 42642 13838 0 outputs.output_gen.pwm_ff
rlabel metal1 40848 13498 40848 13498 0 outputs.output_gen.pwm_unff
rlabel metal1 43240 14518 43240 14518 0 outputs.pwm_output
rlabel metal1 36938 6766 36938 6766 0 outputs.sample_rate.count\[0\]
rlabel metal1 38042 7514 38042 7514 0 outputs.sample_rate.count\[1\]
rlabel metal1 37444 7854 37444 7854 0 outputs.sample_rate.count\[2\]
rlabel metal1 36478 8806 36478 8806 0 outputs.sample_rate.count\[3\]
rlabel metal1 35144 11730 35144 11730 0 outputs.sample_rate.count\[4\]
rlabel metal2 36478 11458 36478 11458 0 outputs.sample_rate.count\[5\]
rlabel metal1 36156 13838 36156 13838 0 outputs.sample_rate.count\[6\]
rlabel metal1 36938 14450 36938 14450 0 outputs.sample_rate.count\[7\]
rlabel metal1 35420 6426 35420 6426 0 outputs.sample_rate.next_count\[0\]
rlabel metal1 38410 6222 38410 6222 0 outputs.sample_rate.next_count\[1\]
rlabel metal1 36938 8398 36938 8398 0 outputs.sample_rate.next_count\[2\]
rlabel metal1 35512 8602 35512 8602 0 outputs.sample_rate.next_count\[3\]
rlabel metal1 33902 11186 33902 11186 0 outputs.sample_rate.next_count\[4\]
rlabel metal1 34904 11322 34904 11322 0 outputs.sample_rate.next_count\[5\]
rlabel metal1 35650 12954 35650 12954 0 outputs.sample_rate.next_count\[6\]
rlabel metal1 35420 15062 35420 15062 0 outputs.sample_rate.next_count\[7\]
rlabel metal1 42826 21556 42826 21556 0 outputs.scaled_buffer\[0\]
rlabel metal2 42918 21250 42918 21250 0 outputs.scaled_buffer\[1\]
rlabel metal1 43240 21658 43240 21658 0 outputs.scaled_buffer\[2\]
rlabel metal1 42826 23630 42826 23630 0 outputs.scaled_buffer\[3\]
rlabel metal1 41814 23766 41814 23766 0 outputs.scaled_buffer\[4\]
rlabel metal1 40250 22066 40250 22066 0 outputs.scaled_buffer\[5\]
rlabel metal1 39330 21590 39330 21590 0 outputs.scaled_buffer\[6\]
rlabel metal2 38318 20672 38318 20672 0 outputs.scaled_buffer\[7\]
rlabel metal2 20700 29988 20700 29988 0 outputs.shaper.count\[0\]
rlabel metal1 11454 39270 11454 39270 0 outputs.shaper.count\[10\]
rlabel metal1 12558 44846 12558 44846 0 outputs.shaper.count\[11\]
rlabel metal1 15180 44302 15180 44302 0 outputs.shaper.count\[12\]
rlabel metal1 17480 44370 17480 44370 0 outputs.shaper.count\[13\]
rlabel metal1 21022 43350 21022 43350 0 outputs.shaper.count\[14\]
rlabel metal1 20148 38930 20148 38930 0 outputs.shaper.count\[15\]
rlabel metal2 20746 33286 20746 33286 0 outputs.shaper.count\[16\]
rlabel metal1 21712 38182 21712 38182 0 outputs.shaper.count\[17\]
rlabel metal1 19550 27608 19550 27608 0 outputs.shaper.count\[1\]
rlabel metal1 21873 28050 21873 28050 0 outputs.shaper.count\[2\]
rlabel metal2 22770 33456 22770 33456 0 outputs.shaper.count\[3\]
rlabel metal1 18216 30022 18216 30022 0 outputs.shaper.count\[4\]
rlabel metal1 20424 35530 20424 35530 0 outputs.shaper.count\[5\]
rlabel metal1 20194 34918 20194 34918 0 outputs.shaper.count\[6\]
rlabel metal1 20516 35666 20516 35666 0 outputs.shaper.count\[7\]
rlabel metal1 13570 36040 13570 36040 0 outputs.shaper.count\[8\]
rlabel metal1 11730 36550 11730 36550 0 outputs.shaper.count\[9\]
rlabel metal1 13202 27472 13202 27472 0 outputs.sig_gen.count\[0\]
rlabel metal1 8924 33082 8924 33082 0 outputs.sig_gen.count\[10\]
rlabel via1 13017 28050 13017 28050 0 outputs.sig_gen.count\[11\]
rlabel metal1 10166 32334 10166 32334 0 outputs.sig_gen.count\[12\]
rlabel metal1 7222 36686 7222 36686 0 outputs.sig_gen.count\[13\]
rlabel metal2 15594 38148 15594 38148 0 outputs.sig_gen.count\[14\]
rlabel metal2 8694 36414 8694 36414 0 outputs.sig_gen.count\[15\]
rlabel metal1 14582 35088 14582 35088 0 outputs.sig_gen.count\[16\]
rlabel metal2 15916 33388 15916 33388 0 outputs.sig_gen.count\[17\]
rlabel metal1 13662 25874 13662 25874 0 outputs.sig_gen.count\[1\]
rlabel metal2 14950 27200 14950 27200 0 outputs.sig_gen.count\[2\]
rlabel metal1 16606 31790 16606 31790 0 outputs.sig_gen.count\[3\]
rlabel metal1 11270 28560 11270 28560 0 outputs.sig_gen.count\[4\]
rlabel metal1 15686 33354 15686 33354 0 outputs.sig_gen.count\[5\]
rlabel metal2 15410 30226 15410 30226 0 outputs.sig_gen.count\[6\]
rlabel metal1 7498 30022 7498 30022 0 outputs.sig_gen.count\[7\]
rlabel metal1 7498 31994 7498 31994 0 outputs.sig_gen.count\[8\]
rlabel metal1 8004 38862 8004 38862 0 outputs.sig_gen.count\[9\]
rlabel metal1 7774 25806 7774 25806 0 outputs.sig_gen.next_count\[0\]
rlabel metal1 7544 32538 7544 32538 0 outputs.sig_gen.next_count\[10\]
rlabel metal1 9522 31450 9522 31450 0 outputs.sig_gen.next_count\[11\]
rlabel metal2 4646 33252 4646 33252 0 outputs.sig_gen.next_count\[12\]
rlabel metal1 5290 36346 5290 36346 0 outputs.sig_gen.next_count\[13\]
rlabel metal1 5520 34986 5520 34986 0 outputs.sig_gen.next_count\[14\]
rlabel metal1 7360 35802 7360 35802 0 outputs.sig_gen.next_count\[15\]
rlabel metal1 9798 34986 9798 34986 0 outputs.sig_gen.next_count\[16\]
rlabel via1 9331 34374 9331 34374 0 outputs.sig_gen.next_count\[17\]
rlabel via1 10724 25466 10724 25466 0 outputs.sig_gen.next_count\[1\]
rlabel metal1 8694 27030 8694 27030 0 outputs.sig_gen.next_count\[2\]
rlabel metal1 9430 29206 9430 29206 0 outputs.sig_gen.next_count\[3\]
rlabel metal1 6660 27642 6660 27642 0 outputs.sig_gen.next_count\[4\]
rlabel metal1 5191 27642 5191 27642 0 outputs.sig_gen.next_count\[5\]
rlabel metal1 4140 29274 4140 29274 0 outputs.sig_gen.next_count\[6\]
rlabel metal1 5060 30770 5060 30770 0 outputs.sig_gen.next_count\[7\]
rlabel metal1 5796 31858 5796 31858 0 outputs.sig_gen.next_count\[8\]
rlabel metal1 8142 29818 8142 29818 0 outputs.sig_gen.next_count\[9\]
rlabel metal1 21206 25330 21206 25330 0 outputs.signal_buffer2\[0\]
rlabel metal1 11316 40562 11316 40562 0 outputs.signal_buffer2\[10\]
rlabel metal2 12926 44132 12926 44132 0 outputs.signal_buffer2\[11\]
rlabel metal1 14214 43418 14214 43418 0 outputs.signal_buffer2\[12\]
rlabel metal1 17112 43826 17112 43826 0 outputs.signal_buffer2\[13\]
rlabel metal1 19918 43384 19918 43384 0 outputs.signal_buffer2\[14\]
rlabel metal1 20286 40018 20286 40018 0 outputs.signal_buffer2\[15\]
rlabel metal1 22586 40698 22586 40698 0 outputs.signal_buffer2\[16\]
rlabel metal2 23598 38692 23598 38692 0 outputs.signal_buffer2\[17\]
rlabel metal1 18492 27098 18492 27098 0 outputs.signal_buffer2\[1\]
rlabel metal2 23046 28356 23046 28356 0 outputs.signal_buffer2\[2\]
rlabel metal2 22034 34068 22034 34068 0 outputs.signal_buffer2\[3\]
rlabel metal1 17480 29138 17480 29138 0 outputs.signal_buffer2\[4\]
rlabel metal2 21758 36788 21758 36788 0 outputs.signal_buffer2\[5\]
rlabel metal1 18722 35258 18722 35258 0 outputs.signal_buffer2\[6\]
rlabel metal1 18722 36788 18722 36788 0 outputs.signal_buffer2\[7\]
rlabel metal2 12282 37060 12282 37060 0 outputs.signal_buffer2\[8\]
rlabel metal1 11316 37978 11316 37978 0 outputs.signal_buffer2\[9\]
rlabel metal2 44206 15793 44206 15793 0 pwm
<< properties >>
string FIXED_BBOX 0 0 45733 47877
<< end >>
