VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO z23
  CLASS BLOCK ;
  FOREIGN z23 ;
  ORIGIN 0.000 0.000 ;
  SIZE 274.825 BY 285.545 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END clk
  PIN interrupt_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END interrupt_gpio_in
  PIN keypad_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END keypad_input[0]
  PIN keypad_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 3.440 274.825 4.040 ;
    END
  END keypad_input[10]
  PIN keypad_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END keypad_input[11]
  PIN keypad_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 281.545 261.190 285.545 ;
    END
  END keypad_input[12]
  PIN keypad_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END keypad_input[13]
  PIN keypad_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 78.240 274.825 78.840 ;
    END
  END keypad_input[14]
  PIN keypad_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END keypad_input[15]
  PIN keypad_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END keypad_input[1]
  PIN keypad_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END keypad_input[2]
  PIN keypad_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 281.545 190.350 285.545 ;
    END
  END keypad_input[3]
  PIN keypad_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END keypad_input[4]
  PIN keypad_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END keypad_input[5]
  PIN keypad_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 281.545 119.510 285.545 ;
    END
  END keypad_input[6]
  PIN keypad_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 51.040 274.825 51.640 ;
    END
  END keypad_input[7]
  PIN keypad_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 176.840 274.825 177.440 ;
    END
  END keypad_input[8]
  PIN keypad_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 281.545 235.430 285.545 ;
    END
  END keypad_input[9]
  PIN memory_address_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 281.545 267.630 285.545 ;
    END
  END memory_address_out[0]
  PIN memory_address_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 281.545 87.310 285.545 ;
    END
  END memory_address_out[10]
  PIN memory_address_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 281.545 142.050 285.545 ;
    END
  END memory_address_out[11]
  PIN memory_address_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 200.640 274.825 201.240 ;
    END
  END memory_address_out[12]
  PIN memory_address_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 251.250 281.545 251.530 285.545 ;
    END
  END memory_address_out[13]
  PIN memory_address_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 37.440 274.825 38.040 ;
    END
  END memory_address_out[14]
  PIN memory_address_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 228.710 281.545 228.990 285.545 ;
    END
  END memory_address_out[15]
  PIN memory_address_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END memory_address_out[1]
  PIN memory_address_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 217.640 274.825 218.240 ;
    END
  END memory_address_out[2]
  PIN memory_address_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 281.545 26.130 285.545 ;
    END
  END memory_address_out[3]
  PIN memory_address_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 281.545 158.150 285.545 ;
    END
  END memory_address_out[4]
  PIN memory_address_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END memory_address_out[5]
  PIN memory_address_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END memory_address_out[6]
  PIN memory_address_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 85.040 274.825 85.640 ;
    END
  END memory_address_out[7]
  PIN memory_address_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END memory_address_out[8]
  PIN memory_address_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END memory_address_out[9]
  PIN memory_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 125.840 274.825 126.440 ;
    END
  END memory_data_in[0]
  PIN memory_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END memory_data_in[1]
  PIN memory_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END memory_data_in[2]
  PIN memory_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 281.545 32.570 285.545 ;
    END
  END memory_data_in[3]
  PIN memory_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END memory_data_in[4]
  PIN memory_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 281.545 180.690 285.545 ;
    END
  END memory_data_in[5]
  PIN memory_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 281.545 135.610 285.545 ;
    END
  END memory_data_in[6]
  PIN memory_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 270.825 193.840 274.825 194.440 ;
    END
  END memory_data_in[7]
  PIN memory_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 227.840 274.825 228.440 ;
    END
  END memory_data_out[0]
  PIN memory_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END memory_data_out[1]
  PIN memory_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 119.040 274.825 119.640 ;
    END
  END memory_data_out[2]
  PIN memory_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END memory_data_out[3]
  PIN memory_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END memory_data_out[4]
  PIN memory_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END memory_data_out[5]
  PIN memory_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 10.240 274.825 10.840 ;
    END
  END memory_data_out[6]
  PIN memory_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END memory_data_out[7]
  PIN memory_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 153.040 274.825 153.640 ;
    END
  END memory_wr
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 281.545 222.550 285.545 ;
    END
  END nrst
  PIN programmable_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END programmable_gpio_in[0]
  PIN programmable_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END programmable_gpio_in[1]
  PIN programmable_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END programmable_gpio_in[2]
  PIN programmable_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 270.825 251.640 274.825 252.240 ;
    END
  END programmable_gpio_in[3]
  PIN programmable_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 270.825 95.240 274.825 95.840 ;
    END
  END programmable_gpio_in[4]
  PIN programmable_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 281.545 80.870 285.545 ;
    END
  END programmable_gpio_in[5]
  PIN programmable_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END programmable_gpio_in[6]
  PIN programmable_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END programmable_gpio_in[7]
  PIN programmable_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 281.545 113.070 285.545 ;
    END
  END programmable_gpio_out[0]
  PIN programmable_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END programmable_gpio_out[1]
  PIN programmable_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 234.640 274.825 235.240 ;
    END
  END programmable_gpio_out[2]
  PIN programmable_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 61.240 274.825 61.840 ;
    END
  END programmable_gpio_out[3]
  PIN programmable_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END programmable_gpio_out[4]
  PIN programmable_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END programmable_gpio_out[5]
  PIN programmable_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END programmable_gpio_out[6]
  PIN programmable_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END programmable_gpio_out[7]
  PIN programmable_gpio_wr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END programmable_gpio_wr[0]
  PIN programmable_gpio_wr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 170.040 274.825 170.640 ;
    END
  END programmable_gpio_wr[1]
  PIN programmable_gpio_wr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 281.545 58.330 285.545 ;
    END
  END programmable_gpio_wr[2]
  PIN programmable_gpio_wr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END programmable_gpio_wr[3]
  PIN programmable_gpio_wr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 268.640 274.825 269.240 ;
    END
  END programmable_gpio_wr[4]
  PIN programmable_gpio_wr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 281.545 125.950 285.545 ;
    END
  END programmable_gpio_wr[5]
  PIN programmable_gpio_wr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 281.545 10.030 285.545 ;
    END
  END programmable_gpio_wr[6]
  PIN programmable_gpio_wr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END programmable_gpio_wr[7]
  PIN ss0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 281.545 96.970 285.545 ;
    END
  END ss0[0]
  PIN ss0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 281.545 64.770 285.545 ;
    END
  END ss0[1]
  PIN ss0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 281.545 42.230 285.545 ;
    END
  END ss0[2]
  PIN ss0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 102.040 274.825 102.640 ;
    END
  END ss0[3]
  PIN ss0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 275.440 274.825 276.040 ;
    END
  END ss0[4]
  PIN ss0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END ss0[5]
  PIN ss0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 20.440 274.825 21.040 ;
    END
  END ss0[6]
  PIN ss0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 108.840 274.825 109.440 ;
    END
  END ss0[7]
  PIN ss1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.970 281.545 174.250 285.545 ;
    END
  END ss1[0]
  PIN ss1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 281.545 16.470 285.545 ;
    END
  END ss1[1]
  PIN ss1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END ss1[2]
  PIN ss1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END ss1[3]
  PIN ss1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END ss1[4]
  PIN ss1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 273.790 281.545 274.070 285.545 ;
    END
  END ss1[5]
  PIN ss1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END ss1[6]
  PIN ss1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END ss1[7]
  PIN ss2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END ss2[0]
  PIN ss2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END ss2[1]
  PIN ss2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 281.545 103.410 285.545 ;
    END
  END ss2[2]
  PIN ss2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END ss2[3]
  PIN ss2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END ss2[4]
  PIN ss2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END ss2[5]
  PIN ss2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 27.240 274.825 27.840 ;
    END
  END ss2[6]
  PIN ss2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 210.840 274.825 211.440 ;
    END
  END ss2[7]
  PIN ss3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 142.840 274.825 143.440 ;
    END
  END ss3[0]
  PIN ss3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END ss3[1]
  PIN ss3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END ss3[2]
  PIN ss3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 270.825 68.040 274.825 68.640 ;
    END
  END ss3[3]
  PIN ss3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END ss3[4]
  PIN ss3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 159.840 274.825 160.440 ;
    END
  END ss3[5]
  PIN ss3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 241.440 274.825 242.040 ;
    END
  END ss3[6]
  PIN ss3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END ss3[7]
  PIN ss4[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 258.440 274.825 259.040 ;
    END
  END ss4[0]
  PIN ss4[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END ss4[1]
  PIN ss4[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END ss4[2]
  PIN ss4[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END ss4[3]
  PIN ss4[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ss4[4]
  PIN ss4[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END ss4[5]
  PIN ss4[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END ss4[6]
  PIN ss4[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 281.545 71.210 285.545 ;
    END
  END ss4[7]
  PIN ss5[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 281.545 167.810 285.545 ;
    END
  END ss5[0]
  PIN ss5[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END ss5[1]
  PIN ss5[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END ss5[2]
  PIN ss5[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END ss5[3]
  PIN ss5[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 212.610 281.545 212.890 285.545 ;
    END
  END ss5[4]
  PIN ss5[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 281.545 151.710 285.545 ;
    END
  END ss5[5]
  PIN ss5[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END ss5[6]
  PIN ss5[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.810 281.545 245.090 285.545 ;
    END
  END ss5[7]
  PIN ss6[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 44.240 274.825 44.840 ;
    END
  END ss6[0]
  PIN ss6[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END ss6[1]
  PIN ss6[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ss6[2]
  PIN ss6[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END ss6[3]
  PIN ss6[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END ss6[4]
  PIN ss6[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END ss6[5]
  PIN ss6[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 183.640 274.825 184.240 ;
    END
  END ss6[6]
  PIN ss6[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END ss6[7]
  PIN ss7[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.170 281.545 206.450 285.545 ;
    END
  END ss7[0]
  PIN ss7[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.510 281.545 196.790 285.545 ;
    END
  END ss7[1]
  PIN ss7[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.310 281.545 3.590 285.545 ;
    END
  END ss7[2]
  PIN ss7[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 281.545 48.670 285.545 ;
    END
  END ss7[3]
  PIN ss7[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END ss7[4]
  PIN ss7[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END ss7[5]
  PIN ss7[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END ss7[6]
  PIN ss7[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 270.825 136.040 274.825 136.640 ;
    END
  END ss7[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 272.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 272.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 269.100 272.085 ;
      LAYER met1 ;
        RECT 0.070 8.880 274.090 274.680 ;
      LAYER met2 ;
        RECT 0.100 281.265 3.030 281.545 ;
        RECT 3.870 281.265 9.470 281.545 ;
        RECT 10.310 281.265 15.910 281.545 ;
        RECT 16.750 281.265 25.570 281.545 ;
        RECT 26.410 281.265 32.010 281.545 ;
        RECT 32.850 281.265 41.670 281.545 ;
        RECT 42.510 281.265 48.110 281.545 ;
        RECT 48.950 281.265 57.770 281.545 ;
        RECT 58.610 281.265 64.210 281.545 ;
        RECT 65.050 281.265 70.650 281.545 ;
        RECT 71.490 281.265 80.310 281.545 ;
        RECT 81.150 281.265 86.750 281.545 ;
        RECT 87.590 281.265 96.410 281.545 ;
        RECT 97.250 281.265 102.850 281.545 ;
        RECT 103.690 281.265 112.510 281.545 ;
        RECT 113.350 281.265 118.950 281.545 ;
        RECT 119.790 281.265 125.390 281.545 ;
        RECT 126.230 281.265 135.050 281.545 ;
        RECT 135.890 281.265 141.490 281.545 ;
        RECT 142.330 281.265 151.150 281.545 ;
        RECT 151.990 281.265 157.590 281.545 ;
        RECT 158.430 281.265 167.250 281.545 ;
        RECT 168.090 281.265 173.690 281.545 ;
        RECT 174.530 281.265 180.130 281.545 ;
        RECT 180.970 281.265 189.790 281.545 ;
        RECT 190.630 281.265 196.230 281.545 ;
        RECT 197.070 281.265 205.890 281.545 ;
        RECT 206.730 281.265 212.330 281.545 ;
        RECT 213.170 281.265 221.990 281.545 ;
        RECT 222.830 281.265 228.430 281.545 ;
        RECT 229.270 281.265 234.870 281.545 ;
        RECT 235.710 281.265 244.530 281.545 ;
        RECT 245.370 281.265 250.970 281.545 ;
        RECT 251.810 281.265 260.630 281.545 ;
        RECT 261.470 281.265 267.070 281.545 ;
        RECT 267.910 281.265 273.510 281.545 ;
        RECT 0.100 4.280 274.060 281.265 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 67.430 4.280 ;
        RECT 68.270 3.555 77.090 4.280 ;
        RECT 77.930 3.555 83.530 4.280 ;
        RECT 84.370 3.555 93.190 4.280 ;
        RECT 94.030 3.555 99.630 4.280 ;
        RECT 100.470 3.555 109.290 4.280 ;
        RECT 110.130 3.555 115.730 4.280 ;
        RECT 116.570 3.555 122.170 4.280 ;
        RECT 123.010 3.555 131.830 4.280 ;
        RECT 132.670 3.555 138.270 4.280 ;
        RECT 139.110 3.555 147.930 4.280 ;
        RECT 148.770 3.555 154.370 4.280 ;
        RECT 155.210 3.555 160.810 4.280 ;
        RECT 161.650 3.555 170.470 4.280 ;
        RECT 171.310 3.555 176.910 4.280 ;
        RECT 177.750 3.555 186.570 4.280 ;
        RECT 187.410 3.555 193.010 4.280 ;
        RECT 193.850 3.555 202.670 4.280 ;
        RECT 203.510 3.555 209.110 4.280 ;
        RECT 209.950 3.555 218.770 4.280 ;
        RECT 219.610 3.555 225.210 4.280 ;
        RECT 226.050 3.555 231.650 4.280 ;
        RECT 232.490 3.555 241.310 4.280 ;
        RECT 242.150 3.555 247.750 4.280 ;
        RECT 248.590 3.555 257.410 4.280 ;
        RECT 258.250 3.555 263.850 4.280 ;
        RECT 264.690 3.555 273.510 4.280 ;
      LAYER met3 ;
        RECT 4.400 278.440 273.635 279.305 ;
        RECT 4.000 276.440 273.635 278.440 ;
        RECT 4.000 275.040 270.425 276.440 ;
        RECT 4.000 273.040 273.635 275.040 ;
        RECT 4.400 271.640 273.635 273.040 ;
        RECT 4.000 269.640 273.635 271.640 ;
        RECT 4.000 268.240 270.425 269.640 ;
        RECT 4.000 262.840 273.635 268.240 ;
        RECT 4.400 261.440 273.635 262.840 ;
        RECT 4.000 259.440 273.635 261.440 ;
        RECT 4.000 258.040 270.425 259.440 ;
        RECT 4.000 256.040 273.635 258.040 ;
        RECT 4.400 254.640 273.635 256.040 ;
        RECT 4.000 252.640 273.635 254.640 ;
        RECT 4.000 251.240 270.425 252.640 ;
        RECT 4.000 245.840 273.635 251.240 ;
        RECT 4.400 244.440 273.635 245.840 ;
        RECT 4.000 242.440 273.635 244.440 ;
        RECT 4.000 241.040 270.425 242.440 ;
        RECT 4.000 239.040 273.635 241.040 ;
        RECT 4.400 237.640 273.635 239.040 ;
        RECT 4.000 235.640 273.635 237.640 ;
        RECT 4.000 234.240 270.425 235.640 ;
        RECT 4.000 228.840 273.635 234.240 ;
        RECT 4.400 227.440 270.425 228.840 ;
        RECT 4.000 222.040 273.635 227.440 ;
        RECT 4.400 220.640 273.635 222.040 ;
        RECT 4.000 218.640 273.635 220.640 ;
        RECT 4.000 217.240 270.425 218.640 ;
        RECT 4.000 215.240 273.635 217.240 ;
        RECT 4.400 213.840 273.635 215.240 ;
        RECT 4.000 211.840 273.635 213.840 ;
        RECT 4.000 210.440 270.425 211.840 ;
        RECT 4.000 205.040 273.635 210.440 ;
        RECT 4.400 203.640 273.635 205.040 ;
        RECT 4.000 201.640 273.635 203.640 ;
        RECT 4.000 200.240 270.425 201.640 ;
        RECT 4.000 198.240 273.635 200.240 ;
        RECT 4.400 196.840 273.635 198.240 ;
        RECT 4.000 194.840 273.635 196.840 ;
        RECT 4.000 193.440 270.425 194.840 ;
        RECT 4.000 188.040 273.635 193.440 ;
        RECT 4.400 186.640 273.635 188.040 ;
        RECT 4.000 184.640 273.635 186.640 ;
        RECT 4.000 183.240 270.425 184.640 ;
        RECT 4.000 181.240 273.635 183.240 ;
        RECT 4.400 179.840 273.635 181.240 ;
        RECT 4.000 177.840 273.635 179.840 ;
        RECT 4.000 176.440 270.425 177.840 ;
        RECT 4.000 171.040 273.635 176.440 ;
        RECT 4.400 169.640 270.425 171.040 ;
        RECT 4.000 164.240 273.635 169.640 ;
        RECT 4.400 162.840 273.635 164.240 ;
        RECT 4.000 160.840 273.635 162.840 ;
        RECT 4.000 159.440 270.425 160.840 ;
        RECT 4.000 157.440 273.635 159.440 ;
        RECT 4.400 156.040 273.635 157.440 ;
        RECT 4.000 154.040 273.635 156.040 ;
        RECT 4.000 152.640 270.425 154.040 ;
        RECT 4.000 147.240 273.635 152.640 ;
        RECT 4.400 145.840 273.635 147.240 ;
        RECT 4.000 143.840 273.635 145.840 ;
        RECT 4.000 142.440 270.425 143.840 ;
        RECT 4.000 140.440 273.635 142.440 ;
        RECT 4.400 139.040 273.635 140.440 ;
        RECT 4.000 137.040 273.635 139.040 ;
        RECT 4.000 135.640 270.425 137.040 ;
        RECT 4.000 130.240 273.635 135.640 ;
        RECT 4.400 128.840 273.635 130.240 ;
        RECT 4.000 126.840 273.635 128.840 ;
        RECT 4.000 125.440 270.425 126.840 ;
        RECT 4.000 123.440 273.635 125.440 ;
        RECT 4.400 122.040 273.635 123.440 ;
        RECT 4.000 120.040 273.635 122.040 ;
        RECT 4.000 118.640 270.425 120.040 ;
        RECT 4.000 113.240 273.635 118.640 ;
        RECT 4.400 111.840 273.635 113.240 ;
        RECT 4.000 109.840 273.635 111.840 ;
        RECT 4.000 108.440 270.425 109.840 ;
        RECT 4.000 106.440 273.635 108.440 ;
        RECT 4.400 105.040 273.635 106.440 ;
        RECT 4.000 103.040 273.635 105.040 ;
        RECT 4.000 101.640 270.425 103.040 ;
        RECT 4.000 99.640 273.635 101.640 ;
        RECT 4.400 98.240 273.635 99.640 ;
        RECT 4.000 96.240 273.635 98.240 ;
        RECT 4.000 94.840 270.425 96.240 ;
        RECT 4.000 89.440 273.635 94.840 ;
        RECT 4.400 88.040 273.635 89.440 ;
        RECT 4.000 86.040 273.635 88.040 ;
        RECT 4.000 84.640 270.425 86.040 ;
        RECT 4.000 82.640 273.635 84.640 ;
        RECT 4.400 81.240 273.635 82.640 ;
        RECT 4.000 79.240 273.635 81.240 ;
        RECT 4.000 77.840 270.425 79.240 ;
        RECT 4.000 72.440 273.635 77.840 ;
        RECT 4.400 71.040 273.635 72.440 ;
        RECT 4.000 69.040 273.635 71.040 ;
        RECT 4.000 67.640 270.425 69.040 ;
        RECT 4.000 65.640 273.635 67.640 ;
        RECT 4.400 64.240 273.635 65.640 ;
        RECT 4.000 62.240 273.635 64.240 ;
        RECT 4.000 60.840 270.425 62.240 ;
        RECT 4.000 55.440 273.635 60.840 ;
        RECT 4.400 54.040 273.635 55.440 ;
        RECT 4.000 52.040 273.635 54.040 ;
        RECT 4.000 50.640 270.425 52.040 ;
        RECT 4.000 48.640 273.635 50.640 ;
        RECT 4.400 47.240 273.635 48.640 ;
        RECT 4.000 45.240 273.635 47.240 ;
        RECT 4.000 43.840 270.425 45.240 ;
        RECT 4.000 41.840 273.635 43.840 ;
        RECT 4.400 40.440 273.635 41.840 ;
        RECT 4.000 38.440 273.635 40.440 ;
        RECT 4.000 37.040 270.425 38.440 ;
        RECT 4.000 31.640 273.635 37.040 ;
        RECT 4.400 30.240 273.635 31.640 ;
        RECT 4.000 28.240 273.635 30.240 ;
        RECT 4.000 26.840 270.425 28.240 ;
        RECT 4.000 24.840 273.635 26.840 ;
        RECT 4.400 23.440 273.635 24.840 ;
        RECT 4.000 21.440 273.635 23.440 ;
        RECT 4.000 20.040 270.425 21.440 ;
        RECT 4.000 14.640 273.635 20.040 ;
        RECT 4.400 13.240 273.635 14.640 ;
        RECT 4.000 11.240 273.635 13.240 ;
        RECT 4.000 9.840 270.425 11.240 ;
        RECT 4.000 7.840 273.635 9.840 ;
        RECT 4.400 6.440 273.635 7.840 ;
        RECT 4.000 4.440 273.635 6.440 ;
        RECT 4.000 3.575 270.425 4.440 ;
      LAYER met4 ;
        RECT 33.415 11.055 97.440 270.465 ;
        RECT 99.840 11.055 174.240 270.465 ;
        RECT 176.640 11.055 251.040 270.465 ;
        RECT 253.440 11.055 261.905 270.465 ;
  END
END z23
END LIBRARY

